/* modified netlist. Source: module AES in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/5-AES_EncRoundBased_PortParallel/4-AGEMA/AES.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module AES_SAUBER_Pipeline_d1 (plaintext_s0_t, key_s0_t, start_t, start_f, key_s0_f, key_s1_t, key_s1_f, plaintext_s0_f, plaintext_s1_t, plaintext_s1_f, ciphertext_s0_t, done_t, ciphertext_s0_f, ciphertext_s1_t, ciphertext_s1_f, done_f);
    input [127:0] plaintext_s0_t ;
    input [127:0] key_s0_t ;
    input start_t ;
    input start_f ;
    input [127:0] key_s0_f ;
    input [127:0] key_s1_t ;
    input [127:0] key_s1_f ;
    input [127:0] plaintext_s0_f ;
    input [127:0] plaintext_s1_t ;
    input [127:0] plaintext_s1_f ;
    output [127:0] ciphertext_s0_t ;
    output done_t ;
    output [127:0] ciphertext_s0_f ;
    output [127:0] ciphertext_s1_t ;
    output [127:0] ciphertext_s1_f ;
    output done_f ;
    wire n283 ;
    wire n285 ;
    wire n577 ;
    wire n585 ;
    wire n586 ;
    wire n588 ;
    wire n589 ;
    wire n591 ;
    wire n592 ;
    wire n593 ;
    wire n594 ;
    wire n595 ;
    wire n596 ;
    wire n597 ;
    wire n598 ;
    wire n599 ;
    wire n600 ;
    wire n601 ;
    wire n602 ;
    wire n603 ;
    wire n604 ;
    wire n605 ;
    wire n606 ;
    wire n607 ;
    wire n608 ;
    wire n609 ;
    wire n610 ;
    wire n611 ;
    wire n612 ;
    wire n613 ;
    wire n614 ;
    wire n615 ;
    wire n616 ;
    wire n617 ;
    wire n618 ;
    wire n619 ;
    wire n620 ;
    wire n621 ;
    wire n622 ;
    wire n623 ;
    wire n624 ;
    wire n625 ;
    wire n626 ;
    wire n627 ;
    wire n628 ;
    wire n629 ;
    wire n630 ;
    wire n631 ;
    wire n632 ;
    wire n633 ;
    wire n634 ;
    wire n635 ;
    wire n636 ;
    wire n637 ;
    wire n638 ;
    wire n639 ;
    wire n640 ;
    wire n641 ;
    wire n642 ;
    wire n643 ;
    wire n644 ;
    wire n645 ;
    wire n646 ;
    wire n647 ;
    wire n648 ;
    wire n649 ;
    wire n650 ;
    wire n651 ;
    wire n652 ;
    wire n653 ;
    wire n654 ;
    wire n655 ;
    wire n656 ;
    wire n657 ;
    wire n658 ;
    wire n659 ;
    wire n660 ;
    wire n661 ;
    wire n662 ;
    wire n663 ;
    wire n664 ;
    wire n665 ;
    wire n666 ;
    wire n667 ;
    wire n668 ;
    wire n669 ;
    wire n670 ;
    wire n671 ;
    wire n672 ;
    wire n673 ;
    wire n674 ;
    wire n675 ;
    wire n676 ;
    wire n677 ;
    wire n678 ;
    wire n679 ;
    wire n680 ;
    wire n681 ;
    wire n682 ;
    wire n683 ;
    wire n684 ;
    wire n685 ;
    wire n686 ;
    wire n687 ;
    wire n688 ;
    wire n689 ;
    wire n690 ;
    wire n691 ;
    wire n692 ;
    wire n693 ;
    wire n694 ;
    wire n695 ;
    wire n696 ;
    wire n697 ;
    wire n698 ;
    wire n699 ;
    wire n700 ;
    wire n701 ;
    wire n702 ;
    wire n703 ;
    wire n704 ;
    wire n705 ;
    wire n706 ;
    wire n707 ;
    wire n708 ;
    wire n709 ;
    wire n710 ;
    wire n711 ;
    wire n712 ;
    wire n713 ;
    wire n714 ;
    wire n715 ;
    wire n716 ;
    wire n717 ;
    wire n718 ;
    wire n719 ;
    wire n720 ;
    wire n721 ;
    wire n722 ;
    wire n723 ;
    wire n724 ;
    wire n725 ;
    wire n726 ;
    wire n727 ;
    wire n728 ;
    wire n729 ;
    wire n730 ;
    wire n731 ;
    wire n732 ;
    wire n733 ;
    wire n734 ;
    wire n735 ;
    wire n736 ;
    wire n737 ;
    wire n738 ;
    wire n739 ;
    wire n740 ;
    wire n741 ;
    wire n742 ;
    wire n743 ;
    wire n744 ;
    wire n745 ;
    wire n746 ;
    wire n747 ;
    wire n748 ;
    wire n749 ;
    wire n750 ;
    wire n751 ;
    wire n752 ;
    wire n753 ;
    wire n754 ;
    wire n755 ;
    wire n756 ;
    wire n757 ;
    wire n758 ;
    wire n759 ;
    wire n760 ;
    wire n761 ;
    wire n762 ;
    wire n763 ;
    wire n764 ;
    wire n765 ;
    wire n766 ;
    wire n767 ;
    wire n768 ;
    wire n769 ;
    wire n770 ;
    wire n771 ;
    wire n772 ;
    wire n773 ;
    wire n774 ;
    wire n775 ;
    wire n776 ;
    wire n777 ;
    wire n778 ;
    wire n779 ;
    wire n780 ;
    wire n781 ;
    wire n782 ;
    wire n783 ;
    wire n784 ;
    wire n785 ;
    wire n786 ;
    wire n787 ;
    wire n788 ;
    wire n789 ;
    wire n790 ;
    wire n791 ;
    wire n792 ;
    wire n793 ;
    wire n794 ;
    wire n795 ;
    wire n796 ;
    wire n797 ;
    wire n798 ;
    wire n799 ;
    wire n800 ;
    wire n801 ;
    wire n802 ;
    wire n803 ;
    wire n804 ;
    wire n805 ;
    wire n806 ;
    wire n807 ;
    wire n808 ;
    wire n809 ;
    wire n810 ;
    wire n811 ;
    wire n812 ;
    wire n813 ;
    wire n814 ;
    wire n815 ;
    wire n816 ;
    wire n817 ;
    wire n818 ;
    wire n819 ;
    wire n820 ;
    wire n821 ;
    wire n822 ;
    wire n823 ;
    wire n824 ;
    wire n825 ;
    wire n826 ;
    wire n827 ;
    wire n828 ;
    wire n829 ;
    wire n830 ;
    wire n831 ;
    wire n832 ;
    wire n833 ;
    wire n834 ;
    wire n835 ;
    wire n836 ;
    wire n837 ;
    wire n838 ;
    wire n839 ;
    wire n840 ;
    wire n841 ;
    wire n842 ;
    wire n843 ;
    wire n844 ;
    wire n845 ;
    wire n846 ;
    wire n847 ;
    wire n848 ;
    wire n849 ;
    wire n850 ;
    wire n851 ;
    wire n852 ;
    wire n853 ;
    wire n855 ;
    wire n856 ;
    wire RoundReg_Inst_ff_SDE_0_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_0_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_1_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_1_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_2_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_2_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_3_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_3_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_4_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_4_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_5_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_5_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_6_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_6_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_7_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_7_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_8_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_8_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_9_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_9_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_10_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_10_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_11_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_11_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_12_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_12_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_13_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_13_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_14_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_14_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_15_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_15_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_16_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_16_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_17_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_17_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_18_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_18_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_19_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_19_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_20_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_20_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_21_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_21_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_22_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_22_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_23_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_23_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_24_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_24_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_25_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_25_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_26_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_26_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_27_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_27_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_28_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_28_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_29_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_29_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_30_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_30_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_31_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_31_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_32_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_32_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_33_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_33_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_34_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_34_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_35_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_35_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_36_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_36_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_37_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_37_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_38_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_38_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_39_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_39_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_40_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_40_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_41_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_41_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_42_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_42_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_43_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_43_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_44_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_44_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_45_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_45_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_46_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_46_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_47_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_47_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_48_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_48_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_49_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_49_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_50_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_50_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_51_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_51_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_52_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_52_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_53_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_53_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_54_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_54_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_55_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_55_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_56_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_56_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_57_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_57_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_58_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_58_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_59_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_59_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_60_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_60_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_61_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_61_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_62_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_62_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_63_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_63_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_64_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_64_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_65_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_65_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_66_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_66_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_67_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_67_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_68_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_68_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_69_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_69_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_70_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_70_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_71_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_71_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_72_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_72_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_73_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_73_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_74_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_74_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_75_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_75_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_76_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_76_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_77_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_77_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_78_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_78_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_79_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_79_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_80_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_80_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_81_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_81_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_82_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_82_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_83_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_83_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_84_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_84_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_85_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_85_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_86_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_86_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_87_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_87_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_88_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_88_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_89_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_89_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_90_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_90_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_91_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_91_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_92_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_92_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_93_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_93_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_94_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_94_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_95_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_95_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_96_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_96_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_97_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_97_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_98_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_98_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_99_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_99_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_100_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_100_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_101_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_101_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_102_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_102_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_103_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_103_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_104_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_104_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_105_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_105_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_106_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_106_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_107_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_107_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_108_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_108_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_109_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_109_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_110_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_110_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_111_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_111_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_112_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_112_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_113_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_113_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_114_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_114_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_115_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_115_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_116_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_116_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_117_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_117_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_118_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_118_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_119_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_119_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_120_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_120_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_121_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_121_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_122_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_122_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_123_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_123_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_124_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_124_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_125_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_125_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_126_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_126_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_127_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_127_MUX_inst_X ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire SubBytesIns_Inst_Sbox_4_L29 ;
    wire SubBytesIns_Inst_Sbox_4_L28 ;
    wire SubBytesIns_Inst_Sbox_4_L27 ;
    wire SubBytesIns_Inst_Sbox_4_L26 ;
    wire SubBytesIns_Inst_Sbox_4_L25 ;
    wire SubBytesIns_Inst_Sbox_4_L24 ;
    wire SubBytesIns_Inst_Sbox_4_L23 ;
    wire SubBytesIns_Inst_Sbox_4_L22 ;
    wire SubBytesIns_Inst_Sbox_4_L21 ;
    wire SubBytesIns_Inst_Sbox_4_L20 ;
    wire SubBytesIns_Inst_Sbox_4_L19 ;
    wire SubBytesIns_Inst_Sbox_4_L18 ;
    wire SubBytesIns_Inst_Sbox_4_L17 ;
    wire SubBytesIns_Inst_Sbox_4_L16 ;
    wire SubBytesIns_Inst_Sbox_4_L15 ;
    wire SubBytesIns_Inst_Sbox_4_L14 ;
    wire SubBytesIns_Inst_Sbox_4_L13 ;
    wire SubBytesIns_Inst_Sbox_4_L12 ;
    wire SubBytesIns_Inst_Sbox_4_L11 ;
    wire SubBytesIns_Inst_Sbox_4_L10 ;
    wire SubBytesIns_Inst_Sbox_4_L9 ;
    wire SubBytesIns_Inst_Sbox_4_L8 ;
    wire SubBytesIns_Inst_Sbox_4_L7 ;
    wire SubBytesIns_Inst_Sbox_4_L6 ;
    wire SubBytesIns_Inst_Sbox_4_L5 ;
    wire SubBytesIns_Inst_Sbox_4_L4 ;
    wire SubBytesIns_Inst_Sbox_4_L3 ;
    wire SubBytesIns_Inst_Sbox_4_L2 ;
    wire SubBytesIns_Inst_Sbox_4_L1 ;
    wire SubBytesIns_Inst_Sbox_4_L0 ;
    wire SubBytesIns_Inst_Sbox_4_M63 ;
    wire SubBytesIns_Inst_Sbox_4_M62 ;
    wire SubBytesIns_Inst_Sbox_4_M61 ;
    wire SubBytesIns_Inst_Sbox_4_M60 ;
    wire SubBytesIns_Inst_Sbox_4_M59 ;
    wire SubBytesIns_Inst_Sbox_4_M58 ;
    wire SubBytesIns_Inst_Sbox_4_M57 ;
    wire SubBytesIns_Inst_Sbox_4_M56 ;
    wire SubBytesIns_Inst_Sbox_4_M55 ;
    wire SubBytesIns_Inst_Sbox_4_M54 ;
    wire SubBytesIns_Inst_Sbox_4_M53 ;
    wire SubBytesIns_Inst_Sbox_4_M52 ;
    wire SubBytesIns_Inst_Sbox_4_M51 ;
    wire SubBytesIns_Inst_Sbox_4_M50 ;
    wire SubBytesIns_Inst_Sbox_4_M49 ;
    wire SubBytesIns_Inst_Sbox_4_M48 ;
    wire SubBytesIns_Inst_Sbox_4_M47 ;
    wire SubBytesIns_Inst_Sbox_4_M46 ;
    wire SubBytesIns_Inst_Sbox_4_M45 ;
    wire SubBytesIns_Inst_Sbox_4_M44 ;
    wire SubBytesIns_Inst_Sbox_4_M43 ;
    wire SubBytesIns_Inst_Sbox_4_M42 ;
    wire SubBytesIns_Inst_Sbox_4_M41 ;
    wire SubBytesIns_Inst_Sbox_4_M40 ;
    wire SubBytesIns_Inst_Sbox_4_M39 ;
    wire SubBytesIns_Inst_Sbox_4_M38 ;
    wire SubBytesIns_Inst_Sbox_4_M37 ;
    wire SubBytesIns_Inst_Sbox_4_M36 ;
    wire SubBytesIns_Inst_Sbox_4_M35 ;
    wire SubBytesIns_Inst_Sbox_4_M34 ;
    wire SubBytesIns_Inst_Sbox_4_M33 ;
    wire SubBytesIns_Inst_Sbox_4_M32 ;
    wire SubBytesIns_Inst_Sbox_4_M31 ;
    wire SubBytesIns_Inst_Sbox_4_M30 ;
    wire SubBytesIns_Inst_Sbox_4_M29 ;
    wire SubBytesIns_Inst_Sbox_4_M28 ;
    wire SubBytesIns_Inst_Sbox_4_M27 ;
    wire SubBytesIns_Inst_Sbox_4_M26 ;
    wire SubBytesIns_Inst_Sbox_4_M25 ;
    wire SubBytesIns_Inst_Sbox_4_M24 ;
    wire SubBytesIns_Inst_Sbox_4_M23 ;
    wire SubBytesIns_Inst_Sbox_4_M22 ;
    wire SubBytesIns_Inst_Sbox_4_M21 ;
    wire SubBytesIns_Inst_Sbox_4_M20 ;
    wire SubBytesIns_Inst_Sbox_4_M19 ;
    wire SubBytesIns_Inst_Sbox_4_M18 ;
    wire SubBytesIns_Inst_Sbox_4_M17 ;
    wire SubBytesIns_Inst_Sbox_4_M16 ;
    wire SubBytesIns_Inst_Sbox_4_M15 ;
    wire SubBytesIns_Inst_Sbox_4_M14 ;
    wire SubBytesIns_Inst_Sbox_4_M13 ;
    wire SubBytesIns_Inst_Sbox_4_M12 ;
    wire SubBytesIns_Inst_Sbox_4_M11 ;
    wire SubBytesIns_Inst_Sbox_4_M10 ;
    wire SubBytesIns_Inst_Sbox_4_M9 ;
    wire SubBytesIns_Inst_Sbox_4_M8 ;
    wire SubBytesIns_Inst_Sbox_4_M7 ;
    wire SubBytesIns_Inst_Sbox_4_M6 ;
    wire SubBytesIns_Inst_Sbox_4_M5 ;
    wire SubBytesIns_Inst_Sbox_4_M4 ;
    wire SubBytesIns_Inst_Sbox_4_M3 ;
    wire SubBytesIns_Inst_Sbox_4_M2 ;
    wire SubBytesIns_Inst_Sbox_4_M1 ;
    wire SubBytesIns_Inst_Sbox_4_T27 ;
    wire SubBytesIns_Inst_Sbox_4_T26 ;
    wire SubBytesIns_Inst_Sbox_4_T25 ;
    wire SubBytesIns_Inst_Sbox_4_T24 ;
    wire SubBytesIns_Inst_Sbox_4_T23 ;
    wire SubBytesIns_Inst_Sbox_4_T22 ;
    wire SubBytesIns_Inst_Sbox_4_T21 ;
    wire SubBytesIns_Inst_Sbox_4_T20 ;
    wire SubBytesIns_Inst_Sbox_4_T19 ;
    wire SubBytesIns_Inst_Sbox_4_T18 ;
    wire SubBytesIns_Inst_Sbox_4_T17 ;
    wire SubBytesIns_Inst_Sbox_4_T16 ;
    wire SubBytesIns_Inst_Sbox_4_T15 ;
    wire SubBytesIns_Inst_Sbox_4_T14 ;
    wire SubBytesIns_Inst_Sbox_4_T13 ;
    wire SubBytesIns_Inst_Sbox_4_T12 ;
    wire SubBytesIns_Inst_Sbox_4_T11 ;
    wire SubBytesIns_Inst_Sbox_4_T10 ;
    wire SubBytesIns_Inst_Sbox_4_T9 ;
    wire SubBytesIns_Inst_Sbox_4_T8 ;
    wire SubBytesIns_Inst_Sbox_4_T7 ;
    wire SubBytesIns_Inst_Sbox_4_T6 ;
    wire SubBytesIns_Inst_Sbox_4_T5 ;
    wire SubBytesIns_Inst_Sbox_4_T4 ;
    wire SubBytesIns_Inst_Sbox_4_T3 ;
    wire SubBytesIns_Inst_Sbox_4_T2 ;
    wire SubBytesIns_Inst_Sbox_4_T1 ;
    wire SubBytesIns_Inst_Sbox_5_L29 ;
    wire SubBytesIns_Inst_Sbox_5_L28 ;
    wire SubBytesIns_Inst_Sbox_5_L27 ;
    wire SubBytesIns_Inst_Sbox_5_L26 ;
    wire SubBytesIns_Inst_Sbox_5_L25 ;
    wire SubBytesIns_Inst_Sbox_5_L24 ;
    wire SubBytesIns_Inst_Sbox_5_L23 ;
    wire SubBytesIns_Inst_Sbox_5_L22 ;
    wire SubBytesIns_Inst_Sbox_5_L21 ;
    wire SubBytesIns_Inst_Sbox_5_L20 ;
    wire SubBytesIns_Inst_Sbox_5_L19 ;
    wire SubBytesIns_Inst_Sbox_5_L18 ;
    wire SubBytesIns_Inst_Sbox_5_L17 ;
    wire SubBytesIns_Inst_Sbox_5_L16 ;
    wire SubBytesIns_Inst_Sbox_5_L15 ;
    wire SubBytesIns_Inst_Sbox_5_L14 ;
    wire SubBytesIns_Inst_Sbox_5_L13 ;
    wire SubBytesIns_Inst_Sbox_5_L12 ;
    wire SubBytesIns_Inst_Sbox_5_L11 ;
    wire SubBytesIns_Inst_Sbox_5_L10 ;
    wire SubBytesIns_Inst_Sbox_5_L9 ;
    wire SubBytesIns_Inst_Sbox_5_L8 ;
    wire SubBytesIns_Inst_Sbox_5_L7 ;
    wire SubBytesIns_Inst_Sbox_5_L6 ;
    wire SubBytesIns_Inst_Sbox_5_L5 ;
    wire SubBytesIns_Inst_Sbox_5_L4 ;
    wire SubBytesIns_Inst_Sbox_5_L3 ;
    wire SubBytesIns_Inst_Sbox_5_L2 ;
    wire SubBytesIns_Inst_Sbox_5_L1 ;
    wire SubBytesIns_Inst_Sbox_5_L0 ;
    wire SubBytesIns_Inst_Sbox_5_M63 ;
    wire SubBytesIns_Inst_Sbox_5_M62 ;
    wire SubBytesIns_Inst_Sbox_5_M61 ;
    wire SubBytesIns_Inst_Sbox_5_M60 ;
    wire SubBytesIns_Inst_Sbox_5_M59 ;
    wire SubBytesIns_Inst_Sbox_5_M58 ;
    wire SubBytesIns_Inst_Sbox_5_M57 ;
    wire SubBytesIns_Inst_Sbox_5_M56 ;
    wire SubBytesIns_Inst_Sbox_5_M55 ;
    wire SubBytesIns_Inst_Sbox_5_M54 ;
    wire SubBytesIns_Inst_Sbox_5_M53 ;
    wire SubBytesIns_Inst_Sbox_5_M52 ;
    wire SubBytesIns_Inst_Sbox_5_M51 ;
    wire SubBytesIns_Inst_Sbox_5_M50 ;
    wire SubBytesIns_Inst_Sbox_5_M49 ;
    wire SubBytesIns_Inst_Sbox_5_M48 ;
    wire SubBytesIns_Inst_Sbox_5_M47 ;
    wire SubBytesIns_Inst_Sbox_5_M46 ;
    wire SubBytesIns_Inst_Sbox_5_M45 ;
    wire SubBytesIns_Inst_Sbox_5_M44 ;
    wire SubBytesIns_Inst_Sbox_5_M43 ;
    wire SubBytesIns_Inst_Sbox_5_M42 ;
    wire SubBytesIns_Inst_Sbox_5_M41 ;
    wire SubBytesIns_Inst_Sbox_5_M40 ;
    wire SubBytesIns_Inst_Sbox_5_M39 ;
    wire SubBytesIns_Inst_Sbox_5_M38 ;
    wire SubBytesIns_Inst_Sbox_5_M37 ;
    wire SubBytesIns_Inst_Sbox_5_M36 ;
    wire SubBytesIns_Inst_Sbox_5_M35 ;
    wire SubBytesIns_Inst_Sbox_5_M34 ;
    wire SubBytesIns_Inst_Sbox_5_M33 ;
    wire SubBytesIns_Inst_Sbox_5_M32 ;
    wire SubBytesIns_Inst_Sbox_5_M31 ;
    wire SubBytesIns_Inst_Sbox_5_M30 ;
    wire SubBytesIns_Inst_Sbox_5_M29 ;
    wire SubBytesIns_Inst_Sbox_5_M28 ;
    wire SubBytesIns_Inst_Sbox_5_M27 ;
    wire SubBytesIns_Inst_Sbox_5_M26 ;
    wire SubBytesIns_Inst_Sbox_5_M25 ;
    wire SubBytesIns_Inst_Sbox_5_M24 ;
    wire SubBytesIns_Inst_Sbox_5_M23 ;
    wire SubBytesIns_Inst_Sbox_5_M22 ;
    wire SubBytesIns_Inst_Sbox_5_M21 ;
    wire SubBytesIns_Inst_Sbox_5_M20 ;
    wire SubBytesIns_Inst_Sbox_5_M19 ;
    wire SubBytesIns_Inst_Sbox_5_M18 ;
    wire SubBytesIns_Inst_Sbox_5_M17 ;
    wire SubBytesIns_Inst_Sbox_5_M16 ;
    wire SubBytesIns_Inst_Sbox_5_M15 ;
    wire SubBytesIns_Inst_Sbox_5_M14 ;
    wire SubBytesIns_Inst_Sbox_5_M13 ;
    wire SubBytesIns_Inst_Sbox_5_M12 ;
    wire SubBytesIns_Inst_Sbox_5_M11 ;
    wire SubBytesIns_Inst_Sbox_5_M10 ;
    wire SubBytesIns_Inst_Sbox_5_M9 ;
    wire SubBytesIns_Inst_Sbox_5_M8 ;
    wire SubBytesIns_Inst_Sbox_5_M7 ;
    wire SubBytesIns_Inst_Sbox_5_M6 ;
    wire SubBytesIns_Inst_Sbox_5_M5 ;
    wire SubBytesIns_Inst_Sbox_5_M4 ;
    wire SubBytesIns_Inst_Sbox_5_M3 ;
    wire SubBytesIns_Inst_Sbox_5_M2 ;
    wire SubBytesIns_Inst_Sbox_5_M1 ;
    wire SubBytesIns_Inst_Sbox_5_T27 ;
    wire SubBytesIns_Inst_Sbox_5_T26 ;
    wire SubBytesIns_Inst_Sbox_5_T25 ;
    wire SubBytesIns_Inst_Sbox_5_T24 ;
    wire SubBytesIns_Inst_Sbox_5_T23 ;
    wire SubBytesIns_Inst_Sbox_5_T22 ;
    wire SubBytesIns_Inst_Sbox_5_T21 ;
    wire SubBytesIns_Inst_Sbox_5_T20 ;
    wire SubBytesIns_Inst_Sbox_5_T19 ;
    wire SubBytesIns_Inst_Sbox_5_T18 ;
    wire SubBytesIns_Inst_Sbox_5_T17 ;
    wire SubBytesIns_Inst_Sbox_5_T16 ;
    wire SubBytesIns_Inst_Sbox_5_T15 ;
    wire SubBytesIns_Inst_Sbox_5_T14 ;
    wire SubBytesIns_Inst_Sbox_5_T13 ;
    wire SubBytesIns_Inst_Sbox_5_T12 ;
    wire SubBytesIns_Inst_Sbox_5_T11 ;
    wire SubBytesIns_Inst_Sbox_5_T10 ;
    wire SubBytesIns_Inst_Sbox_5_T9 ;
    wire SubBytesIns_Inst_Sbox_5_T8 ;
    wire SubBytesIns_Inst_Sbox_5_T7 ;
    wire SubBytesIns_Inst_Sbox_5_T6 ;
    wire SubBytesIns_Inst_Sbox_5_T5 ;
    wire SubBytesIns_Inst_Sbox_5_T4 ;
    wire SubBytesIns_Inst_Sbox_5_T3 ;
    wire SubBytesIns_Inst_Sbox_5_T2 ;
    wire SubBytesIns_Inst_Sbox_5_T1 ;
    wire SubBytesIns_Inst_Sbox_6_L29 ;
    wire SubBytesIns_Inst_Sbox_6_L28 ;
    wire SubBytesIns_Inst_Sbox_6_L27 ;
    wire SubBytesIns_Inst_Sbox_6_L26 ;
    wire SubBytesIns_Inst_Sbox_6_L25 ;
    wire SubBytesIns_Inst_Sbox_6_L24 ;
    wire SubBytesIns_Inst_Sbox_6_L23 ;
    wire SubBytesIns_Inst_Sbox_6_L22 ;
    wire SubBytesIns_Inst_Sbox_6_L21 ;
    wire SubBytesIns_Inst_Sbox_6_L20 ;
    wire SubBytesIns_Inst_Sbox_6_L19 ;
    wire SubBytesIns_Inst_Sbox_6_L18 ;
    wire SubBytesIns_Inst_Sbox_6_L17 ;
    wire SubBytesIns_Inst_Sbox_6_L16 ;
    wire SubBytesIns_Inst_Sbox_6_L15 ;
    wire SubBytesIns_Inst_Sbox_6_L14 ;
    wire SubBytesIns_Inst_Sbox_6_L13 ;
    wire SubBytesIns_Inst_Sbox_6_L12 ;
    wire SubBytesIns_Inst_Sbox_6_L11 ;
    wire SubBytesIns_Inst_Sbox_6_L10 ;
    wire SubBytesIns_Inst_Sbox_6_L9 ;
    wire SubBytesIns_Inst_Sbox_6_L8 ;
    wire SubBytesIns_Inst_Sbox_6_L7 ;
    wire SubBytesIns_Inst_Sbox_6_L6 ;
    wire SubBytesIns_Inst_Sbox_6_L5 ;
    wire SubBytesIns_Inst_Sbox_6_L4 ;
    wire SubBytesIns_Inst_Sbox_6_L3 ;
    wire SubBytesIns_Inst_Sbox_6_L2 ;
    wire SubBytesIns_Inst_Sbox_6_L1 ;
    wire SubBytesIns_Inst_Sbox_6_L0 ;
    wire SubBytesIns_Inst_Sbox_6_M63 ;
    wire SubBytesIns_Inst_Sbox_6_M62 ;
    wire SubBytesIns_Inst_Sbox_6_M61 ;
    wire SubBytesIns_Inst_Sbox_6_M60 ;
    wire SubBytesIns_Inst_Sbox_6_M59 ;
    wire SubBytesIns_Inst_Sbox_6_M58 ;
    wire SubBytesIns_Inst_Sbox_6_M57 ;
    wire SubBytesIns_Inst_Sbox_6_M56 ;
    wire SubBytesIns_Inst_Sbox_6_M55 ;
    wire SubBytesIns_Inst_Sbox_6_M54 ;
    wire SubBytesIns_Inst_Sbox_6_M53 ;
    wire SubBytesIns_Inst_Sbox_6_M52 ;
    wire SubBytesIns_Inst_Sbox_6_M51 ;
    wire SubBytesIns_Inst_Sbox_6_M50 ;
    wire SubBytesIns_Inst_Sbox_6_M49 ;
    wire SubBytesIns_Inst_Sbox_6_M48 ;
    wire SubBytesIns_Inst_Sbox_6_M47 ;
    wire SubBytesIns_Inst_Sbox_6_M46 ;
    wire SubBytesIns_Inst_Sbox_6_M45 ;
    wire SubBytesIns_Inst_Sbox_6_M44 ;
    wire SubBytesIns_Inst_Sbox_6_M43 ;
    wire SubBytesIns_Inst_Sbox_6_M42 ;
    wire SubBytesIns_Inst_Sbox_6_M41 ;
    wire SubBytesIns_Inst_Sbox_6_M40 ;
    wire SubBytesIns_Inst_Sbox_6_M39 ;
    wire SubBytesIns_Inst_Sbox_6_M38 ;
    wire SubBytesIns_Inst_Sbox_6_M37 ;
    wire SubBytesIns_Inst_Sbox_6_M36 ;
    wire SubBytesIns_Inst_Sbox_6_M35 ;
    wire SubBytesIns_Inst_Sbox_6_M34 ;
    wire SubBytesIns_Inst_Sbox_6_M33 ;
    wire SubBytesIns_Inst_Sbox_6_M32 ;
    wire SubBytesIns_Inst_Sbox_6_M31 ;
    wire SubBytesIns_Inst_Sbox_6_M30 ;
    wire SubBytesIns_Inst_Sbox_6_M29 ;
    wire SubBytesIns_Inst_Sbox_6_M28 ;
    wire SubBytesIns_Inst_Sbox_6_M27 ;
    wire SubBytesIns_Inst_Sbox_6_M26 ;
    wire SubBytesIns_Inst_Sbox_6_M25 ;
    wire SubBytesIns_Inst_Sbox_6_M24 ;
    wire SubBytesIns_Inst_Sbox_6_M23 ;
    wire SubBytesIns_Inst_Sbox_6_M22 ;
    wire SubBytesIns_Inst_Sbox_6_M21 ;
    wire SubBytesIns_Inst_Sbox_6_M20 ;
    wire SubBytesIns_Inst_Sbox_6_M19 ;
    wire SubBytesIns_Inst_Sbox_6_M18 ;
    wire SubBytesIns_Inst_Sbox_6_M17 ;
    wire SubBytesIns_Inst_Sbox_6_M16 ;
    wire SubBytesIns_Inst_Sbox_6_M15 ;
    wire SubBytesIns_Inst_Sbox_6_M14 ;
    wire SubBytesIns_Inst_Sbox_6_M13 ;
    wire SubBytesIns_Inst_Sbox_6_M12 ;
    wire SubBytesIns_Inst_Sbox_6_M11 ;
    wire SubBytesIns_Inst_Sbox_6_M10 ;
    wire SubBytesIns_Inst_Sbox_6_M9 ;
    wire SubBytesIns_Inst_Sbox_6_M8 ;
    wire SubBytesIns_Inst_Sbox_6_M7 ;
    wire SubBytesIns_Inst_Sbox_6_M6 ;
    wire SubBytesIns_Inst_Sbox_6_M5 ;
    wire SubBytesIns_Inst_Sbox_6_M4 ;
    wire SubBytesIns_Inst_Sbox_6_M3 ;
    wire SubBytesIns_Inst_Sbox_6_M2 ;
    wire SubBytesIns_Inst_Sbox_6_M1 ;
    wire SubBytesIns_Inst_Sbox_6_T27 ;
    wire SubBytesIns_Inst_Sbox_6_T26 ;
    wire SubBytesIns_Inst_Sbox_6_T25 ;
    wire SubBytesIns_Inst_Sbox_6_T24 ;
    wire SubBytesIns_Inst_Sbox_6_T23 ;
    wire SubBytesIns_Inst_Sbox_6_T22 ;
    wire SubBytesIns_Inst_Sbox_6_T21 ;
    wire SubBytesIns_Inst_Sbox_6_T20 ;
    wire SubBytesIns_Inst_Sbox_6_T19 ;
    wire SubBytesIns_Inst_Sbox_6_T18 ;
    wire SubBytesIns_Inst_Sbox_6_T17 ;
    wire SubBytesIns_Inst_Sbox_6_T16 ;
    wire SubBytesIns_Inst_Sbox_6_T15 ;
    wire SubBytesIns_Inst_Sbox_6_T14 ;
    wire SubBytesIns_Inst_Sbox_6_T13 ;
    wire SubBytesIns_Inst_Sbox_6_T12 ;
    wire SubBytesIns_Inst_Sbox_6_T11 ;
    wire SubBytesIns_Inst_Sbox_6_T10 ;
    wire SubBytesIns_Inst_Sbox_6_T9 ;
    wire SubBytesIns_Inst_Sbox_6_T8 ;
    wire SubBytesIns_Inst_Sbox_6_T7 ;
    wire SubBytesIns_Inst_Sbox_6_T6 ;
    wire SubBytesIns_Inst_Sbox_6_T5 ;
    wire SubBytesIns_Inst_Sbox_6_T4 ;
    wire SubBytesIns_Inst_Sbox_6_T3 ;
    wire SubBytesIns_Inst_Sbox_6_T2 ;
    wire SubBytesIns_Inst_Sbox_6_T1 ;
    wire SubBytesIns_Inst_Sbox_7_L29 ;
    wire SubBytesIns_Inst_Sbox_7_L28 ;
    wire SubBytesIns_Inst_Sbox_7_L27 ;
    wire SubBytesIns_Inst_Sbox_7_L26 ;
    wire SubBytesIns_Inst_Sbox_7_L25 ;
    wire SubBytesIns_Inst_Sbox_7_L24 ;
    wire SubBytesIns_Inst_Sbox_7_L23 ;
    wire SubBytesIns_Inst_Sbox_7_L22 ;
    wire SubBytesIns_Inst_Sbox_7_L21 ;
    wire SubBytesIns_Inst_Sbox_7_L20 ;
    wire SubBytesIns_Inst_Sbox_7_L19 ;
    wire SubBytesIns_Inst_Sbox_7_L18 ;
    wire SubBytesIns_Inst_Sbox_7_L17 ;
    wire SubBytesIns_Inst_Sbox_7_L16 ;
    wire SubBytesIns_Inst_Sbox_7_L15 ;
    wire SubBytesIns_Inst_Sbox_7_L14 ;
    wire SubBytesIns_Inst_Sbox_7_L13 ;
    wire SubBytesIns_Inst_Sbox_7_L12 ;
    wire SubBytesIns_Inst_Sbox_7_L11 ;
    wire SubBytesIns_Inst_Sbox_7_L10 ;
    wire SubBytesIns_Inst_Sbox_7_L9 ;
    wire SubBytesIns_Inst_Sbox_7_L8 ;
    wire SubBytesIns_Inst_Sbox_7_L7 ;
    wire SubBytesIns_Inst_Sbox_7_L6 ;
    wire SubBytesIns_Inst_Sbox_7_L5 ;
    wire SubBytesIns_Inst_Sbox_7_L4 ;
    wire SubBytesIns_Inst_Sbox_7_L3 ;
    wire SubBytesIns_Inst_Sbox_7_L2 ;
    wire SubBytesIns_Inst_Sbox_7_L1 ;
    wire SubBytesIns_Inst_Sbox_7_L0 ;
    wire SubBytesIns_Inst_Sbox_7_M63 ;
    wire SubBytesIns_Inst_Sbox_7_M62 ;
    wire SubBytesIns_Inst_Sbox_7_M61 ;
    wire SubBytesIns_Inst_Sbox_7_M60 ;
    wire SubBytesIns_Inst_Sbox_7_M59 ;
    wire SubBytesIns_Inst_Sbox_7_M58 ;
    wire SubBytesIns_Inst_Sbox_7_M57 ;
    wire SubBytesIns_Inst_Sbox_7_M56 ;
    wire SubBytesIns_Inst_Sbox_7_M55 ;
    wire SubBytesIns_Inst_Sbox_7_M54 ;
    wire SubBytesIns_Inst_Sbox_7_M53 ;
    wire SubBytesIns_Inst_Sbox_7_M52 ;
    wire SubBytesIns_Inst_Sbox_7_M51 ;
    wire SubBytesIns_Inst_Sbox_7_M50 ;
    wire SubBytesIns_Inst_Sbox_7_M49 ;
    wire SubBytesIns_Inst_Sbox_7_M48 ;
    wire SubBytesIns_Inst_Sbox_7_M47 ;
    wire SubBytesIns_Inst_Sbox_7_M46 ;
    wire SubBytesIns_Inst_Sbox_7_M45 ;
    wire SubBytesIns_Inst_Sbox_7_M44 ;
    wire SubBytesIns_Inst_Sbox_7_M43 ;
    wire SubBytesIns_Inst_Sbox_7_M42 ;
    wire SubBytesIns_Inst_Sbox_7_M41 ;
    wire SubBytesIns_Inst_Sbox_7_M40 ;
    wire SubBytesIns_Inst_Sbox_7_M39 ;
    wire SubBytesIns_Inst_Sbox_7_M38 ;
    wire SubBytesIns_Inst_Sbox_7_M37 ;
    wire SubBytesIns_Inst_Sbox_7_M36 ;
    wire SubBytesIns_Inst_Sbox_7_M35 ;
    wire SubBytesIns_Inst_Sbox_7_M34 ;
    wire SubBytesIns_Inst_Sbox_7_M33 ;
    wire SubBytesIns_Inst_Sbox_7_M32 ;
    wire SubBytesIns_Inst_Sbox_7_M31 ;
    wire SubBytesIns_Inst_Sbox_7_M30 ;
    wire SubBytesIns_Inst_Sbox_7_M29 ;
    wire SubBytesIns_Inst_Sbox_7_M28 ;
    wire SubBytesIns_Inst_Sbox_7_M27 ;
    wire SubBytesIns_Inst_Sbox_7_M26 ;
    wire SubBytesIns_Inst_Sbox_7_M25 ;
    wire SubBytesIns_Inst_Sbox_7_M24 ;
    wire SubBytesIns_Inst_Sbox_7_M23 ;
    wire SubBytesIns_Inst_Sbox_7_M22 ;
    wire SubBytesIns_Inst_Sbox_7_M21 ;
    wire SubBytesIns_Inst_Sbox_7_M20 ;
    wire SubBytesIns_Inst_Sbox_7_M19 ;
    wire SubBytesIns_Inst_Sbox_7_M18 ;
    wire SubBytesIns_Inst_Sbox_7_M17 ;
    wire SubBytesIns_Inst_Sbox_7_M16 ;
    wire SubBytesIns_Inst_Sbox_7_M15 ;
    wire SubBytesIns_Inst_Sbox_7_M14 ;
    wire SubBytesIns_Inst_Sbox_7_M13 ;
    wire SubBytesIns_Inst_Sbox_7_M12 ;
    wire SubBytesIns_Inst_Sbox_7_M11 ;
    wire SubBytesIns_Inst_Sbox_7_M10 ;
    wire SubBytesIns_Inst_Sbox_7_M9 ;
    wire SubBytesIns_Inst_Sbox_7_M8 ;
    wire SubBytesIns_Inst_Sbox_7_M7 ;
    wire SubBytesIns_Inst_Sbox_7_M6 ;
    wire SubBytesIns_Inst_Sbox_7_M5 ;
    wire SubBytesIns_Inst_Sbox_7_M4 ;
    wire SubBytesIns_Inst_Sbox_7_M3 ;
    wire SubBytesIns_Inst_Sbox_7_M2 ;
    wire SubBytesIns_Inst_Sbox_7_M1 ;
    wire SubBytesIns_Inst_Sbox_7_T27 ;
    wire SubBytesIns_Inst_Sbox_7_T26 ;
    wire SubBytesIns_Inst_Sbox_7_T25 ;
    wire SubBytesIns_Inst_Sbox_7_T24 ;
    wire SubBytesIns_Inst_Sbox_7_T23 ;
    wire SubBytesIns_Inst_Sbox_7_T22 ;
    wire SubBytesIns_Inst_Sbox_7_T21 ;
    wire SubBytesIns_Inst_Sbox_7_T20 ;
    wire SubBytesIns_Inst_Sbox_7_T19 ;
    wire SubBytesIns_Inst_Sbox_7_T18 ;
    wire SubBytesIns_Inst_Sbox_7_T17 ;
    wire SubBytesIns_Inst_Sbox_7_T16 ;
    wire SubBytesIns_Inst_Sbox_7_T15 ;
    wire SubBytesIns_Inst_Sbox_7_T14 ;
    wire SubBytesIns_Inst_Sbox_7_T13 ;
    wire SubBytesIns_Inst_Sbox_7_T12 ;
    wire SubBytesIns_Inst_Sbox_7_T11 ;
    wire SubBytesIns_Inst_Sbox_7_T10 ;
    wire SubBytesIns_Inst_Sbox_7_T9 ;
    wire SubBytesIns_Inst_Sbox_7_T8 ;
    wire SubBytesIns_Inst_Sbox_7_T7 ;
    wire SubBytesIns_Inst_Sbox_7_T6 ;
    wire SubBytesIns_Inst_Sbox_7_T5 ;
    wire SubBytesIns_Inst_Sbox_7_T4 ;
    wire SubBytesIns_Inst_Sbox_7_T3 ;
    wire SubBytesIns_Inst_Sbox_7_T2 ;
    wire SubBytesIns_Inst_Sbox_7_T1 ;
    wire SubBytesIns_Inst_Sbox_8_L29 ;
    wire SubBytesIns_Inst_Sbox_8_L28 ;
    wire SubBytesIns_Inst_Sbox_8_L27 ;
    wire SubBytesIns_Inst_Sbox_8_L26 ;
    wire SubBytesIns_Inst_Sbox_8_L25 ;
    wire SubBytesIns_Inst_Sbox_8_L24 ;
    wire SubBytesIns_Inst_Sbox_8_L23 ;
    wire SubBytesIns_Inst_Sbox_8_L22 ;
    wire SubBytesIns_Inst_Sbox_8_L21 ;
    wire SubBytesIns_Inst_Sbox_8_L20 ;
    wire SubBytesIns_Inst_Sbox_8_L19 ;
    wire SubBytesIns_Inst_Sbox_8_L18 ;
    wire SubBytesIns_Inst_Sbox_8_L17 ;
    wire SubBytesIns_Inst_Sbox_8_L16 ;
    wire SubBytesIns_Inst_Sbox_8_L15 ;
    wire SubBytesIns_Inst_Sbox_8_L14 ;
    wire SubBytesIns_Inst_Sbox_8_L13 ;
    wire SubBytesIns_Inst_Sbox_8_L12 ;
    wire SubBytesIns_Inst_Sbox_8_L11 ;
    wire SubBytesIns_Inst_Sbox_8_L10 ;
    wire SubBytesIns_Inst_Sbox_8_L9 ;
    wire SubBytesIns_Inst_Sbox_8_L8 ;
    wire SubBytesIns_Inst_Sbox_8_L7 ;
    wire SubBytesIns_Inst_Sbox_8_L6 ;
    wire SubBytesIns_Inst_Sbox_8_L5 ;
    wire SubBytesIns_Inst_Sbox_8_L4 ;
    wire SubBytesIns_Inst_Sbox_8_L3 ;
    wire SubBytesIns_Inst_Sbox_8_L2 ;
    wire SubBytesIns_Inst_Sbox_8_L1 ;
    wire SubBytesIns_Inst_Sbox_8_L0 ;
    wire SubBytesIns_Inst_Sbox_8_M63 ;
    wire SubBytesIns_Inst_Sbox_8_M62 ;
    wire SubBytesIns_Inst_Sbox_8_M61 ;
    wire SubBytesIns_Inst_Sbox_8_M60 ;
    wire SubBytesIns_Inst_Sbox_8_M59 ;
    wire SubBytesIns_Inst_Sbox_8_M58 ;
    wire SubBytesIns_Inst_Sbox_8_M57 ;
    wire SubBytesIns_Inst_Sbox_8_M56 ;
    wire SubBytesIns_Inst_Sbox_8_M55 ;
    wire SubBytesIns_Inst_Sbox_8_M54 ;
    wire SubBytesIns_Inst_Sbox_8_M53 ;
    wire SubBytesIns_Inst_Sbox_8_M52 ;
    wire SubBytesIns_Inst_Sbox_8_M51 ;
    wire SubBytesIns_Inst_Sbox_8_M50 ;
    wire SubBytesIns_Inst_Sbox_8_M49 ;
    wire SubBytesIns_Inst_Sbox_8_M48 ;
    wire SubBytesIns_Inst_Sbox_8_M47 ;
    wire SubBytesIns_Inst_Sbox_8_M46 ;
    wire SubBytesIns_Inst_Sbox_8_M45 ;
    wire SubBytesIns_Inst_Sbox_8_M44 ;
    wire SubBytesIns_Inst_Sbox_8_M43 ;
    wire SubBytesIns_Inst_Sbox_8_M42 ;
    wire SubBytesIns_Inst_Sbox_8_M41 ;
    wire SubBytesIns_Inst_Sbox_8_M40 ;
    wire SubBytesIns_Inst_Sbox_8_M39 ;
    wire SubBytesIns_Inst_Sbox_8_M38 ;
    wire SubBytesIns_Inst_Sbox_8_M37 ;
    wire SubBytesIns_Inst_Sbox_8_M36 ;
    wire SubBytesIns_Inst_Sbox_8_M35 ;
    wire SubBytesIns_Inst_Sbox_8_M34 ;
    wire SubBytesIns_Inst_Sbox_8_M33 ;
    wire SubBytesIns_Inst_Sbox_8_M32 ;
    wire SubBytesIns_Inst_Sbox_8_M31 ;
    wire SubBytesIns_Inst_Sbox_8_M30 ;
    wire SubBytesIns_Inst_Sbox_8_M29 ;
    wire SubBytesIns_Inst_Sbox_8_M28 ;
    wire SubBytesIns_Inst_Sbox_8_M27 ;
    wire SubBytesIns_Inst_Sbox_8_M26 ;
    wire SubBytesIns_Inst_Sbox_8_M25 ;
    wire SubBytesIns_Inst_Sbox_8_M24 ;
    wire SubBytesIns_Inst_Sbox_8_M23 ;
    wire SubBytesIns_Inst_Sbox_8_M22 ;
    wire SubBytesIns_Inst_Sbox_8_M21 ;
    wire SubBytesIns_Inst_Sbox_8_M20 ;
    wire SubBytesIns_Inst_Sbox_8_M19 ;
    wire SubBytesIns_Inst_Sbox_8_M18 ;
    wire SubBytesIns_Inst_Sbox_8_M17 ;
    wire SubBytesIns_Inst_Sbox_8_M16 ;
    wire SubBytesIns_Inst_Sbox_8_M15 ;
    wire SubBytesIns_Inst_Sbox_8_M14 ;
    wire SubBytesIns_Inst_Sbox_8_M13 ;
    wire SubBytesIns_Inst_Sbox_8_M12 ;
    wire SubBytesIns_Inst_Sbox_8_M11 ;
    wire SubBytesIns_Inst_Sbox_8_M10 ;
    wire SubBytesIns_Inst_Sbox_8_M9 ;
    wire SubBytesIns_Inst_Sbox_8_M8 ;
    wire SubBytesIns_Inst_Sbox_8_M7 ;
    wire SubBytesIns_Inst_Sbox_8_M6 ;
    wire SubBytesIns_Inst_Sbox_8_M5 ;
    wire SubBytesIns_Inst_Sbox_8_M4 ;
    wire SubBytesIns_Inst_Sbox_8_M3 ;
    wire SubBytesIns_Inst_Sbox_8_M2 ;
    wire SubBytesIns_Inst_Sbox_8_M1 ;
    wire SubBytesIns_Inst_Sbox_8_T27 ;
    wire SubBytesIns_Inst_Sbox_8_T26 ;
    wire SubBytesIns_Inst_Sbox_8_T25 ;
    wire SubBytesIns_Inst_Sbox_8_T24 ;
    wire SubBytesIns_Inst_Sbox_8_T23 ;
    wire SubBytesIns_Inst_Sbox_8_T22 ;
    wire SubBytesIns_Inst_Sbox_8_T21 ;
    wire SubBytesIns_Inst_Sbox_8_T20 ;
    wire SubBytesIns_Inst_Sbox_8_T19 ;
    wire SubBytesIns_Inst_Sbox_8_T18 ;
    wire SubBytesIns_Inst_Sbox_8_T17 ;
    wire SubBytesIns_Inst_Sbox_8_T16 ;
    wire SubBytesIns_Inst_Sbox_8_T15 ;
    wire SubBytesIns_Inst_Sbox_8_T14 ;
    wire SubBytesIns_Inst_Sbox_8_T13 ;
    wire SubBytesIns_Inst_Sbox_8_T12 ;
    wire SubBytesIns_Inst_Sbox_8_T11 ;
    wire SubBytesIns_Inst_Sbox_8_T10 ;
    wire SubBytesIns_Inst_Sbox_8_T9 ;
    wire SubBytesIns_Inst_Sbox_8_T8 ;
    wire SubBytesIns_Inst_Sbox_8_T7 ;
    wire SubBytesIns_Inst_Sbox_8_T6 ;
    wire SubBytesIns_Inst_Sbox_8_T5 ;
    wire SubBytesIns_Inst_Sbox_8_T4 ;
    wire SubBytesIns_Inst_Sbox_8_T3 ;
    wire SubBytesIns_Inst_Sbox_8_T2 ;
    wire SubBytesIns_Inst_Sbox_8_T1 ;
    wire SubBytesIns_Inst_Sbox_9_L29 ;
    wire SubBytesIns_Inst_Sbox_9_L28 ;
    wire SubBytesIns_Inst_Sbox_9_L27 ;
    wire SubBytesIns_Inst_Sbox_9_L26 ;
    wire SubBytesIns_Inst_Sbox_9_L25 ;
    wire SubBytesIns_Inst_Sbox_9_L24 ;
    wire SubBytesIns_Inst_Sbox_9_L23 ;
    wire SubBytesIns_Inst_Sbox_9_L22 ;
    wire SubBytesIns_Inst_Sbox_9_L21 ;
    wire SubBytesIns_Inst_Sbox_9_L20 ;
    wire SubBytesIns_Inst_Sbox_9_L19 ;
    wire SubBytesIns_Inst_Sbox_9_L18 ;
    wire SubBytesIns_Inst_Sbox_9_L17 ;
    wire SubBytesIns_Inst_Sbox_9_L16 ;
    wire SubBytesIns_Inst_Sbox_9_L15 ;
    wire SubBytesIns_Inst_Sbox_9_L14 ;
    wire SubBytesIns_Inst_Sbox_9_L13 ;
    wire SubBytesIns_Inst_Sbox_9_L12 ;
    wire SubBytesIns_Inst_Sbox_9_L11 ;
    wire SubBytesIns_Inst_Sbox_9_L10 ;
    wire SubBytesIns_Inst_Sbox_9_L9 ;
    wire SubBytesIns_Inst_Sbox_9_L8 ;
    wire SubBytesIns_Inst_Sbox_9_L7 ;
    wire SubBytesIns_Inst_Sbox_9_L6 ;
    wire SubBytesIns_Inst_Sbox_9_L5 ;
    wire SubBytesIns_Inst_Sbox_9_L4 ;
    wire SubBytesIns_Inst_Sbox_9_L3 ;
    wire SubBytesIns_Inst_Sbox_9_L2 ;
    wire SubBytesIns_Inst_Sbox_9_L1 ;
    wire SubBytesIns_Inst_Sbox_9_L0 ;
    wire SubBytesIns_Inst_Sbox_9_M63 ;
    wire SubBytesIns_Inst_Sbox_9_M62 ;
    wire SubBytesIns_Inst_Sbox_9_M61 ;
    wire SubBytesIns_Inst_Sbox_9_M60 ;
    wire SubBytesIns_Inst_Sbox_9_M59 ;
    wire SubBytesIns_Inst_Sbox_9_M58 ;
    wire SubBytesIns_Inst_Sbox_9_M57 ;
    wire SubBytesIns_Inst_Sbox_9_M56 ;
    wire SubBytesIns_Inst_Sbox_9_M55 ;
    wire SubBytesIns_Inst_Sbox_9_M54 ;
    wire SubBytesIns_Inst_Sbox_9_M53 ;
    wire SubBytesIns_Inst_Sbox_9_M52 ;
    wire SubBytesIns_Inst_Sbox_9_M51 ;
    wire SubBytesIns_Inst_Sbox_9_M50 ;
    wire SubBytesIns_Inst_Sbox_9_M49 ;
    wire SubBytesIns_Inst_Sbox_9_M48 ;
    wire SubBytesIns_Inst_Sbox_9_M47 ;
    wire SubBytesIns_Inst_Sbox_9_M46 ;
    wire SubBytesIns_Inst_Sbox_9_M45 ;
    wire SubBytesIns_Inst_Sbox_9_M44 ;
    wire SubBytesIns_Inst_Sbox_9_M43 ;
    wire SubBytesIns_Inst_Sbox_9_M42 ;
    wire SubBytesIns_Inst_Sbox_9_M41 ;
    wire SubBytesIns_Inst_Sbox_9_M40 ;
    wire SubBytesIns_Inst_Sbox_9_M39 ;
    wire SubBytesIns_Inst_Sbox_9_M38 ;
    wire SubBytesIns_Inst_Sbox_9_M37 ;
    wire SubBytesIns_Inst_Sbox_9_M36 ;
    wire SubBytesIns_Inst_Sbox_9_M35 ;
    wire SubBytesIns_Inst_Sbox_9_M34 ;
    wire SubBytesIns_Inst_Sbox_9_M33 ;
    wire SubBytesIns_Inst_Sbox_9_M32 ;
    wire SubBytesIns_Inst_Sbox_9_M31 ;
    wire SubBytesIns_Inst_Sbox_9_M30 ;
    wire SubBytesIns_Inst_Sbox_9_M29 ;
    wire SubBytesIns_Inst_Sbox_9_M28 ;
    wire SubBytesIns_Inst_Sbox_9_M27 ;
    wire SubBytesIns_Inst_Sbox_9_M26 ;
    wire SubBytesIns_Inst_Sbox_9_M25 ;
    wire SubBytesIns_Inst_Sbox_9_M24 ;
    wire SubBytesIns_Inst_Sbox_9_M23 ;
    wire SubBytesIns_Inst_Sbox_9_M22 ;
    wire SubBytesIns_Inst_Sbox_9_M21 ;
    wire SubBytesIns_Inst_Sbox_9_M20 ;
    wire SubBytesIns_Inst_Sbox_9_M19 ;
    wire SubBytesIns_Inst_Sbox_9_M18 ;
    wire SubBytesIns_Inst_Sbox_9_M17 ;
    wire SubBytesIns_Inst_Sbox_9_M16 ;
    wire SubBytesIns_Inst_Sbox_9_M15 ;
    wire SubBytesIns_Inst_Sbox_9_M14 ;
    wire SubBytesIns_Inst_Sbox_9_M13 ;
    wire SubBytesIns_Inst_Sbox_9_M12 ;
    wire SubBytesIns_Inst_Sbox_9_M11 ;
    wire SubBytesIns_Inst_Sbox_9_M10 ;
    wire SubBytesIns_Inst_Sbox_9_M9 ;
    wire SubBytesIns_Inst_Sbox_9_M8 ;
    wire SubBytesIns_Inst_Sbox_9_M7 ;
    wire SubBytesIns_Inst_Sbox_9_M6 ;
    wire SubBytesIns_Inst_Sbox_9_M5 ;
    wire SubBytesIns_Inst_Sbox_9_M4 ;
    wire SubBytesIns_Inst_Sbox_9_M3 ;
    wire SubBytesIns_Inst_Sbox_9_M2 ;
    wire SubBytesIns_Inst_Sbox_9_M1 ;
    wire SubBytesIns_Inst_Sbox_9_T27 ;
    wire SubBytesIns_Inst_Sbox_9_T26 ;
    wire SubBytesIns_Inst_Sbox_9_T25 ;
    wire SubBytesIns_Inst_Sbox_9_T24 ;
    wire SubBytesIns_Inst_Sbox_9_T23 ;
    wire SubBytesIns_Inst_Sbox_9_T22 ;
    wire SubBytesIns_Inst_Sbox_9_T21 ;
    wire SubBytesIns_Inst_Sbox_9_T20 ;
    wire SubBytesIns_Inst_Sbox_9_T19 ;
    wire SubBytesIns_Inst_Sbox_9_T18 ;
    wire SubBytesIns_Inst_Sbox_9_T17 ;
    wire SubBytesIns_Inst_Sbox_9_T16 ;
    wire SubBytesIns_Inst_Sbox_9_T15 ;
    wire SubBytesIns_Inst_Sbox_9_T14 ;
    wire SubBytesIns_Inst_Sbox_9_T13 ;
    wire SubBytesIns_Inst_Sbox_9_T12 ;
    wire SubBytesIns_Inst_Sbox_9_T11 ;
    wire SubBytesIns_Inst_Sbox_9_T10 ;
    wire SubBytesIns_Inst_Sbox_9_T9 ;
    wire SubBytesIns_Inst_Sbox_9_T8 ;
    wire SubBytesIns_Inst_Sbox_9_T7 ;
    wire SubBytesIns_Inst_Sbox_9_T6 ;
    wire SubBytesIns_Inst_Sbox_9_T5 ;
    wire SubBytesIns_Inst_Sbox_9_T4 ;
    wire SubBytesIns_Inst_Sbox_9_T3 ;
    wire SubBytesIns_Inst_Sbox_9_T2 ;
    wire SubBytesIns_Inst_Sbox_9_T1 ;
    wire SubBytesIns_Inst_Sbox_10_L29 ;
    wire SubBytesIns_Inst_Sbox_10_L28 ;
    wire SubBytesIns_Inst_Sbox_10_L27 ;
    wire SubBytesIns_Inst_Sbox_10_L26 ;
    wire SubBytesIns_Inst_Sbox_10_L25 ;
    wire SubBytesIns_Inst_Sbox_10_L24 ;
    wire SubBytesIns_Inst_Sbox_10_L23 ;
    wire SubBytesIns_Inst_Sbox_10_L22 ;
    wire SubBytesIns_Inst_Sbox_10_L21 ;
    wire SubBytesIns_Inst_Sbox_10_L20 ;
    wire SubBytesIns_Inst_Sbox_10_L19 ;
    wire SubBytesIns_Inst_Sbox_10_L18 ;
    wire SubBytesIns_Inst_Sbox_10_L17 ;
    wire SubBytesIns_Inst_Sbox_10_L16 ;
    wire SubBytesIns_Inst_Sbox_10_L15 ;
    wire SubBytesIns_Inst_Sbox_10_L14 ;
    wire SubBytesIns_Inst_Sbox_10_L13 ;
    wire SubBytesIns_Inst_Sbox_10_L12 ;
    wire SubBytesIns_Inst_Sbox_10_L11 ;
    wire SubBytesIns_Inst_Sbox_10_L10 ;
    wire SubBytesIns_Inst_Sbox_10_L9 ;
    wire SubBytesIns_Inst_Sbox_10_L8 ;
    wire SubBytesIns_Inst_Sbox_10_L7 ;
    wire SubBytesIns_Inst_Sbox_10_L6 ;
    wire SubBytesIns_Inst_Sbox_10_L5 ;
    wire SubBytesIns_Inst_Sbox_10_L4 ;
    wire SubBytesIns_Inst_Sbox_10_L3 ;
    wire SubBytesIns_Inst_Sbox_10_L2 ;
    wire SubBytesIns_Inst_Sbox_10_L1 ;
    wire SubBytesIns_Inst_Sbox_10_L0 ;
    wire SubBytesIns_Inst_Sbox_10_M63 ;
    wire SubBytesIns_Inst_Sbox_10_M62 ;
    wire SubBytesIns_Inst_Sbox_10_M61 ;
    wire SubBytesIns_Inst_Sbox_10_M60 ;
    wire SubBytesIns_Inst_Sbox_10_M59 ;
    wire SubBytesIns_Inst_Sbox_10_M58 ;
    wire SubBytesIns_Inst_Sbox_10_M57 ;
    wire SubBytesIns_Inst_Sbox_10_M56 ;
    wire SubBytesIns_Inst_Sbox_10_M55 ;
    wire SubBytesIns_Inst_Sbox_10_M54 ;
    wire SubBytesIns_Inst_Sbox_10_M53 ;
    wire SubBytesIns_Inst_Sbox_10_M52 ;
    wire SubBytesIns_Inst_Sbox_10_M51 ;
    wire SubBytesIns_Inst_Sbox_10_M50 ;
    wire SubBytesIns_Inst_Sbox_10_M49 ;
    wire SubBytesIns_Inst_Sbox_10_M48 ;
    wire SubBytesIns_Inst_Sbox_10_M47 ;
    wire SubBytesIns_Inst_Sbox_10_M46 ;
    wire SubBytesIns_Inst_Sbox_10_M45 ;
    wire SubBytesIns_Inst_Sbox_10_M44 ;
    wire SubBytesIns_Inst_Sbox_10_M43 ;
    wire SubBytesIns_Inst_Sbox_10_M42 ;
    wire SubBytesIns_Inst_Sbox_10_M41 ;
    wire SubBytesIns_Inst_Sbox_10_M40 ;
    wire SubBytesIns_Inst_Sbox_10_M39 ;
    wire SubBytesIns_Inst_Sbox_10_M38 ;
    wire SubBytesIns_Inst_Sbox_10_M37 ;
    wire SubBytesIns_Inst_Sbox_10_M36 ;
    wire SubBytesIns_Inst_Sbox_10_M35 ;
    wire SubBytesIns_Inst_Sbox_10_M34 ;
    wire SubBytesIns_Inst_Sbox_10_M33 ;
    wire SubBytesIns_Inst_Sbox_10_M32 ;
    wire SubBytesIns_Inst_Sbox_10_M31 ;
    wire SubBytesIns_Inst_Sbox_10_M30 ;
    wire SubBytesIns_Inst_Sbox_10_M29 ;
    wire SubBytesIns_Inst_Sbox_10_M28 ;
    wire SubBytesIns_Inst_Sbox_10_M27 ;
    wire SubBytesIns_Inst_Sbox_10_M26 ;
    wire SubBytesIns_Inst_Sbox_10_M25 ;
    wire SubBytesIns_Inst_Sbox_10_M24 ;
    wire SubBytesIns_Inst_Sbox_10_M23 ;
    wire SubBytesIns_Inst_Sbox_10_M22 ;
    wire SubBytesIns_Inst_Sbox_10_M21 ;
    wire SubBytesIns_Inst_Sbox_10_M20 ;
    wire SubBytesIns_Inst_Sbox_10_M19 ;
    wire SubBytesIns_Inst_Sbox_10_M18 ;
    wire SubBytesIns_Inst_Sbox_10_M17 ;
    wire SubBytesIns_Inst_Sbox_10_M16 ;
    wire SubBytesIns_Inst_Sbox_10_M15 ;
    wire SubBytesIns_Inst_Sbox_10_M14 ;
    wire SubBytesIns_Inst_Sbox_10_M13 ;
    wire SubBytesIns_Inst_Sbox_10_M12 ;
    wire SubBytesIns_Inst_Sbox_10_M11 ;
    wire SubBytesIns_Inst_Sbox_10_M10 ;
    wire SubBytesIns_Inst_Sbox_10_M9 ;
    wire SubBytesIns_Inst_Sbox_10_M8 ;
    wire SubBytesIns_Inst_Sbox_10_M7 ;
    wire SubBytesIns_Inst_Sbox_10_M6 ;
    wire SubBytesIns_Inst_Sbox_10_M5 ;
    wire SubBytesIns_Inst_Sbox_10_M4 ;
    wire SubBytesIns_Inst_Sbox_10_M3 ;
    wire SubBytesIns_Inst_Sbox_10_M2 ;
    wire SubBytesIns_Inst_Sbox_10_M1 ;
    wire SubBytesIns_Inst_Sbox_10_T27 ;
    wire SubBytesIns_Inst_Sbox_10_T26 ;
    wire SubBytesIns_Inst_Sbox_10_T25 ;
    wire SubBytesIns_Inst_Sbox_10_T24 ;
    wire SubBytesIns_Inst_Sbox_10_T23 ;
    wire SubBytesIns_Inst_Sbox_10_T22 ;
    wire SubBytesIns_Inst_Sbox_10_T21 ;
    wire SubBytesIns_Inst_Sbox_10_T20 ;
    wire SubBytesIns_Inst_Sbox_10_T19 ;
    wire SubBytesIns_Inst_Sbox_10_T18 ;
    wire SubBytesIns_Inst_Sbox_10_T17 ;
    wire SubBytesIns_Inst_Sbox_10_T16 ;
    wire SubBytesIns_Inst_Sbox_10_T15 ;
    wire SubBytesIns_Inst_Sbox_10_T14 ;
    wire SubBytesIns_Inst_Sbox_10_T13 ;
    wire SubBytesIns_Inst_Sbox_10_T12 ;
    wire SubBytesIns_Inst_Sbox_10_T11 ;
    wire SubBytesIns_Inst_Sbox_10_T10 ;
    wire SubBytesIns_Inst_Sbox_10_T9 ;
    wire SubBytesIns_Inst_Sbox_10_T8 ;
    wire SubBytesIns_Inst_Sbox_10_T7 ;
    wire SubBytesIns_Inst_Sbox_10_T6 ;
    wire SubBytesIns_Inst_Sbox_10_T5 ;
    wire SubBytesIns_Inst_Sbox_10_T4 ;
    wire SubBytesIns_Inst_Sbox_10_T3 ;
    wire SubBytesIns_Inst_Sbox_10_T2 ;
    wire SubBytesIns_Inst_Sbox_10_T1 ;
    wire SubBytesIns_Inst_Sbox_11_L29 ;
    wire SubBytesIns_Inst_Sbox_11_L28 ;
    wire SubBytesIns_Inst_Sbox_11_L27 ;
    wire SubBytesIns_Inst_Sbox_11_L26 ;
    wire SubBytesIns_Inst_Sbox_11_L25 ;
    wire SubBytesIns_Inst_Sbox_11_L24 ;
    wire SubBytesIns_Inst_Sbox_11_L23 ;
    wire SubBytesIns_Inst_Sbox_11_L22 ;
    wire SubBytesIns_Inst_Sbox_11_L21 ;
    wire SubBytesIns_Inst_Sbox_11_L20 ;
    wire SubBytesIns_Inst_Sbox_11_L19 ;
    wire SubBytesIns_Inst_Sbox_11_L18 ;
    wire SubBytesIns_Inst_Sbox_11_L17 ;
    wire SubBytesIns_Inst_Sbox_11_L16 ;
    wire SubBytesIns_Inst_Sbox_11_L15 ;
    wire SubBytesIns_Inst_Sbox_11_L14 ;
    wire SubBytesIns_Inst_Sbox_11_L13 ;
    wire SubBytesIns_Inst_Sbox_11_L12 ;
    wire SubBytesIns_Inst_Sbox_11_L11 ;
    wire SubBytesIns_Inst_Sbox_11_L10 ;
    wire SubBytesIns_Inst_Sbox_11_L9 ;
    wire SubBytesIns_Inst_Sbox_11_L8 ;
    wire SubBytesIns_Inst_Sbox_11_L7 ;
    wire SubBytesIns_Inst_Sbox_11_L6 ;
    wire SubBytesIns_Inst_Sbox_11_L5 ;
    wire SubBytesIns_Inst_Sbox_11_L4 ;
    wire SubBytesIns_Inst_Sbox_11_L3 ;
    wire SubBytesIns_Inst_Sbox_11_L2 ;
    wire SubBytesIns_Inst_Sbox_11_L1 ;
    wire SubBytesIns_Inst_Sbox_11_L0 ;
    wire SubBytesIns_Inst_Sbox_11_M63 ;
    wire SubBytesIns_Inst_Sbox_11_M62 ;
    wire SubBytesIns_Inst_Sbox_11_M61 ;
    wire SubBytesIns_Inst_Sbox_11_M60 ;
    wire SubBytesIns_Inst_Sbox_11_M59 ;
    wire SubBytesIns_Inst_Sbox_11_M58 ;
    wire SubBytesIns_Inst_Sbox_11_M57 ;
    wire SubBytesIns_Inst_Sbox_11_M56 ;
    wire SubBytesIns_Inst_Sbox_11_M55 ;
    wire SubBytesIns_Inst_Sbox_11_M54 ;
    wire SubBytesIns_Inst_Sbox_11_M53 ;
    wire SubBytesIns_Inst_Sbox_11_M52 ;
    wire SubBytesIns_Inst_Sbox_11_M51 ;
    wire SubBytesIns_Inst_Sbox_11_M50 ;
    wire SubBytesIns_Inst_Sbox_11_M49 ;
    wire SubBytesIns_Inst_Sbox_11_M48 ;
    wire SubBytesIns_Inst_Sbox_11_M47 ;
    wire SubBytesIns_Inst_Sbox_11_M46 ;
    wire SubBytesIns_Inst_Sbox_11_M45 ;
    wire SubBytesIns_Inst_Sbox_11_M44 ;
    wire SubBytesIns_Inst_Sbox_11_M43 ;
    wire SubBytesIns_Inst_Sbox_11_M42 ;
    wire SubBytesIns_Inst_Sbox_11_M41 ;
    wire SubBytesIns_Inst_Sbox_11_M40 ;
    wire SubBytesIns_Inst_Sbox_11_M39 ;
    wire SubBytesIns_Inst_Sbox_11_M38 ;
    wire SubBytesIns_Inst_Sbox_11_M37 ;
    wire SubBytesIns_Inst_Sbox_11_M36 ;
    wire SubBytesIns_Inst_Sbox_11_M35 ;
    wire SubBytesIns_Inst_Sbox_11_M34 ;
    wire SubBytesIns_Inst_Sbox_11_M33 ;
    wire SubBytesIns_Inst_Sbox_11_M32 ;
    wire SubBytesIns_Inst_Sbox_11_M31 ;
    wire SubBytesIns_Inst_Sbox_11_M30 ;
    wire SubBytesIns_Inst_Sbox_11_M29 ;
    wire SubBytesIns_Inst_Sbox_11_M28 ;
    wire SubBytesIns_Inst_Sbox_11_M27 ;
    wire SubBytesIns_Inst_Sbox_11_M26 ;
    wire SubBytesIns_Inst_Sbox_11_M25 ;
    wire SubBytesIns_Inst_Sbox_11_M24 ;
    wire SubBytesIns_Inst_Sbox_11_M23 ;
    wire SubBytesIns_Inst_Sbox_11_M22 ;
    wire SubBytesIns_Inst_Sbox_11_M21 ;
    wire SubBytesIns_Inst_Sbox_11_M20 ;
    wire SubBytesIns_Inst_Sbox_11_M19 ;
    wire SubBytesIns_Inst_Sbox_11_M18 ;
    wire SubBytesIns_Inst_Sbox_11_M17 ;
    wire SubBytesIns_Inst_Sbox_11_M16 ;
    wire SubBytesIns_Inst_Sbox_11_M15 ;
    wire SubBytesIns_Inst_Sbox_11_M14 ;
    wire SubBytesIns_Inst_Sbox_11_M13 ;
    wire SubBytesIns_Inst_Sbox_11_M12 ;
    wire SubBytesIns_Inst_Sbox_11_M11 ;
    wire SubBytesIns_Inst_Sbox_11_M10 ;
    wire SubBytesIns_Inst_Sbox_11_M9 ;
    wire SubBytesIns_Inst_Sbox_11_M8 ;
    wire SubBytesIns_Inst_Sbox_11_M7 ;
    wire SubBytesIns_Inst_Sbox_11_M6 ;
    wire SubBytesIns_Inst_Sbox_11_M5 ;
    wire SubBytesIns_Inst_Sbox_11_M4 ;
    wire SubBytesIns_Inst_Sbox_11_M3 ;
    wire SubBytesIns_Inst_Sbox_11_M2 ;
    wire SubBytesIns_Inst_Sbox_11_M1 ;
    wire SubBytesIns_Inst_Sbox_11_T27 ;
    wire SubBytesIns_Inst_Sbox_11_T26 ;
    wire SubBytesIns_Inst_Sbox_11_T25 ;
    wire SubBytesIns_Inst_Sbox_11_T24 ;
    wire SubBytesIns_Inst_Sbox_11_T23 ;
    wire SubBytesIns_Inst_Sbox_11_T22 ;
    wire SubBytesIns_Inst_Sbox_11_T21 ;
    wire SubBytesIns_Inst_Sbox_11_T20 ;
    wire SubBytesIns_Inst_Sbox_11_T19 ;
    wire SubBytesIns_Inst_Sbox_11_T18 ;
    wire SubBytesIns_Inst_Sbox_11_T17 ;
    wire SubBytesIns_Inst_Sbox_11_T16 ;
    wire SubBytesIns_Inst_Sbox_11_T15 ;
    wire SubBytesIns_Inst_Sbox_11_T14 ;
    wire SubBytesIns_Inst_Sbox_11_T13 ;
    wire SubBytesIns_Inst_Sbox_11_T12 ;
    wire SubBytesIns_Inst_Sbox_11_T11 ;
    wire SubBytesIns_Inst_Sbox_11_T10 ;
    wire SubBytesIns_Inst_Sbox_11_T9 ;
    wire SubBytesIns_Inst_Sbox_11_T8 ;
    wire SubBytesIns_Inst_Sbox_11_T7 ;
    wire SubBytesIns_Inst_Sbox_11_T6 ;
    wire SubBytesIns_Inst_Sbox_11_T5 ;
    wire SubBytesIns_Inst_Sbox_11_T4 ;
    wire SubBytesIns_Inst_Sbox_11_T3 ;
    wire SubBytesIns_Inst_Sbox_11_T2 ;
    wire SubBytesIns_Inst_Sbox_11_T1 ;
    wire SubBytesIns_Inst_Sbox_12_L29 ;
    wire SubBytesIns_Inst_Sbox_12_L28 ;
    wire SubBytesIns_Inst_Sbox_12_L27 ;
    wire SubBytesIns_Inst_Sbox_12_L26 ;
    wire SubBytesIns_Inst_Sbox_12_L25 ;
    wire SubBytesIns_Inst_Sbox_12_L24 ;
    wire SubBytesIns_Inst_Sbox_12_L23 ;
    wire SubBytesIns_Inst_Sbox_12_L22 ;
    wire SubBytesIns_Inst_Sbox_12_L21 ;
    wire SubBytesIns_Inst_Sbox_12_L20 ;
    wire SubBytesIns_Inst_Sbox_12_L19 ;
    wire SubBytesIns_Inst_Sbox_12_L18 ;
    wire SubBytesIns_Inst_Sbox_12_L17 ;
    wire SubBytesIns_Inst_Sbox_12_L16 ;
    wire SubBytesIns_Inst_Sbox_12_L15 ;
    wire SubBytesIns_Inst_Sbox_12_L14 ;
    wire SubBytesIns_Inst_Sbox_12_L13 ;
    wire SubBytesIns_Inst_Sbox_12_L12 ;
    wire SubBytesIns_Inst_Sbox_12_L11 ;
    wire SubBytesIns_Inst_Sbox_12_L10 ;
    wire SubBytesIns_Inst_Sbox_12_L9 ;
    wire SubBytesIns_Inst_Sbox_12_L8 ;
    wire SubBytesIns_Inst_Sbox_12_L7 ;
    wire SubBytesIns_Inst_Sbox_12_L6 ;
    wire SubBytesIns_Inst_Sbox_12_L5 ;
    wire SubBytesIns_Inst_Sbox_12_L4 ;
    wire SubBytesIns_Inst_Sbox_12_L3 ;
    wire SubBytesIns_Inst_Sbox_12_L2 ;
    wire SubBytesIns_Inst_Sbox_12_L1 ;
    wire SubBytesIns_Inst_Sbox_12_L0 ;
    wire SubBytesIns_Inst_Sbox_12_M63 ;
    wire SubBytesIns_Inst_Sbox_12_M62 ;
    wire SubBytesIns_Inst_Sbox_12_M61 ;
    wire SubBytesIns_Inst_Sbox_12_M60 ;
    wire SubBytesIns_Inst_Sbox_12_M59 ;
    wire SubBytesIns_Inst_Sbox_12_M58 ;
    wire SubBytesIns_Inst_Sbox_12_M57 ;
    wire SubBytesIns_Inst_Sbox_12_M56 ;
    wire SubBytesIns_Inst_Sbox_12_M55 ;
    wire SubBytesIns_Inst_Sbox_12_M54 ;
    wire SubBytesIns_Inst_Sbox_12_M53 ;
    wire SubBytesIns_Inst_Sbox_12_M52 ;
    wire SubBytesIns_Inst_Sbox_12_M51 ;
    wire SubBytesIns_Inst_Sbox_12_M50 ;
    wire SubBytesIns_Inst_Sbox_12_M49 ;
    wire SubBytesIns_Inst_Sbox_12_M48 ;
    wire SubBytesIns_Inst_Sbox_12_M47 ;
    wire SubBytesIns_Inst_Sbox_12_M46 ;
    wire SubBytesIns_Inst_Sbox_12_M45 ;
    wire SubBytesIns_Inst_Sbox_12_M44 ;
    wire SubBytesIns_Inst_Sbox_12_M43 ;
    wire SubBytesIns_Inst_Sbox_12_M42 ;
    wire SubBytesIns_Inst_Sbox_12_M41 ;
    wire SubBytesIns_Inst_Sbox_12_M40 ;
    wire SubBytesIns_Inst_Sbox_12_M39 ;
    wire SubBytesIns_Inst_Sbox_12_M38 ;
    wire SubBytesIns_Inst_Sbox_12_M37 ;
    wire SubBytesIns_Inst_Sbox_12_M36 ;
    wire SubBytesIns_Inst_Sbox_12_M35 ;
    wire SubBytesIns_Inst_Sbox_12_M34 ;
    wire SubBytesIns_Inst_Sbox_12_M33 ;
    wire SubBytesIns_Inst_Sbox_12_M32 ;
    wire SubBytesIns_Inst_Sbox_12_M31 ;
    wire SubBytesIns_Inst_Sbox_12_M30 ;
    wire SubBytesIns_Inst_Sbox_12_M29 ;
    wire SubBytesIns_Inst_Sbox_12_M28 ;
    wire SubBytesIns_Inst_Sbox_12_M27 ;
    wire SubBytesIns_Inst_Sbox_12_M26 ;
    wire SubBytesIns_Inst_Sbox_12_M25 ;
    wire SubBytesIns_Inst_Sbox_12_M24 ;
    wire SubBytesIns_Inst_Sbox_12_M23 ;
    wire SubBytesIns_Inst_Sbox_12_M22 ;
    wire SubBytesIns_Inst_Sbox_12_M21 ;
    wire SubBytesIns_Inst_Sbox_12_M20 ;
    wire SubBytesIns_Inst_Sbox_12_M19 ;
    wire SubBytesIns_Inst_Sbox_12_M18 ;
    wire SubBytesIns_Inst_Sbox_12_M17 ;
    wire SubBytesIns_Inst_Sbox_12_M16 ;
    wire SubBytesIns_Inst_Sbox_12_M15 ;
    wire SubBytesIns_Inst_Sbox_12_M14 ;
    wire SubBytesIns_Inst_Sbox_12_M13 ;
    wire SubBytesIns_Inst_Sbox_12_M12 ;
    wire SubBytesIns_Inst_Sbox_12_M11 ;
    wire SubBytesIns_Inst_Sbox_12_M10 ;
    wire SubBytesIns_Inst_Sbox_12_M9 ;
    wire SubBytesIns_Inst_Sbox_12_M8 ;
    wire SubBytesIns_Inst_Sbox_12_M7 ;
    wire SubBytesIns_Inst_Sbox_12_M6 ;
    wire SubBytesIns_Inst_Sbox_12_M5 ;
    wire SubBytesIns_Inst_Sbox_12_M4 ;
    wire SubBytesIns_Inst_Sbox_12_M3 ;
    wire SubBytesIns_Inst_Sbox_12_M2 ;
    wire SubBytesIns_Inst_Sbox_12_M1 ;
    wire SubBytesIns_Inst_Sbox_12_T27 ;
    wire SubBytesIns_Inst_Sbox_12_T26 ;
    wire SubBytesIns_Inst_Sbox_12_T25 ;
    wire SubBytesIns_Inst_Sbox_12_T24 ;
    wire SubBytesIns_Inst_Sbox_12_T23 ;
    wire SubBytesIns_Inst_Sbox_12_T22 ;
    wire SubBytesIns_Inst_Sbox_12_T21 ;
    wire SubBytesIns_Inst_Sbox_12_T20 ;
    wire SubBytesIns_Inst_Sbox_12_T19 ;
    wire SubBytesIns_Inst_Sbox_12_T18 ;
    wire SubBytesIns_Inst_Sbox_12_T17 ;
    wire SubBytesIns_Inst_Sbox_12_T16 ;
    wire SubBytesIns_Inst_Sbox_12_T15 ;
    wire SubBytesIns_Inst_Sbox_12_T14 ;
    wire SubBytesIns_Inst_Sbox_12_T13 ;
    wire SubBytesIns_Inst_Sbox_12_T12 ;
    wire SubBytesIns_Inst_Sbox_12_T11 ;
    wire SubBytesIns_Inst_Sbox_12_T10 ;
    wire SubBytesIns_Inst_Sbox_12_T9 ;
    wire SubBytesIns_Inst_Sbox_12_T8 ;
    wire SubBytesIns_Inst_Sbox_12_T7 ;
    wire SubBytesIns_Inst_Sbox_12_T6 ;
    wire SubBytesIns_Inst_Sbox_12_T5 ;
    wire SubBytesIns_Inst_Sbox_12_T4 ;
    wire SubBytesIns_Inst_Sbox_12_T3 ;
    wire SubBytesIns_Inst_Sbox_12_T2 ;
    wire SubBytesIns_Inst_Sbox_12_T1 ;
    wire SubBytesIns_Inst_Sbox_13_L29 ;
    wire SubBytesIns_Inst_Sbox_13_L28 ;
    wire SubBytesIns_Inst_Sbox_13_L27 ;
    wire SubBytesIns_Inst_Sbox_13_L26 ;
    wire SubBytesIns_Inst_Sbox_13_L25 ;
    wire SubBytesIns_Inst_Sbox_13_L24 ;
    wire SubBytesIns_Inst_Sbox_13_L23 ;
    wire SubBytesIns_Inst_Sbox_13_L22 ;
    wire SubBytesIns_Inst_Sbox_13_L21 ;
    wire SubBytesIns_Inst_Sbox_13_L20 ;
    wire SubBytesIns_Inst_Sbox_13_L19 ;
    wire SubBytesIns_Inst_Sbox_13_L18 ;
    wire SubBytesIns_Inst_Sbox_13_L17 ;
    wire SubBytesIns_Inst_Sbox_13_L16 ;
    wire SubBytesIns_Inst_Sbox_13_L15 ;
    wire SubBytesIns_Inst_Sbox_13_L14 ;
    wire SubBytesIns_Inst_Sbox_13_L13 ;
    wire SubBytesIns_Inst_Sbox_13_L12 ;
    wire SubBytesIns_Inst_Sbox_13_L11 ;
    wire SubBytesIns_Inst_Sbox_13_L10 ;
    wire SubBytesIns_Inst_Sbox_13_L9 ;
    wire SubBytesIns_Inst_Sbox_13_L8 ;
    wire SubBytesIns_Inst_Sbox_13_L7 ;
    wire SubBytesIns_Inst_Sbox_13_L6 ;
    wire SubBytesIns_Inst_Sbox_13_L5 ;
    wire SubBytesIns_Inst_Sbox_13_L4 ;
    wire SubBytesIns_Inst_Sbox_13_L3 ;
    wire SubBytesIns_Inst_Sbox_13_L2 ;
    wire SubBytesIns_Inst_Sbox_13_L1 ;
    wire SubBytesIns_Inst_Sbox_13_L0 ;
    wire SubBytesIns_Inst_Sbox_13_M63 ;
    wire SubBytesIns_Inst_Sbox_13_M62 ;
    wire SubBytesIns_Inst_Sbox_13_M61 ;
    wire SubBytesIns_Inst_Sbox_13_M60 ;
    wire SubBytesIns_Inst_Sbox_13_M59 ;
    wire SubBytesIns_Inst_Sbox_13_M58 ;
    wire SubBytesIns_Inst_Sbox_13_M57 ;
    wire SubBytesIns_Inst_Sbox_13_M56 ;
    wire SubBytesIns_Inst_Sbox_13_M55 ;
    wire SubBytesIns_Inst_Sbox_13_M54 ;
    wire SubBytesIns_Inst_Sbox_13_M53 ;
    wire SubBytesIns_Inst_Sbox_13_M52 ;
    wire SubBytesIns_Inst_Sbox_13_M51 ;
    wire SubBytesIns_Inst_Sbox_13_M50 ;
    wire SubBytesIns_Inst_Sbox_13_M49 ;
    wire SubBytesIns_Inst_Sbox_13_M48 ;
    wire SubBytesIns_Inst_Sbox_13_M47 ;
    wire SubBytesIns_Inst_Sbox_13_M46 ;
    wire SubBytesIns_Inst_Sbox_13_M45 ;
    wire SubBytesIns_Inst_Sbox_13_M44 ;
    wire SubBytesIns_Inst_Sbox_13_M43 ;
    wire SubBytesIns_Inst_Sbox_13_M42 ;
    wire SubBytesIns_Inst_Sbox_13_M41 ;
    wire SubBytesIns_Inst_Sbox_13_M40 ;
    wire SubBytesIns_Inst_Sbox_13_M39 ;
    wire SubBytesIns_Inst_Sbox_13_M38 ;
    wire SubBytesIns_Inst_Sbox_13_M37 ;
    wire SubBytesIns_Inst_Sbox_13_M36 ;
    wire SubBytesIns_Inst_Sbox_13_M35 ;
    wire SubBytesIns_Inst_Sbox_13_M34 ;
    wire SubBytesIns_Inst_Sbox_13_M33 ;
    wire SubBytesIns_Inst_Sbox_13_M32 ;
    wire SubBytesIns_Inst_Sbox_13_M31 ;
    wire SubBytesIns_Inst_Sbox_13_M30 ;
    wire SubBytesIns_Inst_Sbox_13_M29 ;
    wire SubBytesIns_Inst_Sbox_13_M28 ;
    wire SubBytesIns_Inst_Sbox_13_M27 ;
    wire SubBytesIns_Inst_Sbox_13_M26 ;
    wire SubBytesIns_Inst_Sbox_13_M25 ;
    wire SubBytesIns_Inst_Sbox_13_M24 ;
    wire SubBytesIns_Inst_Sbox_13_M23 ;
    wire SubBytesIns_Inst_Sbox_13_M22 ;
    wire SubBytesIns_Inst_Sbox_13_M21 ;
    wire SubBytesIns_Inst_Sbox_13_M20 ;
    wire SubBytesIns_Inst_Sbox_13_M19 ;
    wire SubBytesIns_Inst_Sbox_13_M18 ;
    wire SubBytesIns_Inst_Sbox_13_M17 ;
    wire SubBytesIns_Inst_Sbox_13_M16 ;
    wire SubBytesIns_Inst_Sbox_13_M15 ;
    wire SubBytesIns_Inst_Sbox_13_M14 ;
    wire SubBytesIns_Inst_Sbox_13_M13 ;
    wire SubBytesIns_Inst_Sbox_13_M12 ;
    wire SubBytesIns_Inst_Sbox_13_M11 ;
    wire SubBytesIns_Inst_Sbox_13_M10 ;
    wire SubBytesIns_Inst_Sbox_13_M9 ;
    wire SubBytesIns_Inst_Sbox_13_M8 ;
    wire SubBytesIns_Inst_Sbox_13_M7 ;
    wire SubBytesIns_Inst_Sbox_13_M6 ;
    wire SubBytesIns_Inst_Sbox_13_M5 ;
    wire SubBytesIns_Inst_Sbox_13_M4 ;
    wire SubBytesIns_Inst_Sbox_13_M3 ;
    wire SubBytesIns_Inst_Sbox_13_M2 ;
    wire SubBytesIns_Inst_Sbox_13_M1 ;
    wire SubBytesIns_Inst_Sbox_13_T27 ;
    wire SubBytesIns_Inst_Sbox_13_T26 ;
    wire SubBytesIns_Inst_Sbox_13_T25 ;
    wire SubBytesIns_Inst_Sbox_13_T24 ;
    wire SubBytesIns_Inst_Sbox_13_T23 ;
    wire SubBytesIns_Inst_Sbox_13_T22 ;
    wire SubBytesIns_Inst_Sbox_13_T21 ;
    wire SubBytesIns_Inst_Sbox_13_T20 ;
    wire SubBytesIns_Inst_Sbox_13_T19 ;
    wire SubBytesIns_Inst_Sbox_13_T18 ;
    wire SubBytesIns_Inst_Sbox_13_T17 ;
    wire SubBytesIns_Inst_Sbox_13_T16 ;
    wire SubBytesIns_Inst_Sbox_13_T15 ;
    wire SubBytesIns_Inst_Sbox_13_T14 ;
    wire SubBytesIns_Inst_Sbox_13_T13 ;
    wire SubBytesIns_Inst_Sbox_13_T12 ;
    wire SubBytesIns_Inst_Sbox_13_T11 ;
    wire SubBytesIns_Inst_Sbox_13_T10 ;
    wire SubBytesIns_Inst_Sbox_13_T9 ;
    wire SubBytesIns_Inst_Sbox_13_T8 ;
    wire SubBytesIns_Inst_Sbox_13_T7 ;
    wire SubBytesIns_Inst_Sbox_13_T6 ;
    wire SubBytesIns_Inst_Sbox_13_T5 ;
    wire SubBytesIns_Inst_Sbox_13_T4 ;
    wire SubBytesIns_Inst_Sbox_13_T3 ;
    wire SubBytesIns_Inst_Sbox_13_T2 ;
    wire SubBytesIns_Inst_Sbox_13_T1 ;
    wire SubBytesIns_Inst_Sbox_14_L29 ;
    wire SubBytesIns_Inst_Sbox_14_L28 ;
    wire SubBytesIns_Inst_Sbox_14_L27 ;
    wire SubBytesIns_Inst_Sbox_14_L26 ;
    wire SubBytesIns_Inst_Sbox_14_L25 ;
    wire SubBytesIns_Inst_Sbox_14_L24 ;
    wire SubBytesIns_Inst_Sbox_14_L23 ;
    wire SubBytesIns_Inst_Sbox_14_L22 ;
    wire SubBytesIns_Inst_Sbox_14_L21 ;
    wire SubBytesIns_Inst_Sbox_14_L20 ;
    wire SubBytesIns_Inst_Sbox_14_L19 ;
    wire SubBytesIns_Inst_Sbox_14_L18 ;
    wire SubBytesIns_Inst_Sbox_14_L17 ;
    wire SubBytesIns_Inst_Sbox_14_L16 ;
    wire SubBytesIns_Inst_Sbox_14_L15 ;
    wire SubBytesIns_Inst_Sbox_14_L14 ;
    wire SubBytesIns_Inst_Sbox_14_L13 ;
    wire SubBytesIns_Inst_Sbox_14_L12 ;
    wire SubBytesIns_Inst_Sbox_14_L11 ;
    wire SubBytesIns_Inst_Sbox_14_L10 ;
    wire SubBytesIns_Inst_Sbox_14_L9 ;
    wire SubBytesIns_Inst_Sbox_14_L8 ;
    wire SubBytesIns_Inst_Sbox_14_L7 ;
    wire SubBytesIns_Inst_Sbox_14_L6 ;
    wire SubBytesIns_Inst_Sbox_14_L5 ;
    wire SubBytesIns_Inst_Sbox_14_L4 ;
    wire SubBytesIns_Inst_Sbox_14_L3 ;
    wire SubBytesIns_Inst_Sbox_14_L2 ;
    wire SubBytesIns_Inst_Sbox_14_L1 ;
    wire SubBytesIns_Inst_Sbox_14_L0 ;
    wire SubBytesIns_Inst_Sbox_14_M63 ;
    wire SubBytesIns_Inst_Sbox_14_M62 ;
    wire SubBytesIns_Inst_Sbox_14_M61 ;
    wire SubBytesIns_Inst_Sbox_14_M60 ;
    wire SubBytesIns_Inst_Sbox_14_M59 ;
    wire SubBytesIns_Inst_Sbox_14_M58 ;
    wire SubBytesIns_Inst_Sbox_14_M57 ;
    wire SubBytesIns_Inst_Sbox_14_M56 ;
    wire SubBytesIns_Inst_Sbox_14_M55 ;
    wire SubBytesIns_Inst_Sbox_14_M54 ;
    wire SubBytesIns_Inst_Sbox_14_M53 ;
    wire SubBytesIns_Inst_Sbox_14_M52 ;
    wire SubBytesIns_Inst_Sbox_14_M51 ;
    wire SubBytesIns_Inst_Sbox_14_M50 ;
    wire SubBytesIns_Inst_Sbox_14_M49 ;
    wire SubBytesIns_Inst_Sbox_14_M48 ;
    wire SubBytesIns_Inst_Sbox_14_M47 ;
    wire SubBytesIns_Inst_Sbox_14_M46 ;
    wire SubBytesIns_Inst_Sbox_14_M45 ;
    wire SubBytesIns_Inst_Sbox_14_M44 ;
    wire SubBytesIns_Inst_Sbox_14_M43 ;
    wire SubBytesIns_Inst_Sbox_14_M42 ;
    wire SubBytesIns_Inst_Sbox_14_M41 ;
    wire SubBytesIns_Inst_Sbox_14_M40 ;
    wire SubBytesIns_Inst_Sbox_14_M39 ;
    wire SubBytesIns_Inst_Sbox_14_M38 ;
    wire SubBytesIns_Inst_Sbox_14_M37 ;
    wire SubBytesIns_Inst_Sbox_14_M36 ;
    wire SubBytesIns_Inst_Sbox_14_M35 ;
    wire SubBytesIns_Inst_Sbox_14_M34 ;
    wire SubBytesIns_Inst_Sbox_14_M33 ;
    wire SubBytesIns_Inst_Sbox_14_M32 ;
    wire SubBytesIns_Inst_Sbox_14_M31 ;
    wire SubBytesIns_Inst_Sbox_14_M30 ;
    wire SubBytesIns_Inst_Sbox_14_M29 ;
    wire SubBytesIns_Inst_Sbox_14_M28 ;
    wire SubBytesIns_Inst_Sbox_14_M27 ;
    wire SubBytesIns_Inst_Sbox_14_M26 ;
    wire SubBytesIns_Inst_Sbox_14_M25 ;
    wire SubBytesIns_Inst_Sbox_14_M24 ;
    wire SubBytesIns_Inst_Sbox_14_M23 ;
    wire SubBytesIns_Inst_Sbox_14_M22 ;
    wire SubBytesIns_Inst_Sbox_14_M21 ;
    wire SubBytesIns_Inst_Sbox_14_M20 ;
    wire SubBytesIns_Inst_Sbox_14_M19 ;
    wire SubBytesIns_Inst_Sbox_14_M18 ;
    wire SubBytesIns_Inst_Sbox_14_M17 ;
    wire SubBytesIns_Inst_Sbox_14_M16 ;
    wire SubBytesIns_Inst_Sbox_14_M15 ;
    wire SubBytesIns_Inst_Sbox_14_M14 ;
    wire SubBytesIns_Inst_Sbox_14_M13 ;
    wire SubBytesIns_Inst_Sbox_14_M12 ;
    wire SubBytesIns_Inst_Sbox_14_M11 ;
    wire SubBytesIns_Inst_Sbox_14_M10 ;
    wire SubBytesIns_Inst_Sbox_14_M9 ;
    wire SubBytesIns_Inst_Sbox_14_M8 ;
    wire SubBytesIns_Inst_Sbox_14_M7 ;
    wire SubBytesIns_Inst_Sbox_14_M6 ;
    wire SubBytesIns_Inst_Sbox_14_M5 ;
    wire SubBytesIns_Inst_Sbox_14_M4 ;
    wire SubBytesIns_Inst_Sbox_14_M3 ;
    wire SubBytesIns_Inst_Sbox_14_M2 ;
    wire SubBytesIns_Inst_Sbox_14_M1 ;
    wire SubBytesIns_Inst_Sbox_14_T27 ;
    wire SubBytesIns_Inst_Sbox_14_T26 ;
    wire SubBytesIns_Inst_Sbox_14_T25 ;
    wire SubBytesIns_Inst_Sbox_14_T24 ;
    wire SubBytesIns_Inst_Sbox_14_T23 ;
    wire SubBytesIns_Inst_Sbox_14_T22 ;
    wire SubBytesIns_Inst_Sbox_14_T21 ;
    wire SubBytesIns_Inst_Sbox_14_T20 ;
    wire SubBytesIns_Inst_Sbox_14_T19 ;
    wire SubBytesIns_Inst_Sbox_14_T18 ;
    wire SubBytesIns_Inst_Sbox_14_T17 ;
    wire SubBytesIns_Inst_Sbox_14_T16 ;
    wire SubBytesIns_Inst_Sbox_14_T15 ;
    wire SubBytesIns_Inst_Sbox_14_T14 ;
    wire SubBytesIns_Inst_Sbox_14_T13 ;
    wire SubBytesIns_Inst_Sbox_14_T12 ;
    wire SubBytesIns_Inst_Sbox_14_T11 ;
    wire SubBytesIns_Inst_Sbox_14_T10 ;
    wire SubBytesIns_Inst_Sbox_14_T9 ;
    wire SubBytesIns_Inst_Sbox_14_T8 ;
    wire SubBytesIns_Inst_Sbox_14_T7 ;
    wire SubBytesIns_Inst_Sbox_14_T6 ;
    wire SubBytesIns_Inst_Sbox_14_T5 ;
    wire SubBytesIns_Inst_Sbox_14_T4 ;
    wire SubBytesIns_Inst_Sbox_14_T3 ;
    wire SubBytesIns_Inst_Sbox_14_T2 ;
    wire SubBytesIns_Inst_Sbox_14_T1 ;
    wire SubBytesIns_Inst_Sbox_15_L29 ;
    wire SubBytesIns_Inst_Sbox_15_L28 ;
    wire SubBytesIns_Inst_Sbox_15_L27 ;
    wire SubBytesIns_Inst_Sbox_15_L26 ;
    wire SubBytesIns_Inst_Sbox_15_L25 ;
    wire SubBytesIns_Inst_Sbox_15_L24 ;
    wire SubBytesIns_Inst_Sbox_15_L23 ;
    wire SubBytesIns_Inst_Sbox_15_L22 ;
    wire SubBytesIns_Inst_Sbox_15_L21 ;
    wire SubBytesIns_Inst_Sbox_15_L20 ;
    wire SubBytesIns_Inst_Sbox_15_L19 ;
    wire SubBytesIns_Inst_Sbox_15_L18 ;
    wire SubBytesIns_Inst_Sbox_15_L17 ;
    wire SubBytesIns_Inst_Sbox_15_L16 ;
    wire SubBytesIns_Inst_Sbox_15_L15 ;
    wire SubBytesIns_Inst_Sbox_15_L14 ;
    wire SubBytesIns_Inst_Sbox_15_L13 ;
    wire SubBytesIns_Inst_Sbox_15_L12 ;
    wire SubBytesIns_Inst_Sbox_15_L11 ;
    wire SubBytesIns_Inst_Sbox_15_L10 ;
    wire SubBytesIns_Inst_Sbox_15_L9 ;
    wire SubBytesIns_Inst_Sbox_15_L8 ;
    wire SubBytesIns_Inst_Sbox_15_L7 ;
    wire SubBytesIns_Inst_Sbox_15_L6 ;
    wire SubBytesIns_Inst_Sbox_15_L5 ;
    wire SubBytesIns_Inst_Sbox_15_L4 ;
    wire SubBytesIns_Inst_Sbox_15_L3 ;
    wire SubBytesIns_Inst_Sbox_15_L2 ;
    wire SubBytesIns_Inst_Sbox_15_L1 ;
    wire SubBytesIns_Inst_Sbox_15_L0 ;
    wire SubBytesIns_Inst_Sbox_15_M63 ;
    wire SubBytesIns_Inst_Sbox_15_M62 ;
    wire SubBytesIns_Inst_Sbox_15_M61 ;
    wire SubBytesIns_Inst_Sbox_15_M60 ;
    wire SubBytesIns_Inst_Sbox_15_M59 ;
    wire SubBytesIns_Inst_Sbox_15_M58 ;
    wire SubBytesIns_Inst_Sbox_15_M57 ;
    wire SubBytesIns_Inst_Sbox_15_M56 ;
    wire SubBytesIns_Inst_Sbox_15_M55 ;
    wire SubBytesIns_Inst_Sbox_15_M54 ;
    wire SubBytesIns_Inst_Sbox_15_M53 ;
    wire SubBytesIns_Inst_Sbox_15_M52 ;
    wire SubBytesIns_Inst_Sbox_15_M51 ;
    wire SubBytesIns_Inst_Sbox_15_M50 ;
    wire SubBytesIns_Inst_Sbox_15_M49 ;
    wire SubBytesIns_Inst_Sbox_15_M48 ;
    wire SubBytesIns_Inst_Sbox_15_M47 ;
    wire SubBytesIns_Inst_Sbox_15_M46 ;
    wire SubBytesIns_Inst_Sbox_15_M45 ;
    wire SubBytesIns_Inst_Sbox_15_M44 ;
    wire SubBytesIns_Inst_Sbox_15_M43 ;
    wire SubBytesIns_Inst_Sbox_15_M42 ;
    wire SubBytesIns_Inst_Sbox_15_M41 ;
    wire SubBytesIns_Inst_Sbox_15_M40 ;
    wire SubBytesIns_Inst_Sbox_15_M39 ;
    wire SubBytesIns_Inst_Sbox_15_M38 ;
    wire SubBytesIns_Inst_Sbox_15_M37 ;
    wire SubBytesIns_Inst_Sbox_15_M36 ;
    wire SubBytesIns_Inst_Sbox_15_M35 ;
    wire SubBytesIns_Inst_Sbox_15_M34 ;
    wire SubBytesIns_Inst_Sbox_15_M33 ;
    wire SubBytesIns_Inst_Sbox_15_M32 ;
    wire SubBytesIns_Inst_Sbox_15_M31 ;
    wire SubBytesIns_Inst_Sbox_15_M30 ;
    wire SubBytesIns_Inst_Sbox_15_M29 ;
    wire SubBytesIns_Inst_Sbox_15_M28 ;
    wire SubBytesIns_Inst_Sbox_15_M27 ;
    wire SubBytesIns_Inst_Sbox_15_M26 ;
    wire SubBytesIns_Inst_Sbox_15_M25 ;
    wire SubBytesIns_Inst_Sbox_15_M24 ;
    wire SubBytesIns_Inst_Sbox_15_M23 ;
    wire SubBytesIns_Inst_Sbox_15_M22 ;
    wire SubBytesIns_Inst_Sbox_15_M21 ;
    wire SubBytesIns_Inst_Sbox_15_M20 ;
    wire SubBytesIns_Inst_Sbox_15_M19 ;
    wire SubBytesIns_Inst_Sbox_15_M18 ;
    wire SubBytesIns_Inst_Sbox_15_M17 ;
    wire SubBytesIns_Inst_Sbox_15_M16 ;
    wire SubBytesIns_Inst_Sbox_15_M15 ;
    wire SubBytesIns_Inst_Sbox_15_M14 ;
    wire SubBytesIns_Inst_Sbox_15_M13 ;
    wire SubBytesIns_Inst_Sbox_15_M12 ;
    wire SubBytesIns_Inst_Sbox_15_M11 ;
    wire SubBytesIns_Inst_Sbox_15_M10 ;
    wire SubBytesIns_Inst_Sbox_15_M9 ;
    wire SubBytesIns_Inst_Sbox_15_M8 ;
    wire SubBytesIns_Inst_Sbox_15_M7 ;
    wire SubBytesIns_Inst_Sbox_15_M6 ;
    wire SubBytesIns_Inst_Sbox_15_M5 ;
    wire SubBytesIns_Inst_Sbox_15_M4 ;
    wire SubBytesIns_Inst_Sbox_15_M3 ;
    wire SubBytesIns_Inst_Sbox_15_M2 ;
    wire SubBytesIns_Inst_Sbox_15_M1 ;
    wire SubBytesIns_Inst_Sbox_15_T27 ;
    wire SubBytesIns_Inst_Sbox_15_T26 ;
    wire SubBytesIns_Inst_Sbox_15_T25 ;
    wire SubBytesIns_Inst_Sbox_15_T24 ;
    wire SubBytesIns_Inst_Sbox_15_T23 ;
    wire SubBytesIns_Inst_Sbox_15_T22 ;
    wire SubBytesIns_Inst_Sbox_15_T21 ;
    wire SubBytesIns_Inst_Sbox_15_T20 ;
    wire SubBytesIns_Inst_Sbox_15_T19 ;
    wire SubBytesIns_Inst_Sbox_15_T18 ;
    wire SubBytesIns_Inst_Sbox_15_T17 ;
    wire SubBytesIns_Inst_Sbox_15_T16 ;
    wire SubBytesIns_Inst_Sbox_15_T15 ;
    wire SubBytesIns_Inst_Sbox_15_T14 ;
    wire SubBytesIns_Inst_Sbox_15_T13 ;
    wire SubBytesIns_Inst_Sbox_15_T12 ;
    wire SubBytesIns_Inst_Sbox_15_T11 ;
    wire SubBytesIns_Inst_Sbox_15_T10 ;
    wire SubBytesIns_Inst_Sbox_15_T9 ;
    wire SubBytesIns_Inst_Sbox_15_T8 ;
    wire SubBytesIns_Inst_Sbox_15_T7 ;
    wire SubBytesIns_Inst_Sbox_15_T6 ;
    wire SubBytesIns_Inst_Sbox_15_T5 ;
    wire SubBytesIns_Inst_Sbox_15_T4 ;
    wire SubBytesIns_Inst_Sbox_15_T3 ;
    wire SubBytesIns_Inst_Sbox_15_T2 ;
    wire SubBytesIns_Inst_Sbox_15_T1 ;
    wire MixColumnsIns_MixOneColumnInst_0_n192 ;
    wire MixColumnsIns_MixOneColumnInst_0_n191 ;
    wire MixColumnsIns_MixOneColumnInst_0_n190 ;
    wire MixColumnsIns_MixOneColumnInst_0_n189 ;
    wire MixColumnsIns_MixOneColumnInst_0_n188 ;
    wire MixColumnsIns_MixOneColumnInst_0_n187 ;
    wire MixColumnsIns_MixOneColumnInst_0_n186 ;
    wire MixColumnsIns_MixOneColumnInst_0_n185 ;
    wire MixColumnsIns_MixOneColumnInst_0_n184 ;
    wire MixColumnsIns_MixOneColumnInst_0_n183 ;
    wire MixColumnsIns_MixOneColumnInst_0_n182 ;
    wire MixColumnsIns_MixOneColumnInst_0_n181 ;
    wire MixColumnsIns_MixOneColumnInst_0_n180 ;
    wire MixColumnsIns_MixOneColumnInst_0_n179 ;
    wire MixColumnsIns_MixOneColumnInst_0_n178 ;
    wire MixColumnsIns_MixOneColumnInst_0_n177 ;
    wire MixColumnsIns_MixOneColumnInst_0_n176 ;
    wire MixColumnsIns_MixOneColumnInst_0_n175 ;
    wire MixColumnsIns_MixOneColumnInst_0_n174 ;
    wire MixColumnsIns_MixOneColumnInst_0_n173 ;
    wire MixColumnsIns_MixOneColumnInst_0_n172 ;
    wire MixColumnsIns_MixOneColumnInst_0_n171 ;
    wire MixColumnsIns_MixOneColumnInst_0_n170 ;
    wire MixColumnsIns_MixOneColumnInst_0_n169 ;
    wire MixColumnsIns_MixOneColumnInst_0_n168 ;
    wire MixColumnsIns_MixOneColumnInst_0_n167 ;
    wire MixColumnsIns_MixOneColumnInst_0_n166 ;
    wire MixColumnsIns_MixOneColumnInst_0_n165 ;
    wire MixColumnsIns_MixOneColumnInst_0_n164 ;
    wire MixColumnsIns_MixOneColumnInst_0_n163 ;
    wire MixColumnsIns_MixOneColumnInst_0_n162 ;
    wire MixColumnsIns_MixOneColumnInst_0_n161 ;
    wire MixColumnsIns_MixOneColumnInst_0_n160 ;
    wire MixColumnsIns_MixOneColumnInst_0_n159 ;
    wire MixColumnsIns_MixOneColumnInst_0_n158 ;
    wire MixColumnsIns_MixOneColumnInst_0_n157 ;
    wire MixColumnsIns_MixOneColumnInst_0_n156 ;
    wire MixColumnsIns_MixOneColumnInst_0_n155 ;
    wire MixColumnsIns_MixOneColumnInst_0_n154 ;
    wire MixColumnsIns_MixOneColumnInst_0_n153 ;
    wire MixColumnsIns_MixOneColumnInst_0_n152 ;
    wire MixColumnsIns_MixOneColumnInst_0_n151 ;
    wire MixColumnsIns_MixOneColumnInst_0_n150 ;
    wire MixColumnsIns_MixOneColumnInst_0_n149 ;
    wire MixColumnsIns_MixOneColumnInst_0_n148 ;
    wire MixColumnsIns_MixOneColumnInst_0_n147 ;
    wire MixColumnsIns_MixOneColumnInst_0_n146 ;
    wire MixColumnsIns_MixOneColumnInst_0_n145 ;
    wire MixColumnsIns_MixOneColumnInst_0_n144 ;
    wire MixColumnsIns_MixOneColumnInst_0_n143 ;
    wire MixColumnsIns_MixOneColumnInst_0_n142 ;
    wire MixColumnsIns_MixOneColumnInst_0_n141 ;
    wire MixColumnsIns_MixOneColumnInst_0_n140 ;
    wire MixColumnsIns_MixOneColumnInst_0_n139 ;
    wire MixColumnsIns_MixOneColumnInst_0_n138 ;
    wire MixColumnsIns_MixOneColumnInst_0_n137 ;
    wire MixColumnsIns_MixOneColumnInst_0_n136 ;
    wire MixColumnsIns_MixOneColumnInst_0_n135 ;
    wire MixColumnsIns_MixOneColumnInst_0_n134 ;
    wire MixColumnsIns_MixOneColumnInst_0_n133 ;
    wire MixColumnsIns_MixOneColumnInst_0_n132 ;
    wire MixColumnsIns_MixOneColumnInst_0_n131 ;
    wire MixColumnsIns_MixOneColumnInst_0_n130 ;
    wire MixColumnsIns_MixOneColumnInst_0_n129 ;
    wire MixColumnsIns_MixOneColumnInst_1_n192 ;
    wire MixColumnsIns_MixOneColumnInst_1_n191 ;
    wire MixColumnsIns_MixOneColumnInst_1_n190 ;
    wire MixColumnsIns_MixOneColumnInst_1_n189 ;
    wire MixColumnsIns_MixOneColumnInst_1_n188 ;
    wire MixColumnsIns_MixOneColumnInst_1_n187 ;
    wire MixColumnsIns_MixOneColumnInst_1_n186 ;
    wire MixColumnsIns_MixOneColumnInst_1_n185 ;
    wire MixColumnsIns_MixOneColumnInst_1_n184 ;
    wire MixColumnsIns_MixOneColumnInst_1_n183 ;
    wire MixColumnsIns_MixOneColumnInst_1_n182 ;
    wire MixColumnsIns_MixOneColumnInst_1_n181 ;
    wire MixColumnsIns_MixOneColumnInst_1_n180 ;
    wire MixColumnsIns_MixOneColumnInst_1_n179 ;
    wire MixColumnsIns_MixOneColumnInst_1_n178 ;
    wire MixColumnsIns_MixOneColumnInst_1_n177 ;
    wire MixColumnsIns_MixOneColumnInst_1_n176 ;
    wire MixColumnsIns_MixOneColumnInst_1_n175 ;
    wire MixColumnsIns_MixOneColumnInst_1_n174 ;
    wire MixColumnsIns_MixOneColumnInst_1_n173 ;
    wire MixColumnsIns_MixOneColumnInst_1_n172 ;
    wire MixColumnsIns_MixOneColumnInst_1_n171 ;
    wire MixColumnsIns_MixOneColumnInst_1_n170 ;
    wire MixColumnsIns_MixOneColumnInst_1_n169 ;
    wire MixColumnsIns_MixOneColumnInst_1_n168 ;
    wire MixColumnsIns_MixOneColumnInst_1_n167 ;
    wire MixColumnsIns_MixOneColumnInst_1_n166 ;
    wire MixColumnsIns_MixOneColumnInst_1_n165 ;
    wire MixColumnsIns_MixOneColumnInst_1_n164 ;
    wire MixColumnsIns_MixOneColumnInst_1_n163 ;
    wire MixColumnsIns_MixOneColumnInst_1_n162 ;
    wire MixColumnsIns_MixOneColumnInst_1_n161 ;
    wire MixColumnsIns_MixOneColumnInst_1_n160 ;
    wire MixColumnsIns_MixOneColumnInst_1_n159 ;
    wire MixColumnsIns_MixOneColumnInst_1_n158 ;
    wire MixColumnsIns_MixOneColumnInst_1_n157 ;
    wire MixColumnsIns_MixOneColumnInst_1_n156 ;
    wire MixColumnsIns_MixOneColumnInst_1_n155 ;
    wire MixColumnsIns_MixOneColumnInst_1_n154 ;
    wire MixColumnsIns_MixOneColumnInst_1_n153 ;
    wire MixColumnsIns_MixOneColumnInst_1_n152 ;
    wire MixColumnsIns_MixOneColumnInst_1_n151 ;
    wire MixColumnsIns_MixOneColumnInst_1_n150 ;
    wire MixColumnsIns_MixOneColumnInst_1_n149 ;
    wire MixColumnsIns_MixOneColumnInst_1_n148 ;
    wire MixColumnsIns_MixOneColumnInst_1_n147 ;
    wire MixColumnsIns_MixOneColumnInst_1_n146 ;
    wire MixColumnsIns_MixOneColumnInst_1_n145 ;
    wire MixColumnsIns_MixOneColumnInst_1_n144 ;
    wire MixColumnsIns_MixOneColumnInst_1_n143 ;
    wire MixColumnsIns_MixOneColumnInst_1_n142 ;
    wire MixColumnsIns_MixOneColumnInst_1_n141 ;
    wire MixColumnsIns_MixOneColumnInst_1_n140 ;
    wire MixColumnsIns_MixOneColumnInst_1_n139 ;
    wire MixColumnsIns_MixOneColumnInst_1_n138 ;
    wire MixColumnsIns_MixOneColumnInst_1_n137 ;
    wire MixColumnsIns_MixOneColumnInst_1_n136 ;
    wire MixColumnsIns_MixOneColumnInst_1_n135 ;
    wire MixColumnsIns_MixOneColumnInst_1_n134 ;
    wire MixColumnsIns_MixOneColumnInst_1_n133 ;
    wire MixColumnsIns_MixOneColumnInst_1_n132 ;
    wire MixColumnsIns_MixOneColumnInst_1_n131 ;
    wire MixColumnsIns_MixOneColumnInst_1_n130 ;
    wire MixColumnsIns_MixOneColumnInst_1_n129 ;
    wire MixColumnsIns_MixOneColumnInst_2_n192 ;
    wire MixColumnsIns_MixOneColumnInst_2_n191 ;
    wire MixColumnsIns_MixOneColumnInst_2_n190 ;
    wire MixColumnsIns_MixOneColumnInst_2_n189 ;
    wire MixColumnsIns_MixOneColumnInst_2_n188 ;
    wire MixColumnsIns_MixOneColumnInst_2_n187 ;
    wire MixColumnsIns_MixOneColumnInst_2_n186 ;
    wire MixColumnsIns_MixOneColumnInst_2_n185 ;
    wire MixColumnsIns_MixOneColumnInst_2_n184 ;
    wire MixColumnsIns_MixOneColumnInst_2_n183 ;
    wire MixColumnsIns_MixOneColumnInst_2_n182 ;
    wire MixColumnsIns_MixOneColumnInst_2_n181 ;
    wire MixColumnsIns_MixOneColumnInst_2_n180 ;
    wire MixColumnsIns_MixOneColumnInst_2_n179 ;
    wire MixColumnsIns_MixOneColumnInst_2_n178 ;
    wire MixColumnsIns_MixOneColumnInst_2_n177 ;
    wire MixColumnsIns_MixOneColumnInst_2_n176 ;
    wire MixColumnsIns_MixOneColumnInst_2_n175 ;
    wire MixColumnsIns_MixOneColumnInst_2_n174 ;
    wire MixColumnsIns_MixOneColumnInst_2_n173 ;
    wire MixColumnsIns_MixOneColumnInst_2_n172 ;
    wire MixColumnsIns_MixOneColumnInst_2_n171 ;
    wire MixColumnsIns_MixOneColumnInst_2_n170 ;
    wire MixColumnsIns_MixOneColumnInst_2_n169 ;
    wire MixColumnsIns_MixOneColumnInst_2_n168 ;
    wire MixColumnsIns_MixOneColumnInst_2_n167 ;
    wire MixColumnsIns_MixOneColumnInst_2_n166 ;
    wire MixColumnsIns_MixOneColumnInst_2_n165 ;
    wire MixColumnsIns_MixOneColumnInst_2_n164 ;
    wire MixColumnsIns_MixOneColumnInst_2_n163 ;
    wire MixColumnsIns_MixOneColumnInst_2_n162 ;
    wire MixColumnsIns_MixOneColumnInst_2_n161 ;
    wire MixColumnsIns_MixOneColumnInst_2_n160 ;
    wire MixColumnsIns_MixOneColumnInst_2_n159 ;
    wire MixColumnsIns_MixOneColumnInst_2_n158 ;
    wire MixColumnsIns_MixOneColumnInst_2_n157 ;
    wire MixColumnsIns_MixOneColumnInst_2_n156 ;
    wire MixColumnsIns_MixOneColumnInst_2_n155 ;
    wire MixColumnsIns_MixOneColumnInst_2_n154 ;
    wire MixColumnsIns_MixOneColumnInst_2_n153 ;
    wire MixColumnsIns_MixOneColumnInst_2_n152 ;
    wire MixColumnsIns_MixOneColumnInst_2_n151 ;
    wire MixColumnsIns_MixOneColumnInst_2_n150 ;
    wire MixColumnsIns_MixOneColumnInst_2_n149 ;
    wire MixColumnsIns_MixOneColumnInst_2_n148 ;
    wire MixColumnsIns_MixOneColumnInst_2_n147 ;
    wire MixColumnsIns_MixOneColumnInst_2_n146 ;
    wire MixColumnsIns_MixOneColumnInst_2_n145 ;
    wire MixColumnsIns_MixOneColumnInst_2_n144 ;
    wire MixColumnsIns_MixOneColumnInst_2_n143 ;
    wire MixColumnsIns_MixOneColumnInst_2_n142 ;
    wire MixColumnsIns_MixOneColumnInst_2_n141 ;
    wire MixColumnsIns_MixOneColumnInst_2_n140 ;
    wire MixColumnsIns_MixOneColumnInst_2_n139 ;
    wire MixColumnsIns_MixOneColumnInst_2_n138 ;
    wire MixColumnsIns_MixOneColumnInst_2_n137 ;
    wire MixColumnsIns_MixOneColumnInst_2_n136 ;
    wire MixColumnsIns_MixOneColumnInst_2_n135 ;
    wire MixColumnsIns_MixOneColumnInst_2_n134 ;
    wire MixColumnsIns_MixOneColumnInst_2_n133 ;
    wire MixColumnsIns_MixOneColumnInst_2_n132 ;
    wire MixColumnsIns_MixOneColumnInst_2_n131 ;
    wire MixColumnsIns_MixOneColumnInst_2_n130 ;
    wire MixColumnsIns_MixOneColumnInst_2_n129 ;
    wire MixColumnsIns_MixOneColumnInst_3_n192 ;
    wire MixColumnsIns_MixOneColumnInst_3_n191 ;
    wire MixColumnsIns_MixOneColumnInst_3_n190 ;
    wire MixColumnsIns_MixOneColumnInst_3_n189 ;
    wire MixColumnsIns_MixOneColumnInst_3_n188 ;
    wire MixColumnsIns_MixOneColumnInst_3_n187 ;
    wire MixColumnsIns_MixOneColumnInst_3_n186 ;
    wire MixColumnsIns_MixOneColumnInst_3_n185 ;
    wire MixColumnsIns_MixOneColumnInst_3_n184 ;
    wire MixColumnsIns_MixOneColumnInst_3_n183 ;
    wire MixColumnsIns_MixOneColumnInst_3_n182 ;
    wire MixColumnsIns_MixOneColumnInst_3_n181 ;
    wire MixColumnsIns_MixOneColumnInst_3_n180 ;
    wire MixColumnsIns_MixOneColumnInst_3_n179 ;
    wire MixColumnsIns_MixOneColumnInst_3_n178 ;
    wire MixColumnsIns_MixOneColumnInst_3_n177 ;
    wire MixColumnsIns_MixOneColumnInst_3_n176 ;
    wire MixColumnsIns_MixOneColumnInst_3_n175 ;
    wire MixColumnsIns_MixOneColumnInst_3_n174 ;
    wire MixColumnsIns_MixOneColumnInst_3_n173 ;
    wire MixColumnsIns_MixOneColumnInst_3_n172 ;
    wire MixColumnsIns_MixOneColumnInst_3_n171 ;
    wire MixColumnsIns_MixOneColumnInst_3_n170 ;
    wire MixColumnsIns_MixOneColumnInst_3_n169 ;
    wire MixColumnsIns_MixOneColumnInst_3_n168 ;
    wire MixColumnsIns_MixOneColumnInst_3_n167 ;
    wire MixColumnsIns_MixOneColumnInst_3_n166 ;
    wire MixColumnsIns_MixOneColumnInst_3_n165 ;
    wire MixColumnsIns_MixOneColumnInst_3_n164 ;
    wire MixColumnsIns_MixOneColumnInst_3_n163 ;
    wire MixColumnsIns_MixOneColumnInst_3_n162 ;
    wire MixColumnsIns_MixOneColumnInst_3_n161 ;
    wire MixColumnsIns_MixOneColumnInst_3_n160 ;
    wire MixColumnsIns_MixOneColumnInst_3_n159 ;
    wire MixColumnsIns_MixOneColumnInst_3_n158 ;
    wire MixColumnsIns_MixOneColumnInst_3_n157 ;
    wire MixColumnsIns_MixOneColumnInst_3_n156 ;
    wire MixColumnsIns_MixOneColumnInst_3_n155 ;
    wire MixColumnsIns_MixOneColumnInst_3_n154 ;
    wire MixColumnsIns_MixOneColumnInst_3_n153 ;
    wire MixColumnsIns_MixOneColumnInst_3_n152 ;
    wire MixColumnsIns_MixOneColumnInst_3_n151 ;
    wire MixColumnsIns_MixOneColumnInst_3_n150 ;
    wire MixColumnsIns_MixOneColumnInst_3_n149 ;
    wire MixColumnsIns_MixOneColumnInst_3_n148 ;
    wire MixColumnsIns_MixOneColumnInst_3_n147 ;
    wire MixColumnsIns_MixOneColumnInst_3_n146 ;
    wire MixColumnsIns_MixOneColumnInst_3_n145 ;
    wire MixColumnsIns_MixOneColumnInst_3_n144 ;
    wire MixColumnsIns_MixOneColumnInst_3_n143 ;
    wire MixColumnsIns_MixOneColumnInst_3_n142 ;
    wire MixColumnsIns_MixOneColumnInst_3_n141 ;
    wire MixColumnsIns_MixOneColumnInst_3_n140 ;
    wire MixColumnsIns_MixOneColumnInst_3_n139 ;
    wire MixColumnsIns_MixOneColumnInst_3_n138 ;
    wire MixColumnsIns_MixOneColumnInst_3_n137 ;
    wire MixColumnsIns_MixOneColumnInst_3_n136 ;
    wire MixColumnsIns_MixOneColumnInst_3_n135 ;
    wire MixColumnsIns_MixOneColumnInst_3_n134 ;
    wire MixColumnsIns_MixOneColumnInst_3_n133 ;
    wire MixColumnsIns_MixOneColumnInst_3_n132 ;
    wire MixColumnsIns_MixOneColumnInst_3_n131 ;
    wire MixColumnsIns_MixOneColumnInst_3_n130 ;
    wire MixColumnsIns_MixOneColumnInst_3_n129 ;
    wire KeyReg_Inst_ff_SDE_0_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_0_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_1_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_1_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_2_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_2_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_3_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_3_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_4_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_4_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_5_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_5_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_6_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_6_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_7_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_7_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_8_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_8_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_9_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_9_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_10_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_10_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_11_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_11_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_12_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_12_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_13_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_13_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_14_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_14_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_15_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_15_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_16_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_16_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_17_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_17_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_18_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_18_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_19_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_19_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_20_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_20_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_21_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_21_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_22_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_22_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_23_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_23_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_24_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_24_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_25_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_25_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_26_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_26_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_27_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_27_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_28_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_28_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_29_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_29_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_30_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_30_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_31_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_31_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_32_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_32_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_33_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_33_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_34_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_34_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_35_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_35_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_36_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_36_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_37_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_37_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_38_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_38_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_39_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_39_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_40_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_40_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_41_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_41_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_42_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_42_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_43_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_43_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_44_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_44_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_45_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_45_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_46_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_46_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_47_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_47_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_48_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_48_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_49_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_49_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_50_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_50_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_51_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_51_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_52_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_52_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_53_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_53_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_54_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_54_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_55_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_55_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_56_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_56_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_57_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_57_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_58_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_58_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_59_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_59_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_60_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_60_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_61_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_61_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_62_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_62_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_63_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_63_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_64_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_64_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_65_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_65_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_66_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_66_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_67_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_67_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_68_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_68_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_69_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_69_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_70_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_70_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_71_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_71_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_72_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_72_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_73_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_73_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_74_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_74_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_75_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_75_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_76_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_76_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_77_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_77_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_78_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_78_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_79_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_79_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_80_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_80_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_81_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_81_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_82_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_82_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_83_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_83_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_84_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_84_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_85_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_85_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_86_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_86_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_87_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_87_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_88_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_88_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_89_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_89_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_90_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_90_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_91_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_91_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_92_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_92_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_93_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_93_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_94_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_94_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_95_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_95_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_96_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_96_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_97_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_97_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_98_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_98_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_99_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_99_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_100_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_100_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_101_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_101_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_102_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_102_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_103_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_103_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_104_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_104_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_105_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_105_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_106_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_106_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_107_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_107_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_108_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_108_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_109_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_109_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_110_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_110_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_111_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_111_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_112_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_112_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_113_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_113_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_114_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_114_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_115_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_115_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_116_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_116_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_117_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_117_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_118_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_118_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_119_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_119_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_120_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_120_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_121_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_121_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_122_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_122_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_123_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_123_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_124_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_124_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_125_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_125_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_126_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_126_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_127_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_127_MUX_inst_X ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_ ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n3 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n1 ;
    wire [127:0] RoundOutput ;
    wire [127:0] RoundInput ;
    wire [127:0] RoundKey ;
    wire [123:0] MixColumnsInput ;
    wire [127:0] MixColumnsOutput ;
    wire [127:0] KeyExpansionOutput ;
    wire [5:0] Rcon ;
    wire [3:0] RoundCounter ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_0_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_1_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_2_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_3_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10445 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10453 ;
    wire new_AGEMA_signal_10454 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10550 ;
    wire new_AGEMA_signal_10551 ;
    wire new_AGEMA_signal_10552 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10556 ;
    wire new_AGEMA_signal_10557 ;
    wire new_AGEMA_signal_10558 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10562 ;
    wire new_AGEMA_signal_10563 ;
    wire new_AGEMA_signal_10564 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10568 ;
    wire new_AGEMA_signal_10569 ;
    wire new_AGEMA_signal_10570 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10574 ;
    wire new_AGEMA_signal_10575 ;
    wire new_AGEMA_signal_10576 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10589 ;
    wire new_AGEMA_signal_10590 ;
    wire new_AGEMA_signal_10591 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10595 ;
    wire new_AGEMA_signal_10596 ;
    wire new_AGEMA_signal_10597 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10601 ;
    wire new_AGEMA_signal_10602 ;
    wire new_AGEMA_signal_10603 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10607 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10609 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10636 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10642 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10654 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10706 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10730 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10746 ;
    wire new_AGEMA_signal_10747 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10763 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10777 ;
    wire new_AGEMA_signal_10778 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10781 ;
    wire new_AGEMA_signal_10782 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10785 ;
    wire new_AGEMA_signal_10786 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10789 ;
    wire new_AGEMA_signal_10790 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10793 ;
    wire new_AGEMA_signal_10794 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10797 ;
    wire new_AGEMA_signal_10798 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10801 ;
    wire new_AGEMA_signal_10802 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10805 ;
    wire new_AGEMA_signal_10806 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10809 ;
    wire new_AGEMA_signal_10810 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10813 ;
    wire new_AGEMA_signal_10814 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10817 ;
    wire new_AGEMA_signal_10818 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10821 ;
    wire new_AGEMA_signal_10822 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10825 ;
    wire new_AGEMA_signal_10826 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10829 ;
    wire new_AGEMA_signal_10830 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10833 ;
    wire new_AGEMA_signal_10834 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10837 ;
    wire new_AGEMA_signal_10838 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10841 ;
    wire new_AGEMA_signal_10842 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10845 ;
    wire new_AGEMA_signal_10846 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10849 ;
    wire new_AGEMA_signal_10850 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10853 ;
    wire new_AGEMA_signal_10854 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10857 ;
    wire new_AGEMA_signal_10858 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10861 ;
    wire new_AGEMA_signal_10862 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10865 ;
    wire new_AGEMA_signal_10866 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10869 ;
    wire new_AGEMA_signal_10870 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10873 ;
    wire new_AGEMA_signal_10874 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11197 ;
    wire new_AGEMA_signal_11198 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11201 ;
    wire new_AGEMA_signal_11202 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11205 ;
    wire new_AGEMA_signal_11206 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11209 ;
    wire new_AGEMA_signal_11210 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11213 ;
    wire new_AGEMA_signal_11214 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11217 ;
    wire new_AGEMA_signal_11218 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11221 ;
    wire new_AGEMA_signal_11222 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11225 ;
    wire new_AGEMA_signal_11226 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11229 ;
    wire new_AGEMA_signal_11230 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11233 ;
    wire new_AGEMA_signal_11234 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11237 ;
    wire new_AGEMA_signal_11238 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11241 ;
    wire new_AGEMA_signal_11242 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11245 ;
    wire new_AGEMA_signal_11246 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11249 ;
    wire new_AGEMA_signal_11250 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11253 ;
    wire new_AGEMA_signal_11254 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11257 ;
    wire new_AGEMA_signal_11258 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11261 ;
    wire new_AGEMA_signal_11262 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11265 ;
    wire new_AGEMA_signal_11266 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11269 ;
    wire new_AGEMA_signal_11270 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11273 ;
    wire new_AGEMA_signal_11274 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11277 ;
    wire new_AGEMA_signal_11278 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11281 ;
    wire new_AGEMA_signal_11282 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11285 ;
    wire new_AGEMA_signal_11286 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11289 ;
    wire new_AGEMA_signal_11290 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11293 ;
    wire new_AGEMA_signal_11294 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11297 ;
    wire new_AGEMA_signal_11298 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11301 ;
    wire new_AGEMA_signal_11302 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11305 ;
    wire new_AGEMA_signal_11306 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11309 ;
    wire new_AGEMA_signal_11310 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11313 ;
    wire new_AGEMA_signal_11314 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11317 ;
    wire new_AGEMA_signal_11318 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11321 ;
    wire new_AGEMA_signal_11322 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11612 ;
    wire new_AGEMA_signal_11613 ;
    wire new_AGEMA_signal_11614 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11642 ;
    wire new_AGEMA_signal_11643 ;
    wire new_AGEMA_signal_11644 ;
    wire new_AGEMA_signal_11645 ;
    wire new_AGEMA_signal_11646 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11648 ;
    wire new_AGEMA_signal_11649 ;
    wire new_AGEMA_signal_11650 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11653 ;
    wire new_AGEMA_signal_11654 ;
    wire new_AGEMA_signal_11655 ;
    wire new_AGEMA_signal_11656 ;
    wire new_AGEMA_signal_11657 ;
    wire new_AGEMA_signal_11658 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11660 ;
    wire new_AGEMA_signal_11661 ;
    wire new_AGEMA_signal_11662 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11665 ;
    wire new_AGEMA_signal_11666 ;
    wire new_AGEMA_signal_11667 ;
    wire new_AGEMA_signal_11668 ;
    wire new_AGEMA_signal_11669 ;
    wire new_AGEMA_signal_11670 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11672 ;
    wire new_AGEMA_signal_11673 ;
    wire new_AGEMA_signal_11674 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11677 ;
    wire new_AGEMA_signal_11678 ;
    wire new_AGEMA_signal_11679 ;
    wire new_AGEMA_signal_11680 ;
    wire new_AGEMA_signal_11681 ;
    wire new_AGEMA_signal_11682 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11685 ;
    wire new_AGEMA_signal_11686 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11689 ;
    wire new_AGEMA_signal_11690 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11693 ;
    wire new_AGEMA_signal_11694 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11697 ;
    wire new_AGEMA_signal_11698 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11701 ;
    wire new_AGEMA_signal_11702 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11705 ;
    wire new_AGEMA_signal_11706 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11709 ;
    wire new_AGEMA_signal_11710 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11713 ;
    wire new_AGEMA_signal_11714 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11717 ;
    wire new_AGEMA_signal_11718 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11721 ;
    wire new_AGEMA_signal_11722 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11725 ;
    wire new_AGEMA_signal_11726 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11729 ;
    wire new_AGEMA_signal_11730 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11733 ;
    wire new_AGEMA_signal_11734 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11737 ;
    wire new_AGEMA_signal_11738 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11741 ;
    wire new_AGEMA_signal_11742 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11745 ;
    wire new_AGEMA_signal_11746 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11749 ;
    wire new_AGEMA_signal_11750 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11753 ;
    wire new_AGEMA_signal_11754 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11757 ;
    wire new_AGEMA_signal_11758 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11761 ;
    wire new_AGEMA_signal_11762 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11765 ;
    wire new_AGEMA_signal_11766 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11769 ;
    wire new_AGEMA_signal_11770 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;
    wire new_AGEMA_signal_11777 ;
    wire new_AGEMA_signal_11778 ;
    wire new_AGEMA_signal_11779 ;
    wire new_AGEMA_signal_11780 ;
    wire new_AGEMA_signal_11781 ;
    wire new_AGEMA_signal_11782 ;
    wire new_AGEMA_signal_11783 ;
    wire new_AGEMA_signal_11784 ;
    wire new_AGEMA_signal_11785 ;
    wire new_AGEMA_signal_11786 ;
    wire new_AGEMA_signal_11787 ;
    wire new_AGEMA_signal_11788 ;
    wire new_AGEMA_signal_11789 ;
    wire new_AGEMA_signal_11790 ;
    wire new_AGEMA_signal_11791 ;
    wire new_AGEMA_signal_11792 ;
    wire new_AGEMA_signal_11793 ;
    wire new_AGEMA_signal_11794 ;
    wire new_AGEMA_signal_11795 ;
    wire new_AGEMA_signal_11796 ;
    wire new_AGEMA_signal_11797 ;
    wire new_AGEMA_signal_11798 ;
    wire new_AGEMA_signal_11799 ;
    wire new_AGEMA_signal_11800 ;
    wire new_AGEMA_signal_11801 ;
    wire new_AGEMA_signal_11802 ;
    wire new_AGEMA_signal_11803 ;
    wire new_AGEMA_signal_11804 ;
    wire new_AGEMA_signal_11805 ;
    wire new_AGEMA_signal_11806 ;
    wire new_AGEMA_signal_11807 ;
    wire new_AGEMA_signal_11808 ;
    wire new_AGEMA_signal_11809 ;
    wire new_AGEMA_signal_11810 ;
    wire new_AGEMA_signal_11811 ;
    wire new_AGEMA_signal_11812 ;
    wire new_AGEMA_signal_11813 ;
    wire new_AGEMA_signal_11814 ;
    wire new_AGEMA_signal_11815 ;
    wire new_AGEMA_signal_11816 ;
    wire new_AGEMA_signal_11817 ;
    wire new_AGEMA_signal_11818 ;
    wire new_AGEMA_signal_11819 ;
    wire new_AGEMA_signal_11820 ;
    wire new_AGEMA_signal_11821 ;
    wire new_AGEMA_signal_11822 ;
    wire new_AGEMA_signal_11823 ;
    wire new_AGEMA_signal_11824 ;
    wire new_AGEMA_signal_11825 ;
    wire new_AGEMA_signal_11826 ;
    wire new_AGEMA_signal_11827 ;
    wire new_AGEMA_signal_11828 ;
    wire new_AGEMA_signal_11829 ;
    wire new_AGEMA_signal_11830 ;
    wire new_AGEMA_signal_11831 ;
    wire new_AGEMA_signal_11832 ;
    wire new_AGEMA_signal_11833 ;
    wire new_AGEMA_signal_11834 ;
    wire new_AGEMA_signal_11835 ;
    wire new_AGEMA_signal_11836 ;
    wire new_AGEMA_signal_11837 ;
    wire new_AGEMA_signal_11838 ;
    wire new_AGEMA_signal_11839 ;
    wire new_AGEMA_signal_11840 ;
    wire new_AGEMA_signal_11841 ;
    wire new_AGEMA_signal_11842 ;
    wire new_AGEMA_signal_11843 ;
    wire new_AGEMA_signal_11844 ;
    wire new_AGEMA_signal_11845 ;
    wire new_AGEMA_signal_11846 ;
    wire new_AGEMA_signal_11847 ;
    wire new_AGEMA_signal_11848 ;
    wire new_AGEMA_signal_11849 ;
    wire new_AGEMA_signal_11850 ;
    wire new_AGEMA_signal_11851 ;
    wire new_AGEMA_signal_11852 ;
    wire new_AGEMA_signal_11853 ;
    wire new_AGEMA_signal_11854 ;
    wire new_AGEMA_signal_11855 ;
    wire new_AGEMA_signal_11856 ;
    wire new_AGEMA_signal_11857 ;
    wire new_AGEMA_signal_11858 ;
    wire new_AGEMA_signal_11859 ;
    wire new_AGEMA_signal_11860 ;
    wire new_AGEMA_signal_11861 ;
    wire new_AGEMA_signal_11862 ;
    wire new_AGEMA_signal_11863 ;
    wire new_AGEMA_signal_11864 ;
    wire new_AGEMA_signal_11865 ;
    wire new_AGEMA_signal_11866 ;
    wire new_AGEMA_signal_11867 ;
    wire new_AGEMA_signal_11868 ;
    wire new_AGEMA_signal_11869 ;
    wire new_AGEMA_signal_11870 ;
    wire new_AGEMA_signal_11871 ;
    wire new_AGEMA_signal_11872 ;
    wire new_AGEMA_signal_11873 ;
    wire new_AGEMA_signal_11874 ;
    wire new_AGEMA_signal_11875 ;
    wire new_AGEMA_signal_11876 ;
    wire new_AGEMA_signal_11877 ;
    wire new_AGEMA_signal_11878 ;
    wire new_AGEMA_signal_11879 ;
    wire new_AGEMA_signal_11880 ;
    wire new_AGEMA_signal_11881 ;
    wire new_AGEMA_signal_11882 ;
    wire new_AGEMA_signal_11883 ;
    wire new_AGEMA_signal_11884 ;
    wire new_AGEMA_signal_11885 ;
    wire new_AGEMA_signal_11886 ;
    wire new_AGEMA_signal_11887 ;
    wire new_AGEMA_signal_11888 ;
    wire new_AGEMA_signal_11889 ;
    wire new_AGEMA_signal_11890 ;
    wire new_AGEMA_signal_11891 ;
    wire new_AGEMA_signal_11892 ;
    wire new_AGEMA_signal_11893 ;
    wire new_AGEMA_signal_11894 ;
    wire new_AGEMA_signal_11895 ;
    wire new_AGEMA_signal_11896 ;
    wire new_AGEMA_signal_11897 ;
    wire new_AGEMA_signal_11898 ;
    wire new_AGEMA_signal_11899 ;
    wire new_AGEMA_signal_11900 ;
    wire new_AGEMA_signal_11901 ;
    wire new_AGEMA_signal_11902 ;
    wire new_AGEMA_signal_11903 ;
    wire new_AGEMA_signal_11904 ;
    wire new_AGEMA_signal_11905 ;
    wire new_AGEMA_signal_11906 ;
    wire new_AGEMA_signal_11907 ;
    wire new_AGEMA_signal_11908 ;
    wire new_AGEMA_signal_11909 ;
    wire new_AGEMA_signal_11910 ;
    wire new_AGEMA_signal_11911 ;
    wire new_AGEMA_signal_11912 ;
    wire new_AGEMA_signal_11913 ;
    wire new_AGEMA_signal_11914 ;
    wire new_AGEMA_signal_11915 ;
    wire new_AGEMA_signal_11916 ;
    wire new_AGEMA_signal_11917 ;
    wire new_AGEMA_signal_11918 ;
    wire new_AGEMA_signal_11919 ;
    wire new_AGEMA_signal_11920 ;
    wire new_AGEMA_signal_11921 ;
    wire new_AGEMA_signal_11922 ;
    wire new_AGEMA_signal_11923 ;
    wire new_AGEMA_signal_11924 ;
    wire new_AGEMA_signal_11925 ;
    wire new_AGEMA_signal_11926 ;
    wire new_AGEMA_signal_11927 ;
    wire new_AGEMA_signal_11928 ;
    wire new_AGEMA_signal_11929 ;
    wire new_AGEMA_signal_11930 ;
    wire new_AGEMA_signal_11931 ;
    wire new_AGEMA_signal_11932 ;
    wire new_AGEMA_signal_11933 ;
    wire new_AGEMA_signal_11934 ;
    wire new_AGEMA_signal_11935 ;
    wire new_AGEMA_signal_11936 ;
    wire new_AGEMA_signal_11937 ;
    wire new_AGEMA_signal_11938 ;
    wire new_AGEMA_signal_11939 ;
    wire new_AGEMA_signal_11940 ;
    wire new_AGEMA_signal_11941 ;
    wire new_AGEMA_signal_11942 ;
    wire new_AGEMA_signal_11943 ;
    wire new_AGEMA_signal_11944 ;
    wire new_AGEMA_signal_11945 ;
    wire new_AGEMA_signal_11946 ;
    wire new_AGEMA_signal_11947 ;
    wire new_AGEMA_signal_11948 ;
    wire new_AGEMA_signal_11949 ;
    wire new_AGEMA_signal_11950 ;
    wire new_AGEMA_signal_11951 ;
    wire new_AGEMA_signal_11952 ;
    wire new_AGEMA_signal_11953 ;
    wire new_AGEMA_signal_11954 ;
    wire new_AGEMA_signal_11955 ;
    wire new_AGEMA_signal_11956 ;
    wire new_AGEMA_signal_11957 ;
    wire new_AGEMA_signal_11958 ;
    wire new_AGEMA_signal_11959 ;
    wire new_AGEMA_signal_11960 ;
    wire new_AGEMA_signal_11961 ;
    wire new_AGEMA_signal_11962 ;
    wire new_AGEMA_signal_11963 ;
    wire new_AGEMA_signal_11964 ;
    wire new_AGEMA_signal_11965 ;
    wire new_AGEMA_signal_11966 ;
    wire new_AGEMA_signal_11967 ;
    wire new_AGEMA_signal_11968 ;
    wire new_AGEMA_signal_11969 ;
    wire new_AGEMA_signal_11970 ;
    wire new_AGEMA_signal_11971 ;
    wire new_AGEMA_signal_11972 ;
    wire new_AGEMA_signal_11973 ;
    wire new_AGEMA_signal_11974 ;
    wire new_AGEMA_signal_11975 ;
    wire new_AGEMA_signal_11976 ;
    wire new_AGEMA_signal_11977 ;
    wire new_AGEMA_signal_11978 ;
    wire new_AGEMA_signal_11979 ;
    wire new_AGEMA_signal_11980 ;
    wire new_AGEMA_signal_11981 ;
    wire new_AGEMA_signal_11982 ;
    wire new_AGEMA_signal_11983 ;
    wire new_AGEMA_signal_11984 ;
    wire new_AGEMA_signal_11985 ;
    wire new_AGEMA_signal_11986 ;
    wire new_AGEMA_signal_11987 ;
    wire new_AGEMA_signal_11988 ;
    wire new_AGEMA_signal_11989 ;
    wire new_AGEMA_signal_11990 ;
    wire new_AGEMA_signal_11991 ;
    wire new_AGEMA_signal_11992 ;
    wire new_AGEMA_signal_11993 ;
    wire new_AGEMA_signal_11994 ;
    wire new_AGEMA_signal_11995 ;
    wire new_AGEMA_signal_11996 ;
    wire new_AGEMA_signal_11997 ;
    wire new_AGEMA_signal_11998 ;
    wire new_AGEMA_signal_11999 ;
    wire new_AGEMA_signal_12000 ;
    wire new_AGEMA_signal_12001 ;
    wire new_AGEMA_signal_12002 ;
    wire new_AGEMA_signal_12003 ;
    wire new_AGEMA_signal_12004 ;
    wire new_AGEMA_signal_12005 ;
    wire new_AGEMA_signal_12006 ;
    wire new_AGEMA_signal_12007 ;
    wire new_AGEMA_signal_12008 ;
    wire new_AGEMA_signal_12009 ;
    wire new_AGEMA_signal_12010 ;
    wire new_AGEMA_signal_12011 ;
    wire new_AGEMA_signal_12012 ;
    wire new_AGEMA_signal_12013 ;
    wire new_AGEMA_signal_12014 ;
    wire new_AGEMA_signal_12015 ;
    wire new_AGEMA_signal_12016 ;
    wire new_AGEMA_signal_12017 ;
    wire new_AGEMA_signal_12018 ;
    wire new_AGEMA_signal_12019 ;
    wire new_AGEMA_signal_12020 ;
    wire new_AGEMA_signal_12021 ;
    wire new_AGEMA_signal_12022 ;
    wire new_AGEMA_signal_12023 ;
    wire new_AGEMA_signal_12024 ;
    wire new_AGEMA_signal_12025 ;
    wire new_AGEMA_signal_12026 ;
    wire new_AGEMA_signal_12027 ;
    wire new_AGEMA_signal_12028 ;
    wire new_AGEMA_signal_12029 ;
    wire new_AGEMA_signal_12030 ;
    wire new_AGEMA_signal_12031 ;
    wire new_AGEMA_signal_12032 ;
    wire new_AGEMA_signal_12033 ;
    wire new_AGEMA_signal_12034 ;
    wire new_AGEMA_signal_12035 ;
    wire new_AGEMA_signal_12036 ;
    wire new_AGEMA_signal_12037 ;
    wire new_AGEMA_signal_12038 ;
    wire new_AGEMA_signal_12039 ;
    wire new_AGEMA_signal_12040 ;
    wire new_AGEMA_signal_12041 ;
    wire new_AGEMA_signal_12042 ;
    wire new_AGEMA_signal_12043 ;
    wire new_AGEMA_signal_12044 ;
    wire new_AGEMA_signal_12045 ;
    wire new_AGEMA_signal_12046 ;
    wire new_AGEMA_signal_12047 ;
    wire new_AGEMA_signal_12048 ;
    wire new_AGEMA_signal_12049 ;
    wire new_AGEMA_signal_12050 ;
    wire new_AGEMA_signal_12051 ;
    wire new_AGEMA_signal_12052 ;
    wire new_AGEMA_signal_12053 ;
    wire new_AGEMA_signal_12054 ;
    wire new_AGEMA_signal_12055 ;
    wire new_AGEMA_signal_12056 ;
    wire new_AGEMA_signal_12057 ;
    wire new_AGEMA_signal_12058 ;
    wire new_AGEMA_signal_12059 ;
    wire new_AGEMA_signal_12060 ;
    wire new_AGEMA_signal_12061 ;
    wire new_AGEMA_signal_12062 ;
    wire new_AGEMA_signal_12063 ;
    wire new_AGEMA_signal_12064 ;
    wire new_AGEMA_signal_12065 ;
    wire new_AGEMA_signal_12066 ;
    wire new_AGEMA_signal_12067 ;
    wire new_AGEMA_signal_12068 ;
    wire new_AGEMA_signal_12069 ;
    wire new_AGEMA_signal_12070 ;
    wire new_AGEMA_signal_12071 ;
    wire new_AGEMA_signal_12072 ;
    wire new_AGEMA_signal_12073 ;
    wire new_AGEMA_signal_12074 ;
    wire new_AGEMA_signal_12075 ;
    wire new_AGEMA_signal_12076 ;
    wire new_AGEMA_signal_12077 ;
    wire new_AGEMA_signal_12078 ;
    wire new_AGEMA_signal_12079 ;
    wire new_AGEMA_signal_12080 ;
    wire new_AGEMA_signal_12081 ;
    wire new_AGEMA_signal_12082 ;
    wire new_AGEMA_signal_12083 ;
    wire new_AGEMA_signal_12084 ;
    wire new_AGEMA_signal_12085 ;
    wire new_AGEMA_signal_12086 ;
    wire new_AGEMA_signal_12087 ;
    wire new_AGEMA_signal_12088 ;
    wire new_AGEMA_signal_12089 ;
    wire new_AGEMA_signal_12090 ;
    wire new_AGEMA_signal_12091 ;
    wire new_AGEMA_signal_12092 ;
    wire new_AGEMA_signal_12093 ;
    wire new_AGEMA_signal_12094 ;
    wire new_AGEMA_signal_12095 ;
    wire new_AGEMA_signal_12096 ;
    wire new_AGEMA_signal_12097 ;
    wire new_AGEMA_signal_12098 ;
    wire new_AGEMA_signal_12099 ;
    wire new_AGEMA_signal_12100 ;
    wire new_AGEMA_signal_12101 ;
    wire new_AGEMA_signal_12102 ;
    wire new_AGEMA_signal_12103 ;
    wire new_AGEMA_signal_12104 ;
    wire new_AGEMA_signal_12105 ;
    wire new_AGEMA_signal_12106 ;
    wire new_AGEMA_signal_12107 ;
    wire new_AGEMA_signal_12108 ;
    wire new_AGEMA_signal_12109 ;
    wire new_AGEMA_signal_12110 ;
    wire new_AGEMA_signal_12111 ;
    wire new_AGEMA_signal_12112 ;
    wire new_AGEMA_signal_12113 ;
    wire new_AGEMA_signal_12114 ;
    wire new_AGEMA_signal_12115 ;
    wire new_AGEMA_signal_12116 ;
    wire new_AGEMA_signal_12117 ;
    wire new_AGEMA_signal_12118 ;
    wire new_AGEMA_signal_12119 ;
    wire new_AGEMA_signal_12120 ;
    wire new_AGEMA_signal_12121 ;
    wire new_AGEMA_signal_12122 ;
    wire new_AGEMA_signal_12123 ;
    wire new_AGEMA_signal_12124 ;
    wire new_AGEMA_signal_12125 ;
    wire new_AGEMA_signal_12126 ;
    wire new_AGEMA_signal_12127 ;
    wire new_AGEMA_signal_12128 ;
    wire new_AGEMA_signal_12129 ;
    wire new_AGEMA_signal_12130 ;
    wire new_AGEMA_signal_12131 ;
    wire new_AGEMA_signal_12132 ;
    wire new_AGEMA_signal_12133 ;
    wire new_AGEMA_signal_12134 ;
    wire new_AGEMA_signal_12135 ;
    wire new_AGEMA_signal_12136 ;
    wire new_AGEMA_signal_12137 ;
    wire new_AGEMA_signal_12138 ;
    wire new_AGEMA_signal_12139 ;
    wire new_AGEMA_signal_12140 ;
    wire new_AGEMA_signal_12141 ;
    wire new_AGEMA_signal_12142 ;
    wire new_AGEMA_signal_12143 ;
    wire new_AGEMA_signal_12144 ;
    wire new_AGEMA_signal_12145 ;
    wire new_AGEMA_signal_12146 ;
    wire new_AGEMA_signal_12147 ;
    wire new_AGEMA_signal_12148 ;
    wire new_AGEMA_signal_12149 ;
    wire new_AGEMA_signal_12150 ;
    wire new_AGEMA_signal_12151 ;
    wire new_AGEMA_signal_12152 ;
    wire new_AGEMA_signal_12153 ;
    wire new_AGEMA_signal_12154 ;
    wire new_AGEMA_signal_12155 ;
    wire new_AGEMA_signal_12156 ;
    wire new_AGEMA_signal_12157 ;
    wire new_AGEMA_signal_12158 ;
    wire new_AGEMA_signal_12159 ;
    wire new_AGEMA_signal_12160 ;
    wire new_AGEMA_signal_12161 ;
    wire new_AGEMA_signal_12162 ;
    wire new_AGEMA_signal_12163 ;
    wire new_AGEMA_signal_12164 ;
    wire new_AGEMA_signal_12165 ;
    wire new_AGEMA_signal_12166 ;
    wire new_AGEMA_signal_12167 ;
    wire new_AGEMA_signal_12168 ;
    wire new_AGEMA_signal_12169 ;
    wire new_AGEMA_signal_12170 ;
    wire new_AGEMA_signal_12171 ;
    wire new_AGEMA_signal_12172 ;
    wire new_AGEMA_signal_12173 ;
    wire new_AGEMA_signal_12174 ;
    wire new_AGEMA_signal_12175 ;
    wire new_AGEMA_signal_12176 ;
    wire new_AGEMA_signal_12177 ;
    wire new_AGEMA_signal_12178 ;
    wire new_AGEMA_signal_12179 ;
    wire new_AGEMA_signal_12180 ;
    wire new_AGEMA_signal_12181 ;
    wire new_AGEMA_signal_12182 ;
    wire new_AGEMA_signal_12183 ;
    wire new_AGEMA_signal_12184 ;
    wire new_AGEMA_signal_12185 ;
    wire new_AGEMA_signal_12186 ;
    wire new_AGEMA_signal_12187 ;
    wire new_AGEMA_signal_12188 ;
    wire new_AGEMA_signal_12189 ;
    wire new_AGEMA_signal_12190 ;
    wire new_AGEMA_signal_12191 ;
    wire new_AGEMA_signal_12192 ;
    wire new_AGEMA_signal_12193 ;
    wire new_AGEMA_signal_12194 ;
    wire new_AGEMA_signal_12195 ;
    wire new_AGEMA_signal_12196 ;
    wire new_AGEMA_signal_12197 ;
    wire new_AGEMA_signal_12198 ;
    wire new_AGEMA_signal_12199 ;
    wire new_AGEMA_signal_12200 ;
    wire new_AGEMA_signal_12201 ;
    wire new_AGEMA_signal_12202 ;
    wire new_AGEMA_signal_12203 ;
    wire new_AGEMA_signal_12204 ;
    wire new_AGEMA_signal_12205 ;
    wire new_AGEMA_signal_12206 ;
    wire new_AGEMA_signal_12207 ;
    wire new_AGEMA_signal_12208 ;
    wire new_AGEMA_signal_12209 ;
    wire new_AGEMA_signal_12210 ;
    wire new_AGEMA_signal_12211 ;
    wire new_AGEMA_signal_12212 ;
    wire new_AGEMA_signal_12213 ;
    wire new_AGEMA_signal_12214 ;
    wire new_AGEMA_signal_12215 ;
    wire new_AGEMA_signal_12216 ;
    wire new_AGEMA_signal_12217 ;
    wire new_AGEMA_signal_12218 ;
    wire new_AGEMA_signal_12219 ;
    wire new_AGEMA_signal_12220 ;
    wire new_AGEMA_signal_12221 ;
    wire new_AGEMA_signal_12222 ;
    wire new_AGEMA_signal_12223 ;
    wire new_AGEMA_signal_12224 ;
    wire new_AGEMA_signal_12225 ;
    wire new_AGEMA_signal_12226 ;
    wire new_AGEMA_signal_12227 ;
    wire new_AGEMA_signal_12228 ;
    wire new_AGEMA_signal_12229 ;
    wire new_AGEMA_signal_12230 ;
    wire new_AGEMA_signal_12231 ;
    wire new_AGEMA_signal_12232 ;
    wire new_AGEMA_signal_12233 ;
    wire new_AGEMA_signal_12234 ;
    wire new_AGEMA_signal_12235 ;
    wire new_AGEMA_signal_12236 ;
    wire new_AGEMA_signal_12237 ;
    wire new_AGEMA_signal_12238 ;
    wire new_AGEMA_signal_12239 ;
    wire new_AGEMA_signal_12240 ;
    wire new_AGEMA_signal_12241 ;
    wire new_AGEMA_signal_12242 ;
    wire new_AGEMA_signal_12243 ;
    wire new_AGEMA_signal_12244 ;
    wire new_AGEMA_signal_12245 ;
    wire new_AGEMA_signal_12246 ;
    wire new_AGEMA_signal_12247 ;
    wire new_AGEMA_signal_12248 ;
    wire new_AGEMA_signal_12249 ;
    wire new_AGEMA_signal_12250 ;
    wire new_AGEMA_signal_12251 ;
    wire new_AGEMA_signal_12252 ;
    wire new_AGEMA_signal_12253 ;
    wire new_AGEMA_signal_12254 ;
    wire new_AGEMA_signal_12255 ;
    wire new_AGEMA_signal_12256 ;
    wire new_AGEMA_signal_12257 ;
    wire new_AGEMA_signal_12258 ;
    wire new_AGEMA_signal_12259 ;
    wire new_AGEMA_signal_12260 ;
    wire new_AGEMA_signal_12261 ;
    wire new_AGEMA_signal_12262 ;
    wire new_AGEMA_signal_12263 ;
    wire new_AGEMA_signal_12264 ;
    wire new_AGEMA_signal_12265 ;
    wire new_AGEMA_signal_12266 ;
    wire new_AGEMA_signal_12267 ;
    wire new_AGEMA_signal_12268 ;
    wire new_AGEMA_signal_12269 ;
    wire new_AGEMA_signal_12270 ;
    wire new_AGEMA_signal_12271 ;
    wire new_AGEMA_signal_12272 ;
    wire new_AGEMA_signal_12273 ;
    wire new_AGEMA_signal_12274 ;
    wire new_AGEMA_signal_12275 ;
    wire new_AGEMA_signal_12276 ;
    wire new_AGEMA_signal_12277 ;
    wire new_AGEMA_signal_12278 ;
    wire new_AGEMA_signal_12279 ;
    wire new_AGEMA_signal_12280 ;
    wire new_AGEMA_signal_12281 ;
    wire new_AGEMA_signal_12282 ;
    wire new_AGEMA_signal_12283 ;
    wire new_AGEMA_signal_12284 ;
    wire new_AGEMA_signal_12285 ;
    wire new_AGEMA_signal_12286 ;
    wire new_AGEMA_signal_12287 ;
    wire new_AGEMA_signal_12288 ;
    wire new_AGEMA_signal_12289 ;
    wire new_AGEMA_signal_12290 ;
    wire new_AGEMA_signal_12291 ;
    wire new_AGEMA_signal_12292 ;
    wire new_AGEMA_signal_12293 ;
    wire new_AGEMA_signal_12294 ;
    wire new_AGEMA_signal_12295 ;
    wire new_AGEMA_signal_12296 ;
    wire new_AGEMA_signal_12297 ;
    wire new_AGEMA_signal_12298 ;
    wire new_AGEMA_signal_12299 ;
    wire new_AGEMA_signal_12300 ;
    wire new_AGEMA_signal_12301 ;
    wire new_AGEMA_signal_12302 ;
    wire new_AGEMA_signal_12303 ;
    wire new_AGEMA_signal_12304 ;
    wire new_AGEMA_signal_12305 ;
    wire new_AGEMA_signal_12306 ;
    wire new_AGEMA_signal_12307 ;
    wire new_AGEMA_signal_12308 ;
    wire new_AGEMA_signal_12309 ;
    wire new_AGEMA_signal_12310 ;
    wire new_AGEMA_signal_12311 ;
    wire new_AGEMA_signal_12312 ;
    wire new_AGEMA_signal_12313 ;
    wire new_AGEMA_signal_12314 ;
    wire new_AGEMA_signal_12315 ;
    wire new_AGEMA_signal_12316 ;
    wire new_AGEMA_signal_12317 ;
    wire new_AGEMA_signal_12318 ;
    wire new_AGEMA_signal_12319 ;
    wire new_AGEMA_signal_12320 ;
    wire new_AGEMA_signal_12321 ;
    wire new_AGEMA_signal_12322 ;
    wire new_AGEMA_signal_12323 ;
    wire new_AGEMA_signal_12324 ;
    wire new_AGEMA_signal_12325 ;
    wire new_AGEMA_signal_12326 ;
    wire new_AGEMA_signal_12327 ;
    wire new_AGEMA_signal_12328 ;
    wire new_AGEMA_signal_12329 ;
    wire new_AGEMA_signal_12330 ;
    wire new_AGEMA_signal_12331 ;
    wire new_AGEMA_signal_12332 ;
    wire new_AGEMA_signal_12333 ;
    wire new_AGEMA_signal_12334 ;
    wire new_AGEMA_signal_12335 ;
    wire new_AGEMA_signal_12336 ;
    wire new_AGEMA_signal_12337 ;
    wire new_AGEMA_signal_12338 ;
    wire new_AGEMA_signal_12339 ;
    wire new_AGEMA_signal_12340 ;
    wire new_AGEMA_signal_12341 ;
    wire new_AGEMA_signal_12342 ;
    wire new_AGEMA_signal_12343 ;
    wire new_AGEMA_signal_12344 ;
    wire new_AGEMA_signal_12345 ;
    wire new_AGEMA_signal_12346 ;
    wire new_AGEMA_signal_12347 ;
    wire new_AGEMA_signal_12348 ;
    wire new_AGEMA_signal_12349 ;
    wire new_AGEMA_signal_12350 ;
    wire new_AGEMA_signal_12351 ;
    wire new_AGEMA_signal_12352 ;
    wire new_AGEMA_signal_12353 ;
    wire new_AGEMA_signal_12354 ;
    wire new_AGEMA_signal_12355 ;
    wire new_AGEMA_signal_12356 ;
    wire new_AGEMA_signal_12357 ;
    wire new_AGEMA_signal_12358 ;
    wire new_AGEMA_signal_12359 ;
    wire new_AGEMA_signal_12360 ;
    wire new_AGEMA_signal_12361 ;
    wire new_AGEMA_signal_12362 ;
    wire new_AGEMA_signal_12363 ;
    wire new_AGEMA_signal_12364 ;
    wire new_AGEMA_signal_12365 ;
    wire new_AGEMA_signal_12366 ;
    wire new_AGEMA_signal_12367 ;
    wire new_AGEMA_signal_12368 ;
    wire new_AGEMA_signal_12369 ;
    wire new_AGEMA_signal_12370 ;
    wire new_AGEMA_signal_12371 ;
    wire new_AGEMA_signal_12372 ;
    wire new_AGEMA_signal_12373 ;
    wire new_AGEMA_signal_12374 ;
    wire new_AGEMA_signal_12375 ;
    wire new_AGEMA_signal_12376 ;
    wire new_AGEMA_signal_12377 ;
    wire new_AGEMA_signal_12378 ;
    wire new_AGEMA_signal_12379 ;
    wire new_AGEMA_signal_12380 ;
    wire new_AGEMA_signal_12381 ;
    wire new_AGEMA_signal_12382 ;
    wire new_AGEMA_signal_12383 ;
    wire new_AGEMA_signal_12384 ;
    wire new_AGEMA_signal_12385 ;
    wire new_AGEMA_signal_12386 ;
    wire new_AGEMA_signal_12387 ;
    wire new_AGEMA_signal_12388 ;
    wire new_AGEMA_signal_12389 ;
    wire new_AGEMA_signal_12390 ;
    wire new_AGEMA_signal_12391 ;
    wire new_AGEMA_signal_12392 ;
    wire new_AGEMA_signal_12393 ;
    wire new_AGEMA_signal_12394 ;
    wire new_AGEMA_signal_12395 ;
    wire new_AGEMA_signal_12396 ;
    wire new_AGEMA_signal_12397 ;
    wire new_AGEMA_signal_12398 ;
    wire new_AGEMA_signal_12399 ;
    wire new_AGEMA_signal_12400 ;
    wire new_AGEMA_signal_12401 ;
    wire new_AGEMA_signal_12402 ;
    wire new_AGEMA_signal_12403 ;
    wire new_AGEMA_signal_12404 ;
    wire new_AGEMA_signal_12405 ;
    wire new_AGEMA_signal_12406 ;
    wire new_AGEMA_signal_12407 ;
    wire new_AGEMA_signal_12408 ;
    wire new_AGEMA_signal_12409 ;
    wire new_AGEMA_signal_12410 ;
    wire new_AGEMA_signal_12411 ;
    wire new_AGEMA_signal_12412 ;
    wire new_AGEMA_signal_12413 ;
    wire new_AGEMA_signal_12414 ;
    wire new_AGEMA_signal_12415 ;
    wire new_AGEMA_signal_12416 ;
    wire new_AGEMA_signal_12417 ;
    wire new_AGEMA_signal_12418 ;
    wire new_AGEMA_signal_12419 ;
    wire new_AGEMA_signal_12420 ;
    wire new_AGEMA_signal_12421 ;
    wire new_AGEMA_signal_12422 ;
    wire new_AGEMA_signal_12423 ;
    wire new_AGEMA_signal_12424 ;
    wire new_AGEMA_signal_12425 ;
    wire new_AGEMA_signal_12426 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12429 ;
    wire new_AGEMA_signal_12430 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12433 ;
    wire new_AGEMA_signal_12434 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12437 ;
    wire new_AGEMA_signal_12438 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12441 ;
    wire new_AGEMA_signal_12442 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12445 ;
    wire new_AGEMA_signal_12446 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12449 ;
    wire new_AGEMA_signal_12450 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12453 ;
    wire new_AGEMA_signal_12454 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12457 ;
    wire new_AGEMA_signal_12458 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12461 ;
    wire new_AGEMA_signal_12462 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12465 ;
    wire new_AGEMA_signal_12466 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12469 ;
    wire new_AGEMA_signal_12470 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12473 ;
    wire new_AGEMA_signal_12474 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12477 ;
    wire new_AGEMA_signal_12478 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12481 ;
    wire new_AGEMA_signal_12482 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12485 ;
    wire new_AGEMA_signal_12486 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12489 ;
    wire new_AGEMA_signal_12490 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12493 ;
    wire new_AGEMA_signal_12494 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12497 ;
    wire new_AGEMA_signal_12498 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12501 ;
    wire new_AGEMA_signal_12502 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12505 ;
    wire new_AGEMA_signal_12506 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12509 ;
    wire new_AGEMA_signal_12510 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12513 ;
    wire new_AGEMA_signal_12514 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12517 ;
    wire new_AGEMA_signal_12518 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12521 ;
    wire new_AGEMA_signal_12522 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12525 ;
    wire new_AGEMA_signal_12526 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12529 ;
    wire new_AGEMA_signal_12530 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12533 ;
    wire new_AGEMA_signal_12534 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12537 ;
    wire new_AGEMA_signal_12538 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12541 ;
    wire new_AGEMA_signal_12542 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12545 ;
    wire new_AGEMA_signal_12546 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12549 ;
    wire new_AGEMA_signal_12550 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12553 ;
    wire new_AGEMA_signal_12554 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12557 ;
    wire new_AGEMA_signal_12558 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12561 ;
    wire new_AGEMA_signal_12562 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12565 ;
    wire new_AGEMA_signal_12566 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12569 ;
    wire new_AGEMA_signal_12570 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12573 ;
    wire new_AGEMA_signal_12574 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12577 ;
    wire new_AGEMA_signal_12578 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12581 ;
    wire new_AGEMA_signal_12582 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12585 ;
    wire new_AGEMA_signal_12586 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12589 ;
    wire new_AGEMA_signal_12590 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12593 ;
    wire new_AGEMA_signal_12594 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12597 ;
    wire new_AGEMA_signal_12598 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12601 ;
    wire new_AGEMA_signal_12602 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12605 ;
    wire new_AGEMA_signal_12606 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12609 ;
    wire new_AGEMA_signal_12610 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12613 ;
    wire new_AGEMA_signal_12614 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12617 ;
    wire new_AGEMA_signal_12618 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12621 ;
    wire new_AGEMA_signal_12622 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12625 ;
    wire new_AGEMA_signal_12626 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12629 ;
    wire new_AGEMA_signal_12630 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12633 ;
    wire new_AGEMA_signal_12634 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12637 ;
    wire new_AGEMA_signal_12638 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12641 ;
    wire new_AGEMA_signal_12642 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12645 ;
    wire new_AGEMA_signal_12646 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12649 ;
    wire new_AGEMA_signal_12650 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12653 ;
    wire new_AGEMA_signal_12654 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12657 ;
    wire new_AGEMA_signal_12658 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12661 ;
    wire new_AGEMA_signal_12662 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12665 ;
    wire new_AGEMA_signal_12666 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12669 ;
    wire new_AGEMA_signal_12670 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12673 ;
    wire new_AGEMA_signal_12674 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12677 ;
    wire new_AGEMA_signal_12678 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12681 ;
    wire new_AGEMA_signal_12682 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12685 ;
    wire new_AGEMA_signal_12686 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12689 ;
    wire new_AGEMA_signal_12690 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12693 ;
    wire new_AGEMA_signal_12694 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12697 ;
    wire new_AGEMA_signal_12698 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12701 ;
    wire new_AGEMA_signal_12702 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12705 ;
    wire new_AGEMA_signal_12706 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12709 ;
    wire new_AGEMA_signal_12710 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12713 ;
    wire new_AGEMA_signal_12714 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12717 ;
    wire new_AGEMA_signal_12718 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12721 ;
    wire new_AGEMA_signal_12722 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12725 ;
    wire new_AGEMA_signal_12726 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12729 ;
    wire new_AGEMA_signal_12730 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12733 ;
    wire new_AGEMA_signal_12734 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12737 ;
    wire new_AGEMA_signal_12738 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12741 ;
    wire new_AGEMA_signal_12742 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12745 ;
    wire new_AGEMA_signal_12746 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12749 ;
    wire new_AGEMA_signal_12750 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12753 ;
    wire new_AGEMA_signal_12754 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12757 ;
    wire new_AGEMA_signal_12758 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12761 ;
    wire new_AGEMA_signal_12762 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12765 ;
    wire new_AGEMA_signal_12766 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12769 ;
    wire new_AGEMA_signal_12770 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12773 ;
    wire new_AGEMA_signal_12774 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12777 ;
    wire new_AGEMA_signal_12778 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12781 ;
    wire new_AGEMA_signal_12782 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12785 ;
    wire new_AGEMA_signal_12786 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12789 ;
    wire new_AGEMA_signal_12790 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12793 ;
    wire new_AGEMA_signal_12794 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12797 ;
    wire new_AGEMA_signal_12798 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12801 ;
    wire new_AGEMA_signal_12802 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12805 ;
    wire new_AGEMA_signal_12806 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12809 ;
    wire new_AGEMA_signal_12810 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12813 ;
    wire new_AGEMA_signal_12814 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12817 ;
    wire new_AGEMA_signal_12818 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12821 ;
    wire new_AGEMA_signal_12822 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12825 ;
    wire new_AGEMA_signal_12826 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12829 ;
    wire new_AGEMA_signal_12830 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12833 ;
    wire new_AGEMA_signal_12834 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12837 ;
    wire new_AGEMA_signal_12838 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12841 ;
    wire new_AGEMA_signal_12842 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12845 ;
    wire new_AGEMA_signal_12846 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12849 ;
    wire new_AGEMA_signal_12850 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire new_AGEMA_signal_12853 ;
    wire new_AGEMA_signal_12854 ;
    wire new_AGEMA_signal_12855 ;
    wire new_AGEMA_signal_12856 ;
    wire new_AGEMA_signal_12857 ;
    wire new_AGEMA_signal_12858 ;
    wire new_AGEMA_signal_12859 ;
    wire new_AGEMA_signal_12860 ;
    wire new_AGEMA_signal_12861 ;
    wire new_AGEMA_signal_12862 ;
    wire new_AGEMA_signal_12863 ;
    wire new_AGEMA_signal_12864 ;
    wire new_AGEMA_signal_12865 ;
    wire new_AGEMA_signal_12866 ;
    wire new_AGEMA_signal_12867 ;
    wire new_AGEMA_signal_12868 ;
    wire new_AGEMA_signal_12869 ;
    wire new_AGEMA_signal_12870 ;
    wire new_AGEMA_signal_12871 ;
    wire new_AGEMA_signal_12872 ;
    wire new_AGEMA_signal_12873 ;
    wire new_AGEMA_signal_12874 ;
    wire new_AGEMA_signal_12875 ;
    wire new_AGEMA_signal_12876 ;
    wire new_AGEMA_signal_12877 ;
    wire new_AGEMA_signal_12878 ;
    wire new_AGEMA_signal_12879 ;
    wire new_AGEMA_signal_12880 ;
    wire new_AGEMA_signal_12881 ;
    wire new_AGEMA_signal_12882 ;
    wire new_AGEMA_signal_12883 ;
    wire new_AGEMA_signal_12884 ;
    wire new_AGEMA_signal_12885 ;
    wire new_AGEMA_signal_12886 ;
    wire new_AGEMA_signal_12887 ;
    wire new_AGEMA_signal_12888 ;
    wire new_AGEMA_signal_12889 ;
    wire new_AGEMA_signal_12890 ;
    wire new_AGEMA_signal_12891 ;
    wire new_AGEMA_signal_12892 ;
    wire new_AGEMA_signal_12893 ;
    wire new_AGEMA_signal_12894 ;
    wire new_AGEMA_signal_12895 ;
    wire new_AGEMA_signal_12896 ;
    wire new_AGEMA_signal_12897 ;
    wire new_AGEMA_signal_12898 ;
    wire new_AGEMA_signal_12899 ;
    wire new_AGEMA_signal_12900 ;
    wire new_AGEMA_signal_12901 ;
    wire new_AGEMA_signal_12902 ;
    wire new_AGEMA_signal_12903 ;
    wire new_AGEMA_signal_12904 ;
    wire new_AGEMA_signal_12905 ;
    wire new_AGEMA_signal_12906 ;
    wire new_AGEMA_signal_12907 ;
    wire new_AGEMA_signal_12908 ;
    wire new_AGEMA_signal_12909 ;
    wire new_AGEMA_signal_12910 ;
    wire new_AGEMA_signal_12911 ;
    wire new_AGEMA_signal_12912 ;
    wire new_AGEMA_signal_12913 ;
    wire new_AGEMA_signal_12914 ;
    wire new_AGEMA_signal_12915 ;
    wire new_AGEMA_signal_12916 ;
    wire new_AGEMA_signal_12917 ;
    wire new_AGEMA_signal_12918 ;
    wire new_AGEMA_signal_12919 ;
    wire new_AGEMA_signal_12920 ;
    wire new_AGEMA_signal_12921 ;
    wire new_AGEMA_signal_12922 ;
    wire new_AGEMA_signal_12923 ;
    wire new_AGEMA_signal_12924 ;
    wire new_AGEMA_signal_12925 ;
    wire new_AGEMA_signal_12926 ;
    wire new_AGEMA_signal_12927 ;
    wire new_AGEMA_signal_12928 ;
    wire new_AGEMA_signal_12929 ;
    wire new_AGEMA_signal_12930 ;
    wire new_AGEMA_signal_12931 ;
    wire new_AGEMA_signal_12932 ;
    wire new_AGEMA_signal_12933 ;
    wire new_AGEMA_signal_12934 ;
    wire new_AGEMA_signal_12935 ;
    wire new_AGEMA_signal_12936 ;
    wire new_AGEMA_signal_12937 ;
    wire new_AGEMA_signal_12938 ;
    wire new_AGEMA_signal_12939 ;
    wire new_AGEMA_signal_12940 ;
    wire new_AGEMA_signal_12941 ;
    wire new_AGEMA_signal_12942 ;
    wire new_AGEMA_signal_12943 ;
    wire new_AGEMA_signal_12944 ;
    wire new_AGEMA_signal_12945 ;
    wire new_AGEMA_signal_12946 ;
    wire new_AGEMA_signal_12947 ;
    wire new_AGEMA_signal_12948 ;
    wire new_AGEMA_signal_12949 ;
    wire new_AGEMA_signal_12950 ;
    wire new_AGEMA_signal_12951 ;
    wire new_AGEMA_signal_12952 ;
    wire new_AGEMA_signal_12953 ;
    wire new_AGEMA_signal_12954 ;
    wire new_AGEMA_signal_12955 ;
    wire new_AGEMA_signal_12956 ;
    wire new_AGEMA_signal_12957 ;
    wire new_AGEMA_signal_12958 ;
    wire new_AGEMA_signal_12959 ;
    wire new_AGEMA_signal_12960 ;
    wire new_AGEMA_signal_12961 ;
    wire new_AGEMA_signal_12962 ;
    wire new_AGEMA_signal_12963 ;
    wire new_AGEMA_signal_12964 ;
    wire new_AGEMA_signal_12965 ;
    wire new_AGEMA_signal_12966 ;
    wire new_AGEMA_signal_12967 ;
    wire new_AGEMA_signal_12968 ;
    wire new_AGEMA_signal_12969 ;
    wire new_AGEMA_signal_12970 ;
    wire new_AGEMA_signal_12971 ;
    wire new_AGEMA_signal_12972 ;
    wire new_AGEMA_signal_12973 ;
    wire new_AGEMA_signal_12974 ;
    wire new_AGEMA_signal_12975 ;
    wire new_AGEMA_signal_12976 ;
    wire new_AGEMA_signal_12977 ;
    wire new_AGEMA_signal_12978 ;
    wire new_AGEMA_signal_12979 ;
    wire new_AGEMA_signal_12980 ;
    wire new_AGEMA_signal_12981 ;
    wire new_AGEMA_signal_12982 ;
    wire new_AGEMA_signal_12983 ;
    wire new_AGEMA_signal_12984 ;
    wire new_AGEMA_signal_12985 ;
    wire new_AGEMA_signal_12986 ;
    wire new_AGEMA_signal_12987 ;
    wire new_AGEMA_signal_12988 ;
    wire new_AGEMA_signal_12989 ;
    wire new_AGEMA_signal_12990 ;
    wire new_AGEMA_signal_12991 ;
    wire new_AGEMA_signal_12992 ;
    wire new_AGEMA_signal_12993 ;
    wire new_AGEMA_signal_12994 ;
    wire new_AGEMA_signal_12995 ;
    wire new_AGEMA_signal_12996 ;
    wire new_AGEMA_signal_12997 ;
    wire new_AGEMA_signal_12998 ;
    wire new_AGEMA_signal_12999 ;
    wire new_AGEMA_signal_13000 ;
    wire new_AGEMA_signal_13001 ;
    wire new_AGEMA_signal_13002 ;
    wire new_AGEMA_signal_13003 ;
    wire new_AGEMA_signal_13004 ;
    wire new_AGEMA_signal_13005 ;
    wire new_AGEMA_signal_13006 ;
    wire new_AGEMA_signal_13007 ;
    wire new_AGEMA_signal_13008 ;
    wire new_AGEMA_signal_13009 ;
    wire new_AGEMA_signal_13010 ;
    wire new_AGEMA_signal_13011 ;
    wire new_AGEMA_signal_13012 ;
    wire new_AGEMA_signal_13013 ;
    wire new_AGEMA_signal_13014 ;
    wire new_AGEMA_signal_13015 ;
    wire new_AGEMA_signal_13016 ;
    wire new_AGEMA_signal_13017 ;
    wire new_AGEMA_signal_13018 ;
    wire new_AGEMA_signal_13019 ;
    wire new_AGEMA_signal_13020 ;
    wire new_AGEMA_signal_13021 ;
    wire new_AGEMA_signal_13022 ;
    wire new_AGEMA_signal_13023 ;
    wire new_AGEMA_signal_13024 ;
    wire new_AGEMA_signal_13025 ;
    wire new_AGEMA_signal_13026 ;
    wire new_AGEMA_signal_13027 ;
    wire new_AGEMA_signal_13028 ;
    wire new_AGEMA_signal_13029 ;
    wire new_AGEMA_signal_13030 ;
    wire new_AGEMA_signal_13031 ;
    wire new_AGEMA_signal_13032 ;
    wire new_AGEMA_signal_13033 ;
    wire new_AGEMA_signal_13034 ;
    wire new_AGEMA_signal_13035 ;
    wire new_AGEMA_signal_13036 ;
    wire new_AGEMA_signal_13037 ;
    wire new_AGEMA_signal_13038 ;
    wire new_AGEMA_signal_13039 ;
    wire new_AGEMA_signal_13040 ;
    wire new_AGEMA_signal_13041 ;
    wire new_AGEMA_signal_13042 ;
    wire new_AGEMA_signal_13043 ;
    wire new_AGEMA_signal_13044 ;
    wire new_AGEMA_signal_13045 ;
    wire new_AGEMA_signal_13046 ;
    wire new_AGEMA_signal_13047 ;
    wire new_AGEMA_signal_13048 ;
    wire new_AGEMA_signal_13049 ;
    wire new_AGEMA_signal_13050 ;
    wire new_AGEMA_signal_13051 ;
    wire new_AGEMA_signal_13052 ;
    wire new_AGEMA_signal_13053 ;
    wire new_AGEMA_signal_13054 ;
    wire new_AGEMA_signal_13055 ;
    wire new_AGEMA_signal_13056 ;
    wire new_AGEMA_signal_13057 ;
    wire new_AGEMA_signal_13058 ;
    wire new_AGEMA_signal_13059 ;
    wire new_AGEMA_signal_13060 ;
    wire new_AGEMA_signal_13061 ;
    wire new_AGEMA_signal_13062 ;
    wire new_AGEMA_signal_13063 ;
    wire new_AGEMA_signal_13064 ;
    wire new_AGEMA_signal_13065 ;
    wire new_AGEMA_signal_13066 ;
    wire new_AGEMA_signal_13067 ;
    wire new_AGEMA_signal_13068 ;
    wire new_AGEMA_signal_13069 ;
    wire new_AGEMA_signal_13070 ;
    wire new_AGEMA_signal_13071 ;
    wire new_AGEMA_signal_13072 ;
    wire new_AGEMA_signal_13073 ;
    wire new_AGEMA_signal_13074 ;
    wire new_AGEMA_signal_13075 ;
    wire new_AGEMA_signal_13076 ;
    wire new_AGEMA_signal_13077 ;
    wire new_AGEMA_signal_13078 ;
    wire new_AGEMA_signal_13079 ;
    wire new_AGEMA_signal_13080 ;
    wire new_AGEMA_signal_13081 ;
    wire new_AGEMA_signal_13082 ;
    wire new_AGEMA_signal_13083 ;
    wire new_AGEMA_signal_13084 ;
    wire new_AGEMA_signal_13085 ;
    wire new_AGEMA_signal_13086 ;
    wire new_AGEMA_signal_13087 ;
    wire new_AGEMA_signal_13088 ;
    wire new_AGEMA_signal_13089 ;
    wire new_AGEMA_signal_13090 ;
    wire new_AGEMA_signal_13091 ;
    wire new_AGEMA_signal_13092 ;
    wire new_AGEMA_signal_13093 ;
    wire new_AGEMA_signal_13094 ;
    wire new_AGEMA_signal_13095 ;
    wire new_AGEMA_signal_13096 ;
    wire new_AGEMA_signal_13097 ;
    wire new_AGEMA_signal_13098 ;
    wire new_AGEMA_signal_13099 ;
    wire new_AGEMA_signal_13100 ;
    wire new_AGEMA_signal_13101 ;
    wire new_AGEMA_signal_13102 ;
    wire new_AGEMA_signal_13103 ;
    wire new_AGEMA_signal_13104 ;
    wire new_AGEMA_signal_13105 ;
    wire new_AGEMA_signal_13106 ;
    wire new_AGEMA_signal_13107 ;
    wire new_AGEMA_signal_13108 ;
    wire new_AGEMA_signal_13109 ;
    wire new_AGEMA_signal_13110 ;
    wire new_AGEMA_signal_13111 ;
    wire new_AGEMA_signal_13112 ;
    wire new_AGEMA_signal_13113 ;
    wire new_AGEMA_signal_13114 ;
    wire new_AGEMA_signal_13115 ;
    wire new_AGEMA_signal_13116 ;
    wire new_AGEMA_signal_13117 ;
    wire new_AGEMA_signal_13118 ;
    wire new_AGEMA_signal_13119 ;
    wire new_AGEMA_signal_13120 ;
    wire new_AGEMA_signal_13121 ;
    wire new_AGEMA_signal_13122 ;
    wire new_AGEMA_signal_13123 ;
    wire new_AGEMA_signal_13124 ;
    wire new_AGEMA_signal_13125 ;
    wire new_AGEMA_signal_13126 ;
    wire new_AGEMA_signal_13127 ;
    wire new_AGEMA_signal_13128 ;
    wire new_AGEMA_signal_13129 ;
    wire new_AGEMA_signal_13130 ;
    wire new_AGEMA_signal_13131 ;
    wire new_AGEMA_signal_13132 ;
    wire new_AGEMA_signal_13133 ;
    wire new_AGEMA_signal_13134 ;
    wire new_AGEMA_signal_13135 ;
    wire new_AGEMA_signal_13136 ;
    wire new_AGEMA_signal_13137 ;
    wire new_AGEMA_signal_13138 ;
    wire new_AGEMA_signal_13139 ;
    wire new_AGEMA_signal_13140 ;
    wire new_AGEMA_signal_13141 ;
    wire new_AGEMA_signal_13142 ;
    wire new_AGEMA_signal_13143 ;
    wire new_AGEMA_signal_13144 ;
    wire new_AGEMA_signal_13145 ;
    wire new_AGEMA_signal_13146 ;
    wire new_AGEMA_signal_13147 ;
    wire new_AGEMA_signal_13148 ;
    wire new_AGEMA_signal_13149 ;
    wire new_AGEMA_signal_13150 ;
    wire new_AGEMA_signal_13151 ;
    wire new_AGEMA_signal_13152 ;
    wire new_AGEMA_signal_13153 ;
    wire new_AGEMA_signal_13154 ;
    wire new_AGEMA_signal_13155 ;
    wire new_AGEMA_signal_13156 ;
    wire new_AGEMA_signal_13157 ;
    wire new_AGEMA_signal_13158 ;
    wire new_AGEMA_signal_13159 ;
    wire new_AGEMA_signal_13160 ;
    wire new_AGEMA_signal_13161 ;
    wire new_AGEMA_signal_13162 ;
    wire new_AGEMA_signal_13163 ;
    wire new_AGEMA_signal_13164 ;
    wire new_AGEMA_signal_13165 ;
    wire new_AGEMA_signal_13166 ;
    wire new_AGEMA_signal_13167 ;
    wire new_AGEMA_signal_13168 ;
    wire new_AGEMA_signal_13169 ;
    wire new_AGEMA_signal_13170 ;
    wire new_AGEMA_signal_13171 ;
    wire new_AGEMA_signal_13172 ;
    wire new_AGEMA_signal_13173 ;
    wire new_AGEMA_signal_13174 ;
    wire new_AGEMA_signal_13175 ;
    wire new_AGEMA_signal_13176 ;
    wire new_AGEMA_signal_13177 ;
    wire new_AGEMA_signal_13178 ;
    wire new_AGEMA_signal_13179 ;
    wire new_AGEMA_signal_13180 ;
    wire new_AGEMA_signal_13181 ;
    wire new_AGEMA_signal_13182 ;
    wire new_AGEMA_signal_13183 ;
    wire new_AGEMA_signal_13184 ;
    wire new_AGEMA_signal_13185 ;
    wire new_AGEMA_signal_13186 ;
    wire new_AGEMA_signal_13187 ;
    wire new_AGEMA_signal_13188 ;
    wire new_AGEMA_signal_13189 ;
    wire new_AGEMA_signal_13190 ;
    wire new_AGEMA_signal_13191 ;
    wire new_AGEMA_signal_13192 ;
    wire new_AGEMA_signal_13193 ;
    wire new_AGEMA_signal_13194 ;
    wire new_AGEMA_signal_13195 ;
    wire new_AGEMA_signal_13196 ;
    wire new_AGEMA_signal_13197 ;
    wire new_AGEMA_signal_13198 ;
    wire new_AGEMA_signal_13199 ;
    wire new_AGEMA_signal_13200 ;
    wire new_AGEMA_signal_13201 ;
    wire new_AGEMA_signal_13202 ;
    wire new_AGEMA_signal_13203 ;
    wire new_AGEMA_signal_13204 ;
    wire new_AGEMA_signal_13205 ;
    wire new_AGEMA_signal_13206 ;
    wire new_AGEMA_signal_13207 ;
    wire new_AGEMA_signal_13208 ;
    wire new_AGEMA_signal_13209 ;
    wire new_AGEMA_signal_13210 ;
    wire new_AGEMA_signal_13211 ;
    wire new_AGEMA_signal_13212 ;
    wire new_AGEMA_signal_13213 ;
    wire new_AGEMA_signal_13214 ;
    wire new_AGEMA_signal_13215 ;
    wire new_AGEMA_signal_13216 ;
    wire new_AGEMA_signal_13217 ;
    wire new_AGEMA_signal_13218 ;
    wire new_AGEMA_signal_13219 ;
    wire new_AGEMA_signal_13220 ;
    wire new_AGEMA_signal_13221 ;
    wire new_AGEMA_signal_13222 ;
    wire new_AGEMA_signal_13223 ;
    wire new_AGEMA_signal_13224 ;
    wire new_AGEMA_signal_13225 ;
    wire new_AGEMA_signal_13226 ;
    wire new_AGEMA_signal_13227 ;
    wire new_AGEMA_signal_13228 ;
    wire new_AGEMA_signal_13229 ;
    wire new_AGEMA_signal_13230 ;
    wire new_AGEMA_signal_13231 ;
    wire new_AGEMA_signal_13232 ;
    wire new_AGEMA_signal_13233 ;
    wire new_AGEMA_signal_13234 ;
    wire new_AGEMA_signal_13235 ;
    wire new_AGEMA_signal_13236 ;
    wire new_AGEMA_signal_13237 ;
    wire new_AGEMA_signal_13238 ;
    wire new_AGEMA_signal_13239 ;
    wire new_AGEMA_signal_13240 ;
    wire new_AGEMA_signal_13241 ;
    wire new_AGEMA_signal_13242 ;
    wire new_AGEMA_signal_13243 ;
    wire new_AGEMA_signal_13244 ;
    wire new_AGEMA_signal_13245 ;
    wire new_AGEMA_signal_13246 ;
    wire new_AGEMA_signal_13247 ;
    wire new_AGEMA_signal_13248 ;
    wire new_AGEMA_signal_13249 ;
    wire new_AGEMA_signal_13250 ;
    wire new_AGEMA_signal_13251 ;
    wire new_AGEMA_signal_13252 ;
    wire new_AGEMA_signal_13253 ;
    wire new_AGEMA_signal_13254 ;
    wire new_AGEMA_signal_13255 ;
    wire new_AGEMA_signal_13256 ;
    wire new_AGEMA_signal_13257 ;
    wire new_AGEMA_signal_13258 ;
    wire new_AGEMA_signal_13259 ;
    wire new_AGEMA_signal_13260 ;
    wire new_AGEMA_signal_13261 ;
    wire new_AGEMA_signal_13262 ;
    wire new_AGEMA_signal_13263 ;
    wire new_AGEMA_signal_13264 ;
    wire new_AGEMA_signal_13265 ;
    wire new_AGEMA_signal_13266 ;
    wire new_AGEMA_signal_13267 ;
    wire new_AGEMA_signal_13268 ;
    wire new_AGEMA_signal_13269 ;
    wire new_AGEMA_signal_13270 ;
    wire new_AGEMA_signal_13271 ;
    wire new_AGEMA_signal_13272 ;
    wire new_AGEMA_signal_13273 ;
    wire new_AGEMA_signal_13274 ;
    wire new_AGEMA_signal_13275 ;
    wire new_AGEMA_signal_13276 ;
    wire new_AGEMA_signal_13277 ;
    wire new_AGEMA_signal_13278 ;
    wire new_AGEMA_signal_13279 ;
    wire new_AGEMA_signal_13280 ;
    wire new_AGEMA_signal_13281 ;
    wire new_AGEMA_signal_13282 ;
    wire new_AGEMA_signal_13283 ;
    wire new_AGEMA_signal_13284 ;
    wire new_AGEMA_signal_13285 ;
    wire new_AGEMA_signal_13286 ;
    wire new_AGEMA_signal_13287 ;
    wire new_AGEMA_signal_13288 ;
    wire new_AGEMA_signal_13289 ;
    wire new_AGEMA_signal_13290 ;
    wire new_AGEMA_signal_13291 ;
    wire new_AGEMA_signal_13292 ;
    wire new_AGEMA_signal_13293 ;
    wire new_AGEMA_signal_13294 ;
    wire new_AGEMA_signal_13295 ;
    wire new_AGEMA_signal_13296 ;
    wire new_AGEMA_signal_13297 ;
    wire new_AGEMA_signal_13298 ;
    wire new_AGEMA_signal_13299 ;
    wire new_AGEMA_signal_13300 ;
    wire new_AGEMA_signal_13301 ;
    wire new_AGEMA_signal_13302 ;
    wire new_AGEMA_signal_13303 ;
    wire new_AGEMA_signal_13304 ;
    wire new_AGEMA_signal_13305 ;
    wire new_AGEMA_signal_13306 ;
    wire new_AGEMA_signal_13307 ;
    wire new_AGEMA_signal_13308 ;
    wire new_AGEMA_signal_13309 ;
    wire new_AGEMA_signal_13310 ;
    wire new_AGEMA_signal_13311 ;
    wire new_AGEMA_signal_13312 ;
    wire new_AGEMA_signal_13313 ;
    wire new_AGEMA_signal_13314 ;
    wire new_AGEMA_signal_13315 ;
    wire new_AGEMA_signal_13316 ;
    wire new_AGEMA_signal_13317 ;
    wire new_AGEMA_signal_13318 ;
    wire new_AGEMA_signal_13319 ;
    wire new_AGEMA_signal_13320 ;
    wire new_AGEMA_signal_13321 ;
    wire new_AGEMA_signal_13322 ;
    wire new_AGEMA_signal_13323 ;
    wire new_AGEMA_signal_13324 ;
    wire new_AGEMA_signal_13325 ;
    wire new_AGEMA_signal_13326 ;
    wire new_AGEMA_signal_13327 ;
    wire new_AGEMA_signal_13328 ;
    wire new_AGEMA_signal_13329 ;
    wire new_AGEMA_signal_13330 ;
    wire new_AGEMA_signal_13331 ;
    wire new_AGEMA_signal_13332 ;
    wire new_AGEMA_signal_13333 ;
    wire new_AGEMA_signal_13334 ;
    wire new_AGEMA_signal_13335 ;
    wire new_AGEMA_signal_13336 ;
    wire new_AGEMA_signal_13337 ;
    wire new_AGEMA_signal_13338 ;
    wire new_AGEMA_signal_13339 ;
    wire new_AGEMA_signal_13340 ;
    wire new_AGEMA_signal_13341 ;
    wire new_AGEMA_signal_13342 ;
    wire new_AGEMA_signal_13343 ;
    wire new_AGEMA_signal_13344 ;
    wire new_AGEMA_signal_13345 ;
    wire new_AGEMA_signal_13346 ;
    wire new_AGEMA_signal_13347 ;
    wire new_AGEMA_signal_13348 ;
    wire new_AGEMA_signal_13349 ;
    wire new_AGEMA_signal_13350 ;
    wire new_AGEMA_signal_13351 ;
    wire new_AGEMA_signal_13352 ;
    wire new_AGEMA_signal_13353 ;
    wire new_AGEMA_signal_13354 ;
    wire new_AGEMA_signal_13355 ;
    wire new_AGEMA_signal_13356 ;
    wire new_AGEMA_signal_13357 ;
    wire new_AGEMA_signal_13358 ;
    wire new_AGEMA_signal_13359 ;
    wire new_AGEMA_signal_13360 ;
    wire new_AGEMA_signal_13361 ;
    wire new_AGEMA_signal_13362 ;
    wire new_AGEMA_signal_13363 ;
    wire new_AGEMA_signal_13364 ;
    wire new_AGEMA_signal_13365 ;
    wire new_AGEMA_signal_13366 ;
    wire new_AGEMA_signal_13367 ;
    wire new_AGEMA_signal_13368 ;
    wire new_AGEMA_signal_13369 ;
    wire new_AGEMA_signal_13370 ;
    wire new_AGEMA_signal_13371 ;
    wire new_AGEMA_signal_13372 ;
    wire new_AGEMA_signal_13373 ;
    wire new_AGEMA_signal_13374 ;
    wire new_AGEMA_signal_13375 ;
    wire new_AGEMA_signal_13376 ;
    wire new_AGEMA_signal_13377 ;
    wire new_AGEMA_signal_13378 ;
    wire new_AGEMA_signal_13379 ;
    wire new_AGEMA_signal_13380 ;
    wire new_AGEMA_signal_13381 ;
    wire new_AGEMA_signal_13382 ;
    wire new_AGEMA_signal_13383 ;
    wire new_AGEMA_signal_13384 ;
    wire new_AGEMA_signal_13385 ;
    wire new_AGEMA_signal_13386 ;
    wire new_AGEMA_signal_13387 ;
    wire new_AGEMA_signal_13388 ;
    wire new_AGEMA_signal_13389 ;
    wire new_AGEMA_signal_13390 ;
    wire new_AGEMA_signal_13391 ;
    wire new_AGEMA_signal_13392 ;
    wire new_AGEMA_signal_13393 ;
    wire new_AGEMA_signal_13394 ;
    wire new_AGEMA_signal_13395 ;
    wire new_AGEMA_signal_13396 ;
    wire new_AGEMA_signal_13397 ;
    wire new_AGEMA_signal_13398 ;
    wire new_AGEMA_signal_13399 ;
    wire new_AGEMA_signal_13400 ;
    wire new_AGEMA_signal_13401 ;
    wire new_AGEMA_signal_13402 ;
    wire new_AGEMA_signal_13403 ;
    wire new_AGEMA_signal_13404 ;
    wire new_AGEMA_signal_13405 ;
    wire new_AGEMA_signal_13406 ;
    wire new_AGEMA_signal_13407 ;
    wire new_AGEMA_signal_13408 ;
    wire new_AGEMA_signal_13409 ;
    wire new_AGEMA_signal_13410 ;
    wire new_AGEMA_signal_13411 ;
    wire new_AGEMA_signal_13412 ;
    wire new_AGEMA_signal_13413 ;
    wire new_AGEMA_signal_13414 ;
    wire new_AGEMA_signal_13415 ;
    wire new_AGEMA_signal_13416 ;
    wire new_AGEMA_signal_13417 ;
    wire new_AGEMA_signal_13418 ;
    wire new_AGEMA_signal_13419 ;
    wire new_AGEMA_signal_13420 ;
    wire new_AGEMA_signal_13421 ;
    wire new_AGEMA_signal_13422 ;
    wire new_AGEMA_signal_13423 ;
    wire new_AGEMA_signal_13424 ;
    wire new_AGEMA_signal_13425 ;
    wire new_AGEMA_signal_13426 ;
    wire new_AGEMA_signal_13427 ;
    wire new_AGEMA_signal_13428 ;
    wire new_AGEMA_signal_13429 ;
    wire new_AGEMA_signal_13430 ;
    wire new_AGEMA_signal_13431 ;
    wire new_AGEMA_signal_13432 ;
    wire new_AGEMA_signal_13433 ;
    wire new_AGEMA_signal_13434 ;
    wire new_AGEMA_signal_13435 ;
    wire new_AGEMA_signal_13436 ;
    wire new_AGEMA_signal_13437 ;
    wire new_AGEMA_signal_13438 ;
    wire new_AGEMA_signal_13439 ;
    wire new_AGEMA_signal_13440 ;
    wire new_AGEMA_signal_13441 ;
    wire new_AGEMA_signal_13442 ;
    wire new_AGEMA_signal_13443 ;
    wire new_AGEMA_signal_13444 ;
    wire new_AGEMA_signal_13445 ;
    wire new_AGEMA_signal_13446 ;
    wire new_AGEMA_signal_13447 ;
    wire new_AGEMA_signal_13448 ;
    wire new_AGEMA_signal_13449 ;
    wire new_AGEMA_signal_13450 ;
    wire new_AGEMA_signal_13451 ;
    wire new_AGEMA_signal_13452 ;
    wire new_AGEMA_signal_13453 ;
    wire new_AGEMA_signal_13454 ;
    wire new_AGEMA_signal_13455 ;
    wire new_AGEMA_signal_13456 ;
    wire new_AGEMA_signal_13457 ;
    wire new_AGEMA_signal_13458 ;
    wire new_AGEMA_signal_13459 ;
    wire new_AGEMA_signal_13460 ;
    wire new_AGEMA_signal_13461 ;
    wire new_AGEMA_signal_13462 ;
    wire new_AGEMA_signal_13463 ;
    wire new_AGEMA_signal_13464 ;
    wire new_AGEMA_signal_13465 ;
    wire new_AGEMA_signal_13466 ;
    wire new_AGEMA_signal_13467 ;
    wire new_AGEMA_signal_13468 ;
    wire new_AGEMA_signal_13469 ;
    wire new_AGEMA_signal_13470 ;
    wire new_AGEMA_signal_13471 ;
    wire new_AGEMA_signal_13472 ;
    wire new_AGEMA_signal_13473 ;
    wire new_AGEMA_signal_13474 ;
    wire new_AGEMA_signal_13475 ;
    wire new_AGEMA_signal_13476 ;
    wire new_AGEMA_signal_13477 ;
    wire new_AGEMA_signal_13478 ;
    wire new_AGEMA_signal_13479 ;
    wire new_AGEMA_signal_13480 ;
    wire new_AGEMA_signal_13481 ;
    wire new_AGEMA_signal_13482 ;
    wire new_AGEMA_signal_13483 ;
    wire new_AGEMA_signal_13484 ;
    wire new_AGEMA_signal_13485 ;
    wire new_AGEMA_signal_13486 ;
    wire new_AGEMA_signal_13487 ;
    wire new_AGEMA_signal_13488 ;
    wire new_AGEMA_signal_13489 ;
    wire new_AGEMA_signal_13490 ;
    wire new_AGEMA_signal_13491 ;
    wire new_AGEMA_signal_13492 ;
    wire new_AGEMA_signal_13493 ;
    wire new_AGEMA_signal_13494 ;
    wire new_AGEMA_signal_13495 ;
    wire new_AGEMA_signal_13496 ;
    wire new_AGEMA_signal_13497 ;
    wire new_AGEMA_signal_13498 ;
    wire new_AGEMA_signal_13499 ;
    wire new_AGEMA_signal_13500 ;
    wire new_AGEMA_signal_13501 ;
    wire new_AGEMA_signal_13502 ;
    wire new_AGEMA_signal_13503 ;
    wire new_AGEMA_signal_13504 ;
    wire new_AGEMA_signal_13505 ;
    wire new_AGEMA_signal_13506 ;
    wire new_AGEMA_signal_13507 ;
    wire new_AGEMA_signal_13508 ;
    wire new_AGEMA_signal_13509 ;
    wire new_AGEMA_signal_13510 ;
    wire new_AGEMA_signal_13511 ;
    wire new_AGEMA_signal_13512 ;
    wire new_AGEMA_signal_13513 ;
    wire new_AGEMA_signal_13514 ;
    wire new_AGEMA_signal_13515 ;
    wire new_AGEMA_signal_13516 ;
    wire new_AGEMA_signal_13517 ;
    wire new_AGEMA_signal_13518 ;
    wire new_AGEMA_signal_13519 ;
    wire new_AGEMA_signal_13520 ;
    wire new_AGEMA_signal_13521 ;
    wire new_AGEMA_signal_13522 ;
    wire new_AGEMA_signal_13523 ;
    wire new_AGEMA_signal_13524 ;
    wire new_AGEMA_signal_13525 ;
    wire new_AGEMA_signal_13526 ;
    wire new_AGEMA_signal_13527 ;
    wire new_AGEMA_signal_13528 ;
    wire new_AGEMA_signal_13529 ;
    wire new_AGEMA_signal_13530 ;
    wire new_AGEMA_signal_13531 ;
    wire new_AGEMA_signal_13532 ;
    wire new_AGEMA_signal_13533 ;
    wire new_AGEMA_signal_13534 ;
    wire new_AGEMA_signal_13535 ;
    wire new_AGEMA_signal_13536 ;
    wire new_AGEMA_signal_13537 ;
    wire new_AGEMA_signal_13538 ;
    wire new_AGEMA_signal_13539 ;
    wire new_AGEMA_signal_13540 ;
    wire new_AGEMA_signal_13541 ;
    wire new_AGEMA_signal_13542 ;
    wire new_AGEMA_signal_13543 ;
    wire new_AGEMA_signal_13544 ;
    wire new_AGEMA_signal_13545 ;
    wire new_AGEMA_signal_13546 ;
    wire new_AGEMA_signal_13547 ;
    wire new_AGEMA_signal_13548 ;
    wire new_AGEMA_signal_13549 ;
    wire new_AGEMA_signal_13550 ;
    wire new_AGEMA_signal_13551 ;
    wire new_AGEMA_signal_13552 ;
    wire new_AGEMA_signal_13553 ;
    wire new_AGEMA_signal_13554 ;
    wire new_AGEMA_signal_13555 ;
    wire new_AGEMA_signal_13556 ;
    wire new_AGEMA_signal_13557 ;
    wire new_AGEMA_signal_13558 ;
    wire new_AGEMA_signal_13559 ;
    wire new_AGEMA_signal_13560 ;
    wire new_AGEMA_signal_13561 ;
    wire new_AGEMA_signal_13562 ;
    wire new_AGEMA_signal_13563 ;
    wire new_AGEMA_signal_13564 ;
    wire new_AGEMA_signal_13565 ;
    wire new_AGEMA_signal_13566 ;
    wire new_AGEMA_signal_13567 ;
    wire new_AGEMA_signal_13568 ;
    wire new_AGEMA_signal_13569 ;
    wire new_AGEMA_signal_13570 ;
    wire new_AGEMA_signal_13571 ;
    wire new_AGEMA_signal_13572 ;
    wire new_AGEMA_signal_13573 ;
    wire new_AGEMA_signal_13574 ;
    wire new_AGEMA_signal_13575 ;
    wire new_AGEMA_signal_13576 ;
    wire new_AGEMA_signal_13577 ;
    wire new_AGEMA_signal_13578 ;
    wire new_AGEMA_signal_13579 ;
    wire new_AGEMA_signal_13580 ;
    wire new_AGEMA_signal_13581 ;
    wire new_AGEMA_signal_13582 ;
    wire new_AGEMA_signal_13583 ;
    wire new_AGEMA_signal_13584 ;
    wire new_AGEMA_signal_13585 ;
    wire new_AGEMA_signal_13586 ;
    wire new_AGEMA_signal_13587 ;
    wire new_AGEMA_signal_13588 ;
    wire new_AGEMA_signal_13589 ;
    wire new_AGEMA_signal_13590 ;
    wire new_AGEMA_signal_13591 ;
    wire new_AGEMA_signal_13592 ;
    wire new_AGEMA_signal_13593 ;
    wire new_AGEMA_signal_13594 ;
    wire new_AGEMA_signal_13595 ;
    wire new_AGEMA_signal_13596 ;
    wire new_AGEMA_signal_13597 ;
    wire new_AGEMA_signal_13598 ;
    wire new_AGEMA_signal_13599 ;
    wire new_AGEMA_signal_13600 ;
    wire new_AGEMA_signal_13601 ;
    wire new_AGEMA_signal_13602 ;
    wire new_AGEMA_signal_13603 ;
    wire new_AGEMA_signal_13604 ;
    wire new_AGEMA_signal_13605 ;
    wire new_AGEMA_signal_13606 ;
    wire new_AGEMA_signal_13607 ;
    wire new_AGEMA_signal_13608 ;
    wire new_AGEMA_signal_13609 ;
    wire new_AGEMA_signal_13610 ;
    wire new_AGEMA_signal_13611 ;
    wire new_AGEMA_signal_13612 ;
    wire new_AGEMA_signal_13613 ;
    wire new_AGEMA_signal_13614 ;
    wire new_AGEMA_signal_13615 ;
    wire new_AGEMA_signal_13616 ;
    wire new_AGEMA_signal_13617 ;
    wire new_AGEMA_signal_13618 ;
    wire new_AGEMA_signal_13619 ;
    wire new_AGEMA_signal_13620 ;
    wire new_AGEMA_signal_13621 ;
    wire new_AGEMA_signal_13622 ;
    wire new_AGEMA_signal_13623 ;
    wire new_AGEMA_signal_13624 ;
    wire new_AGEMA_signal_13625 ;
    wire new_AGEMA_signal_13626 ;
    wire new_AGEMA_signal_13627 ;
    wire new_AGEMA_signal_13628 ;
    wire new_AGEMA_signal_13629 ;
    wire new_AGEMA_signal_13630 ;
    wire new_AGEMA_signal_13631 ;
    wire new_AGEMA_signal_13632 ;
    wire new_AGEMA_signal_13633 ;
    wire new_AGEMA_signal_13634 ;
    wire new_AGEMA_signal_13635 ;
    wire new_AGEMA_signal_13636 ;
    wire new_AGEMA_signal_13637 ;
    wire new_AGEMA_signal_13638 ;
    wire new_AGEMA_signal_13639 ;
    wire new_AGEMA_signal_13640 ;
    wire new_AGEMA_signal_13641 ;
    wire new_AGEMA_signal_13642 ;
    wire new_AGEMA_signal_13643 ;
    wire new_AGEMA_signal_13644 ;
    wire new_AGEMA_signal_13645 ;
    wire new_AGEMA_signal_13646 ;
    wire new_AGEMA_signal_13647 ;
    wire new_AGEMA_signal_13648 ;
    wire new_AGEMA_signal_13649 ;
    wire new_AGEMA_signal_13650 ;
    wire new_AGEMA_signal_13651 ;
    wire new_AGEMA_signal_13652 ;
    wire new_AGEMA_signal_13653 ;
    wire new_AGEMA_signal_13654 ;
    wire new_AGEMA_signal_13655 ;
    wire new_AGEMA_signal_13656 ;
    wire new_AGEMA_signal_13657 ;
    wire new_AGEMA_signal_13658 ;
    wire new_AGEMA_signal_13659 ;
    wire new_AGEMA_signal_13660 ;
    wire new_AGEMA_signal_13661 ;
    wire new_AGEMA_signal_13662 ;
    wire new_AGEMA_signal_13663 ;
    wire new_AGEMA_signal_13664 ;
    wire new_AGEMA_signal_13665 ;
    wire new_AGEMA_signal_13666 ;
    wire new_AGEMA_signal_13667 ;
    wire new_AGEMA_signal_13668 ;
    wire new_AGEMA_signal_13669 ;
    wire new_AGEMA_signal_13670 ;
    wire new_AGEMA_signal_13671 ;
    wire new_AGEMA_signal_13672 ;
    wire new_AGEMA_signal_13673 ;
    wire new_AGEMA_signal_13674 ;
    wire new_AGEMA_signal_13675 ;
    wire new_AGEMA_signal_13676 ;
    wire new_AGEMA_signal_13677 ;
    wire new_AGEMA_signal_13678 ;
    wire new_AGEMA_signal_13679 ;
    wire new_AGEMA_signal_13680 ;
    wire new_AGEMA_signal_13681 ;
    wire new_AGEMA_signal_13682 ;
    wire new_AGEMA_signal_13683 ;
    wire new_AGEMA_signal_13684 ;
    wire new_AGEMA_signal_13685 ;
    wire new_AGEMA_signal_13686 ;
    wire new_AGEMA_signal_13687 ;
    wire new_AGEMA_signal_13688 ;
    wire new_AGEMA_signal_13689 ;
    wire new_AGEMA_signal_13690 ;
    wire new_AGEMA_signal_13691 ;
    wire new_AGEMA_signal_13692 ;
    wire new_AGEMA_signal_13693 ;
    wire new_AGEMA_signal_13694 ;
    wire new_AGEMA_signal_13695 ;
    wire new_AGEMA_signal_13696 ;
    wire new_AGEMA_signal_13697 ;
    wire new_AGEMA_signal_13698 ;
    wire new_AGEMA_signal_13699 ;
    wire new_AGEMA_signal_13700 ;
    wire new_AGEMA_signal_13701 ;
    wire new_AGEMA_signal_13702 ;
    wire new_AGEMA_signal_13703 ;
    wire new_AGEMA_signal_13704 ;
    wire new_AGEMA_signal_13705 ;
    wire new_AGEMA_signal_13706 ;
    wire new_AGEMA_signal_13707 ;
    wire new_AGEMA_signal_13708 ;
    wire new_AGEMA_signal_13709 ;
    wire new_AGEMA_signal_13710 ;
    wire new_AGEMA_signal_13711 ;
    wire new_AGEMA_signal_13712 ;
    wire new_AGEMA_signal_13713 ;
    wire new_AGEMA_signal_13714 ;
    wire new_AGEMA_signal_13715 ;
    wire new_AGEMA_signal_13716 ;
    wire new_AGEMA_signal_13717 ;
    wire new_AGEMA_signal_13718 ;
    wire new_AGEMA_signal_13719 ;
    wire new_AGEMA_signal_13720 ;
    wire new_AGEMA_signal_13721 ;
    wire new_AGEMA_signal_13722 ;
    wire new_AGEMA_signal_13723 ;
    wire new_AGEMA_signal_13724 ;
    wire new_AGEMA_signal_13725 ;
    wire new_AGEMA_signal_13726 ;
    wire new_AGEMA_signal_13727 ;
    wire new_AGEMA_signal_13728 ;
    wire new_AGEMA_signal_13729 ;
    wire new_AGEMA_signal_13730 ;
    wire new_AGEMA_signal_13731 ;
    wire new_AGEMA_signal_13732 ;
    wire new_AGEMA_signal_13733 ;
    wire new_AGEMA_signal_13734 ;
    wire new_AGEMA_signal_13735 ;
    wire new_AGEMA_signal_13736 ;
    wire new_AGEMA_signal_13737 ;
    wire new_AGEMA_signal_13738 ;
    wire new_AGEMA_signal_13739 ;
    wire new_AGEMA_signal_13740 ;
    wire new_AGEMA_signal_13741 ;
    wire new_AGEMA_signal_13742 ;
    wire new_AGEMA_signal_13743 ;
    wire new_AGEMA_signal_13744 ;
    wire new_AGEMA_signal_13745 ;
    wire new_AGEMA_signal_13746 ;
    wire new_AGEMA_signal_13747 ;
    wire new_AGEMA_signal_13748 ;
    wire new_AGEMA_signal_13749 ;
    wire new_AGEMA_signal_13750 ;
    wire new_AGEMA_signal_13751 ;
    wire new_AGEMA_signal_13752 ;
    wire new_AGEMA_signal_13753 ;
    wire new_AGEMA_signal_13754 ;
    wire new_AGEMA_signal_13755 ;
    wire new_AGEMA_signal_13756 ;
    wire new_AGEMA_signal_13757 ;
    wire new_AGEMA_signal_13758 ;
    wire new_AGEMA_signal_13759 ;
    wire new_AGEMA_signal_13760 ;
    wire new_AGEMA_signal_13761 ;
    wire new_AGEMA_signal_13762 ;
    wire new_AGEMA_signal_13763 ;
    wire new_AGEMA_signal_13764 ;
    wire new_AGEMA_signal_13765 ;
    wire new_AGEMA_signal_13766 ;
    wire new_AGEMA_signal_13767 ;
    wire new_AGEMA_signal_13768 ;
    wire new_AGEMA_signal_13769 ;
    wire new_AGEMA_signal_13770 ;
    wire new_AGEMA_signal_13771 ;
    wire new_AGEMA_signal_13772 ;
    wire new_AGEMA_signal_13773 ;
    wire new_AGEMA_signal_13774 ;
    wire new_AGEMA_signal_13775 ;
    wire new_AGEMA_signal_13776 ;
    wire new_AGEMA_signal_13777 ;
    wire new_AGEMA_signal_13778 ;
    wire new_AGEMA_signal_13779 ;
    wire new_AGEMA_signal_13780 ;
    wire new_AGEMA_signal_13781 ;
    wire new_AGEMA_signal_13782 ;
    wire new_AGEMA_signal_13783 ;
    wire new_AGEMA_signal_13784 ;
    wire new_AGEMA_signal_13785 ;
    wire new_AGEMA_signal_13786 ;
    wire new_AGEMA_signal_13787 ;
    wire new_AGEMA_signal_13788 ;
    wire new_AGEMA_signal_13789 ;
    wire new_AGEMA_signal_13790 ;
    wire new_AGEMA_signal_13791 ;
    wire new_AGEMA_signal_13792 ;
    wire new_AGEMA_signal_13793 ;
    wire new_AGEMA_signal_13794 ;
    wire new_AGEMA_signal_13795 ;
    wire new_AGEMA_signal_13796 ;
    wire new_AGEMA_signal_13797 ;
    wire new_AGEMA_signal_13798 ;
    wire new_AGEMA_signal_13799 ;
    wire new_AGEMA_signal_13800 ;
    wire new_AGEMA_signal_13801 ;
    wire new_AGEMA_signal_13802 ;
    wire new_AGEMA_signal_13803 ;
    wire new_AGEMA_signal_13804 ;
    wire new_AGEMA_signal_13805 ;
    wire new_AGEMA_signal_13806 ;
    wire new_AGEMA_signal_13807 ;
    wire new_AGEMA_signal_13808 ;
    wire new_AGEMA_signal_13809 ;
    wire new_AGEMA_signal_13810 ;
    wire new_AGEMA_signal_13811 ;
    wire new_AGEMA_signal_13812 ;
    wire new_AGEMA_signal_13813 ;
    wire new_AGEMA_signal_13814 ;
    wire new_AGEMA_signal_13815 ;
    wire new_AGEMA_signal_13816 ;
    wire new_AGEMA_signal_13817 ;
    wire new_AGEMA_signal_13818 ;
    wire new_AGEMA_signal_13819 ;
    wire new_AGEMA_signal_13820 ;
    wire new_AGEMA_signal_13821 ;
    wire new_AGEMA_signal_13822 ;
    wire new_AGEMA_signal_13823 ;
    wire new_AGEMA_signal_13824 ;
    wire new_AGEMA_signal_13825 ;
    wire new_AGEMA_signal_13826 ;
    wire new_AGEMA_signal_13827 ;
    wire new_AGEMA_signal_13828 ;
    wire new_AGEMA_signal_13829 ;
    wire new_AGEMA_signal_13830 ;
    wire new_AGEMA_signal_13831 ;
    wire new_AGEMA_signal_13832 ;
    wire new_AGEMA_signal_13833 ;
    wire new_AGEMA_signal_13834 ;
    wire new_AGEMA_signal_13835 ;
    wire new_AGEMA_signal_13836 ;
    wire new_AGEMA_signal_13837 ;
    wire new_AGEMA_signal_13838 ;
    wire new_AGEMA_signal_13839 ;
    wire new_AGEMA_signal_13840 ;
    wire new_AGEMA_signal_13841 ;
    wire new_AGEMA_signal_13842 ;
    wire new_AGEMA_signal_13843 ;
    wire new_AGEMA_signal_13844 ;
    wire new_AGEMA_signal_13845 ;
    wire new_AGEMA_signal_13846 ;
    wire new_AGEMA_signal_13847 ;
    wire new_AGEMA_signal_13848 ;
    wire new_AGEMA_signal_13849 ;
    wire new_AGEMA_signal_13850 ;
    wire new_AGEMA_signal_13851 ;
    wire new_AGEMA_signal_13852 ;
    wire new_AGEMA_signal_13853 ;
    wire new_AGEMA_signal_13854 ;
    wire new_AGEMA_signal_13855 ;
    wire new_AGEMA_signal_13856 ;
    wire new_AGEMA_signal_13857 ;
    wire new_AGEMA_signal_13858 ;
    wire new_AGEMA_signal_13859 ;
    wire new_AGEMA_signal_13860 ;
    wire new_AGEMA_signal_13861 ;
    wire new_AGEMA_signal_13862 ;
    wire new_AGEMA_signal_13863 ;
    wire new_AGEMA_signal_13864 ;
    wire new_AGEMA_signal_13865 ;
    wire new_AGEMA_signal_13866 ;
    wire new_AGEMA_signal_13867 ;
    wire new_AGEMA_signal_13868 ;
    wire new_AGEMA_signal_13869 ;
    wire new_AGEMA_signal_13870 ;
    wire new_AGEMA_signal_13871 ;
    wire new_AGEMA_signal_13872 ;
    wire new_AGEMA_signal_13873 ;
    wire new_AGEMA_signal_13874 ;
    wire new_AGEMA_signal_13875 ;
    wire new_AGEMA_signal_13876 ;
    wire new_AGEMA_signal_13877 ;
    wire new_AGEMA_signal_13878 ;
    wire new_AGEMA_signal_13879 ;
    wire new_AGEMA_signal_13880 ;
    wire new_AGEMA_signal_13881 ;
    wire new_AGEMA_signal_13882 ;
    wire new_AGEMA_signal_13883 ;
    wire new_AGEMA_signal_13884 ;
    wire new_AGEMA_signal_13885 ;
    wire new_AGEMA_signal_13886 ;
    wire new_AGEMA_signal_13887 ;
    wire new_AGEMA_signal_13888 ;
    wire new_AGEMA_signal_13889 ;
    wire new_AGEMA_signal_13890 ;
    wire new_AGEMA_signal_13891 ;
    wire new_AGEMA_signal_13892 ;
    wire new_AGEMA_signal_13893 ;
    wire new_AGEMA_signal_13894 ;
    wire new_AGEMA_signal_13895 ;
    wire new_AGEMA_signal_13896 ;
    wire new_AGEMA_signal_13897 ;
    wire new_AGEMA_signal_13898 ;
    wire new_AGEMA_signal_13899 ;
    wire new_AGEMA_signal_13900 ;
    wire new_AGEMA_signal_13901 ;
    wire new_AGEMA_signal_13902 ;
    wire new_AGEMA_signal_13903 ;
    wire new_AGEMA_signal_13904 ;
    wire new_AGEMA_signal_13905 ;
    wire new_AGEMA_signal_13906 ;
    wire new_AGEMA_signal_13907 ;
    wire new_AGEMA_signal_13908 ;
    wire new_AGEMA_signal_13909 ;
    wire new_AGEMA_signal_13910 ;
    wire new_AGEMA_signal_13911 ;
    wire new_AGEMA_signal_13912 ;
    wire new_AGEMA_signal_13913 ;
    wire new_AGEMA_signal_13914 ;
    wire new_AGEMA_signal_13915 ;
    wire new_AGEMA_signal_13916 ;
    wire new_AGEMA_signal_13917 ;
    wire new_AGEMA_signal_13918 ;
    wire new_AGEMA_signal_13919 ;
    wire new_AGEMA_signal_13920 ;
    wire new_AGEMA_signal_13921 ;
    wire new_AGEMA_signal_13922 ;
    wire new_AGEMA_signal_13923 ;
    wire new_AGEMA_signal_13924 ;
    wire new_AGEMA_signal_13925 ;
    wire new_AGEMA_signal_13926 ;
    wire new_AGEMA_signal_13927 ;
    wire new_AGEMA_signal_13928 ;
    wire new_AGEMA_signal_13929 ;
    wire new_AGEMA_signal_13930 ;
    wire new_AGEMA_signal_13931 ;
    wire new_AGEMA_signal_13932 ;
    wire new_AGEMA_signal_13933 ;
    wire new_AGEMA_signal_13934 ;
    wire new_AGEMA_signal_13935 ;
    wire new_AGEMA_signal_13936 ;
    wire new_AGEMA_signal_13937 ;
    wire new_AGEMA_signal_13938 ;
    wire new_AGEMA_signal_13939 ;
    wire new_AGEMA_signal_13940 ;
    wire new_AGEMA_signal_13941 ;
    wire new_AGEMA_signal_13942 ;
    wire new_AGEMA_signal_13943 ;
    wire new_AGEMA_signal_13944 ;
    wire new_AGEMA_signal_13945 ;
    wire new_AGEMA_signal_13946 ;
    wire new_AGEMA_signal_13947 ;
    wire new_AGEMA_signal_13948 ;
    wire new_AGEMA_signal_13949 ;
    wire new_AGEMA_signal_13950 ;
    wire new_AGEMA_signal_13951 ;
    wire new_AGEMA_signal_13952 ;
    wire new_AGEMA_signal_13953 ;
    wire new_AGEMA_signal_13954 ;
    wire new_AGEMA_signal_13955 ;
    wire new_AGEMA_signal_13956 ;
    wire new_AGEMA_signal_13957 ;
    wire new_AGEMA_signal_13958 ;
    wire new_AGEMA_signal_13959 ;
    wire new_AGEMA_signal_13960 ;
    wire new_AGEMA_signal_13961 ;
    wire new_AGEMA_signal_13962 ;
    wire new_AGEMA_signal_13963 ;
    wire new_AGEMA_signal_13964 ;
    wire new_AGEMA_signal_13965 ;
    wire new_AGEMA_signal_13966 ;
    wire new_AGEMA_signal_13967 ;
    wire new_AGEMA_signal_13968 ;
    wire new_AGEMA_signal_13969 ;
    wire new_AGEMA_signal_13970 ;
    wire new_AGEMA_signal_13971 ;
    wire new_AGEMA_signal_13972 ;
    wire new_AGEMA_signal_13973 ;
    wire new_AGEMA_signal_13974 ;
    wire new_AGEMA_signal_13975 ;
    wire new_AGEMA_signal_13979 ;
    wire new_AGEMA_signal_13980 ;
    wire new_AGEMA_signal_13981 ;
    wire new_AGEMA_signal_13985 ;
    wire new_AGEMA_signal_13986 ;
    wire new_AGEMA_signal_13987 ;
    wire new_AGEMA_signal_13991 ;
    wire new_AGEMA_signal_13992 ;
    wire new_AGEMA_signal_13993 ;
    wire new_AGEMA_signal_13994 ;
    wire new_AGEMA_signal_13995 ;
    wire new_AGEMA_signal_13996 ;
    wire new_AGEMA_signal_13997 ;
    wire new_AGEMA_signal_13998 ;
    wire new_AGEMA_signal_13999 ;
    wire new_AGEMA_signal_14000 ;
    wire new_AGEMA_signal_14001 ;
    wire new_AGEMA_signal_14002 ;
    wire new_AGEMA_signal_14003 ;
    wire new_AGEMA_signal_14004 ;
    wire new_AGEMA_signal_14005 ;
    wire new_AGEMA_signal_14006 ;
    wire new_AGEMA_signal_14007 ;
    wire new_AGEMA_signal_14008 ;
    wire new_AGEMA_signal_14009 ;
    wire new_AGEMA_signal_14010 ;
    wire new_AGEMA_signal_14011 ;
    wire new_AGEMA_signal_14012 ;
    wire new_AGEMA_signal_14013 ;
    wire new_AGEMA_signal_14014 ;
    wire new_AGEMA_signal_14015 ;
    wire new_AGEMA_signal_14016 ;
    wire new_AGEMA_signal_14017 ;
    wire new_AGEMA_signal_14018 ;
    wire new_AGEMA_signal_14019 ;
    wire new_AGEMA_signal_14020 ;
    wire new_AGEMA_signal_14021 ;
    wire new_AGEMA_signal_14022 ;
    wire new_AGEMA_signal_14023 ;
    wire new_AGEMA_signal_14024 ;
    wire new_AGEMA_signal_14025 ;
    wire new_AGEMA_signal_14026 ;
    wire new_AGEMA_signal_14027 ;
    wire new_AGEMA_signal_14028 ;
    wire new_AGEMA_signal_14029 ;
    wire new_AGEMA_signal_14030 ;
    wire new_AGEMA_signal_14031 ;
    wire new_AGEMA_signal_14032 ;
    wire new_AGEMA_signal_14033 ;
    wire new_AGEMA_signal_14034 ;
    wire new_AGEMA_signal_14035 ;
    wire new_AGEMA_signal_14036 ;
    wire new_AGEMA_signal_14037 ;
    wire new_AGEMA_signal_14038 ;
    wire new_AGEMA_signal_14039 ;
    wire new_AGEMA_signal_14040 ;
    wire new_AGEMA_signal_14041 ;
    wire new_AGEMA_signal_14042 ;
    wire new_AGEMA_signal_14043 ;
    wire new_AGEMA_signal_14044 ;
    wire new_AGEMA_signal_14045 ;
    wire new_AGEMA_signal_14046 ;
    wire new_AGEMA_signal_14047 ;
    wire new_AGEMA_signal_14048 ;
    wire new_AGEMA_signal_14049 ;
    wire new_AGEMA_signal_14050 ;
    wire new_AGEMA_signal_14051 ;
    wire new_AGEMA_signal_14052 ;
    wire new_AGEMA_signal_14053 ;
    wire new_AGEMA_signal_14054 ;
    wire new_AGEMA_signal_14055 ;
    wire new_AGEMA_signal_14056 ;
    wire new_AGEMA_signal_14057 ;
    wire new_AGEMA_signal_14058 ;
    wire new_AGEMA_signal_14059 ;
    wire new_AGEMA_signal_14060 ;
    wire new_AGEMA_signal_14061 ;
    wire new_AGEMA_signal_14062 ;
    wire new_AGEMA_signal_14063 ;
    wire new_AGEMA_signal_14064 ;
    wire new_AGEMA_signal_14065 ;
    wire new_AGEMA_signal_14066 ;
    wire new_AGEMA_signal_14067 ;
    wire new_AGEMA_signal_14068 ;
    wire new_AGEMA_signal_14069 ;
    wire new_AGEMA_signal_14070 ;
    wire new_AGEMA_signal_14071 ;
    wire new_AGEMA_signal_14072 ;
    wire new_AGEMA_signal_14073 ;
    wire new_AGEMA_signal_14074 ;
    wire new_AGEMA_signal_14075 ;
    wire new_AGEMA_signal_14076 ;
    wire new_AGEMA_signal_14077 ;
    wire new_AGEMA_signal_14078 ;
    wire new_AGEMA_signal_14079 ;
    wire new_AGEMA_signal_14080 ;
    wire new_AGEMA_signal_14081 ;
    wire new_AGEMA_signal_14082 ;
    wire new_AGEMA_signal_14083 ;
    wire new_AGEMA_signal_14084 ;
    wire new_AGEMA_signal_14085 ;
    wire new_AGEMA_signal_14086 ;
    wire new_AGEMA_signal_14087 ;
    wire new_AGEMA_signal_14088 ;
    wire new_AGEMA_signal_14089 ;
    wire new_AGEMA_signal_14090 ;
    wire new_AGEMA_signal_14091 ;
    wire new_AGEMA_signal_14092 ;
    wire new_AGEMA_signal_14093 ;
    wire new_AGEMA_signal_14094 ;
    wire new_AGEMA_signal_14095 ;
    wire new_AGEMA_signal_14096 ;
    wire new_AGEMA_signal_14097 ;
    wire new_AGEMA_signal_14098 ;
    wire new_AGEMA_signal_14099 ;
    wire new_AGEMA_signal_14100 ;
    wire new_AGEMA_signal_14101 ;
    wire new_AGEMA_signal_14102 ;
    wire new_AGEMA_signal_14103 ;
    wire new_AGEMA_signal_14104 ;
    wire new_AGEMA_signal_14105 ;
    wire new_AGEMA_signal_14106 ;
    wire new_AGEMA_signal_14107 ;
    wire new_AGEMA_signal_14108 ;
    wire new_AGEMA_signal_14109 ;
    wire new_AGEMA_signal_14110 ;
    wire new_AGEMA_signal_14111 ;
    wire new_AGEMA_signal_14112 ;
    wire new_AGEMA_signal_14113 ;
    wire new_AGEMA_signal_14114 ;
    wire new_AGEMA_signal_14115 ;
    wire new_AGEMA_signal_14116 ;
    wire new_AGEMA_signal_14117 ;
    wire new_AGEMA_signal_14118 ;
    wire new_AGEMA_signal_14119 ;
    wire new_AGEMA_signal_14120 ;
    wire new_AGEMA_signal_14121 ;
    wire new_AGEMA_signal_14122 ;
    wire new_AGEMA_signal_14123 ;
    wire new_AGEMA_signal_14124 ;
    wire new_AGEMA_signal_14125 ;
    wire new_AGEMA_signal_14126 ;
    wire new_AGEMA_signal_14127 ;
    wire new_AGEMA_signal_14128 ;
    wire new_AGEMA_signal_14129 ;
    wire new_AGEMA_signal_14130 ;
    wire new_AGEMA_signal_14131 ;
    wire new_AGEMA_signal_14132 ;
    wire new_AGEMA_signal_14133 ;
    wire new_AGEMA_signal_14134 ;
    wire new_AGEMA_signal_14135 ;
    wire new_AGEMA_signal_14136 ;
    wire new_AGEMA_signal_14137 ;
    wire new_AGEMA_signal_14138 ;
    wire new_AGEMA_signal_14139 ;
    wire new_AGEMA_signal_14140 ;
    wire new_AGEMA_signal_14141 ;
    wire new_AGEMA_signal_14142 ;
    wire new_AGEMA_signal_14143 ;
    wire new_AGEMA_signal_14144 ;
    wire new_AGEMA_signal_14145 ;
    wire new_AGEMA_signal_14146 ;
    wire new_AGEMA_signal_14147 ;
    wire new_AGEMA_signal_14148 ;
    wire new_AGEMA_signal_14149 ;
    wire new_AGEMA_signal_14150 ;
    wire new_AGEMA_signal_14151 ;
    wire new_AGEMA_signal_14152 ;
    wire new_AGEMA_signal_14153 ;
    wire new_AGEMA_signal_14154 ;
    wire new_AGEMA_signal_14155 ;
    wire new_AGEMA_signal_14156 ;
    wire new_AGEMA_signal_14157 ;
    wire new_AGEMA_signal_14158 ;
    wire new_AGEMA_signal_14159 ;
    wire new_AGEMA_signal_14160 ;
    wire new_AGEMA_signal_14161 ;
    wire new_AGEMA_signal_14162 ;
    wire new_AGEMA_signal_14163 ;
    wire new_AGEMA_signal_14164 ;
    wire new_AGEMA_signal_14165 ;
    wire new_AGEMA_signal_14166 ;
    wire new_AGEMA_signal_14167 ;
    wire new_AGEMA_signal_14168 ;
    wire new_AGEMA_signal_14169 ;
    wire new_AGEMA_signal_14170 ;
    wire new_AGEMA_signal_14171 ;
    wire new_AGEMA_signal_14172 ;
    wire new_AGEMA_signal_14173 ;
    wire new_AGEMA_signal_14174 ;
    wire new_AGEMA_signal_14175 ;
    wire new_AGEMA_signal_14176 ;
    wire new_AGEMA_signal_14177 ;
    wire new_AGEMA_signal_14178 ;
    wire new_AGEMA_signal_14179 ;
    wire new_AGEMA_signal_14180 ;
    wire new_AGEMA_signal_14181 ;
    wire new_AGEMA_signal_14182 ;
    wire new_AGEMA_signal_14183 ;
    wire new_AGEMA_signal_14184 ;
    wire new_AGEMA_signal_14185 ;
    wire new_AGEMA_signal_14186 ;
    wire new_AGEMA_signal_14187 ;
    wire new_AGEMA_signal_14188 ;
    wire new_AGEMA_signal_14189 ;
    wire new_AGEMA_signal_14190 ;
    wire new_AGEMA_signal_14191 ;
    wire new_AGEMA_signal_14192 ;
    wire new_AGEMA_signal_14193 ;
    wire new_AGEMA_signal_14194 ;
    wire new_AGEMA_signal_14195 ;
    wire new_AGEMA_signal_14196 ;
    wire new_AGEMA_signal_14197 ;
    wire new_AGEMA_signal_14198 ;
    wire new_AGEMA_signal_14199 ;
    wire new_AGEMA_signal_14200 ;
    wire new_AGEMA_signal_14201 ;
    wire new_AGEMA_signal_14202 ;
    wire new_AGEMA_signal_14203 ;
    wire new_AGEMA_signal_14204 ;
    wire new_AGEMA_signal_14205 ;
    wire new_AGEMA_signal_14206 ;
    wire new_AGEMA_signal_14207 ;
    wire new_AGEMA_signal_14208 ;
    wire new_AGEMA_signal_14209 ;
    wire new_AGEMA_signal_14210 ;
    wire new_AGEMA_signal_14211 ;
    wire new_AGEMA_signal_14212 ;
    wire new_AGEMA_signal_14213 ;
    wire new_AGEMA_signal_14214 ;
    wire new_AGEMA_signal_14215 ;
    wire new_AGEMA_signal_14216 ;
    wire new_AGEMA_signal_14217 ;
    wire new_AGEMA_signal_14218 ;
    wire new_AGEMA_signal_14219 ;
    wire new_AGEMA_signal_14220 ;
    wire new_AGEMA_signal_14221 ;
    wire new_AGEMA_signal_14222 ;
    wire new_AGEMA_signal_14223 ;
    wire new_AGEMA_signal_14224 ;
    wire new_AGEMA_signal_14225 ;
    wire new_AGEMA_signal_14226 ;
    wire new_AGEMA_signal_14227 ;
    wire new_AGEMA_signal_14228 ;
    wire new_AGEMA_signal_14229 ;
    wire new_AGEMA_signal_14230 ;
    wire new_AGEMA_signal_14231 ;
    wire new_AGEMA_signal_14232 ;
    wire new_AGEMA_signal_14233 ;
    wire new_AGEMA_signal_14234 ;
    wire new_AGEMA_signal_14235 ;
    wire new_AGEMA_signal_14236 ;
    wire new_AGEMA_signal_14237 ;
    wire new_AGEMA_signal_14238 ;
    wire new_AGEMA_signal_14239 ;
    wire new_AGEMA_signal_14240 ;
    wire new_AGEMA_signal_14241 ;
    wire new_AGEMA_signal_14242 ;
    wire new_AGEMA_signal_14243 ;
    wire new_AGEMA_signal_14244 ;
    wire new_AGEMA_signal_14245 ;
    wire new_AGEMA_signal_14246 ;
    wire new_AGEMA_signal_14247 ;
    wire new_AGEMA_signal_14248 ;
    wire new_AGEMA_signal_14249 ;
    wire new_AGEMA_signal_14250 ;
    wire new_AGEMA_signal_14251 ;
    wire new_AGEMA_signal_14252 ;
    wire new_AGEMA_signal_14253 ;
    wire new_AGEMA_signal_14254 ;
    wire new_AGEMA_signal_14255 ;
    wire new_AGEMA_signal_14256 ;
    wire new_AGEMA_signal_14257 ;
    wire new_AGEMA_signal_14258 ;
    wire new_AGEMA_signal_14259 ;
    wire new_AGEMA_signal_14260 ;
    wire new_AGEMA_signal_14261 ;
    wire new_AGEMA_signal_14262 ;
    wire new_AGEMA_signal_14263 ;
    wire new_AGEMA_signal_14264 ;
    wire new_AGEMA_signal_14265 ;
    wire new_AGEMA_signal_14266 ;
    wire new_AGEMA_signal_14267 ;
    wire new_AGEMA_signal_14268 ;
    wire new_AGEMA_signal_14269 ;
    wire new_AGEMA_signal_14270 ;
    wire new_AGEMA_signal_14271 ;
    wire new_AGEMA_signal_14272 ;
    wire new_AGEMA_signal_14273 ;
    wire new_AGEMA_signal_14274 ;
    wire new_AGEMA_signal_14275 ;
    wire new_AGEMA_signal_14276 ;
    wire new_AGEMA_signal_14277 ;
    wire new_AGEMA_signal_14278 ;
    wire new_AGEMA_signal_14279 ;
    wire new_AGEMA_signal_14280 ;
    wire new_AGEMA_signal_14281 ;
    wire new_AGEMA_signal_14282 ;
    wire new_AGEMA_signal_14283 ;
    wire new_AGEMA_signal_14284 ;
    wire new_AGEMA_signal_14285 ;
    wire new_AGEMA_signal_14286 ;
    wire new_AGEMA_signal_14287 ;
    wire new_AGEMA_signal_14288 ;
    wire new_AGEMA_signal_14289 ;
    wire new_AGEMA_signal_14290 ;
    wire new_AGEMA_signal_14291 ;
    wire new_AGEMA_signal_14292 ;
    wire new_AGEMA_signal_14293 ;
    wire new_AGEMA_signal_14294 ;
    wire new_AGEMA_signal_14295 ;
    wire new_AGEMA_signal_14296 ;
    wire new_AGEMA_signal_14297 ;
    wire new_AGEMA_signal_14298 ;
    wire new_AGEMA_signal_14299 ;
    wire new_AGEMA_signal_14300 ;
    wire new_AGEMA_signal_14301 ;
    wire new_AGEMA_signal_14302 ;
    wire new_AGEMA_signal_14303 ;
    wire new_AGEMA_signal_14304 ;
    wire new_AGEMA_signal_14305 ;
    wire new_AGEMA_signal_14306 ;
    wire new_AGEMA_signal_14307 ;
    wire new_AGEMA_signal_14308 ;
    wire new_AGEMA_signal_14309 ;
    wire new_AGEMA_signal_14310 ;
    wire new_AGEMA_signal_14311 ;
    wire new_AGEMA_signal_14312 ;
    wire new_AGEMA_signal_14313 ;
    wire new_AGEMA_signal_14314 ;
    wire new_AGEMA_signal_14315 ;
    wire new_AGEMA_signal_14316 ;
    wire new_AGEMA_signal_14317 ;
    wire new_AGEMA_signal_14318 ;
    wire new_AGEMA_signal_14319 ;
    wire new_AGEMA_signal_14320 ;
    wire new_AGEMA_signal_14321 ;
    wire new_AGEMA_signal_14322 ;
    wire new_AGEMA_signal_14323 ;
    wire new_AGEMA_signal_14324 ;
    wire new_AGEMA_signal_14325 ;
    wire new_AGEMA_signal_14326 ;
    wire new_AGEMA_signal_14327 ;
    wire new_AGEMA_signal_14328 ;
    wire new_AGEMA_signal_14329 ;
    wire new_AGEMA_signal_14330 ;
    wire new_AGEMA_signal_14331 ;
    wire new_AGEMA_signal_14332 ;
    wire new_AGEMA_signal_14333 ;
    wire new_AGEMA_signal_14334 ;
    wire new_AGEMA_signal_14335 ;
    wire new_AGEMA_signal_14336 ;
    wire new_AGEMA_signal_14337 ;
    wire new_AGEMA_signal_14338 ;
    wire new_AGEMA_signal_14339 ;
    wire new_AGEMA_signal_14340 ;
    wire new_AGEMA_signal_14341 ;
    wire new_AGEMA_signal_14342 ;
    wire new_AGEMA_signal_14343 ;
    wire new_AGEMA_signal_14344 ;
    wire new_AGEMA_signal_14345 ;
    wire new_AGEMA_signal_14346 ;
    wire new_AGEMA_signal_14347 ;
    wire new_AGEMA_signal_14348 ;
    wire new_AGEMA_signal_14349 ;
    wire new_AGEMA_signal_14350 ;
    wire new_AGEMA_signal_14351 ;
    wire new_AGEMA_signal_14352 ;
    wire new_AGEMA_signal_14353 ;
    wire new_AGEMA_signal_14354 ;
    wire new_AGEMA_signal_14355 ;
    wire new_AGEMA_signal_14356 ;
    wire new_AGEMA_signal_14357 ;
    wire new_AGEMA_signal_14358 ;
    wire new_AGEMA_signal_14359 ;
    wire new_AGEMA_signal_14360 ;
    wire new_AGEMA_signal_14361 ;
    wire new_AGEMA_signal_14362 ;
    wire new_AGEMA_signal_14363 ;
    wire new_AGEMA_signal_14364 ;
    wire new_AGEMA_signal_14365 ;
    wire new_AGEMA_signal_14366 ;
    wire new_AGEMA_signal_14367 ;
    wire new_AGEMA_signal_14368 ;
    wire new_AGEMA_signal_14369 ;
    wire new_AGEMA_signal_14370 ;
    wire new_AGEMA_signal_14371 ;
    wire new_AGEMA_signal_14372 ;
    wire new_AGEMA_signal_14373 ;
    wire new_AGEMA_signal_14374 ;
    wire new_AGEMA_signal_14375 ;
    wire new_AGEMA_signal_14376 ;
    wire new_AGEMA_signal_14377 ;
    wire new_AGEMA_signal_14378 ;
    wire new_AGEMA_signal_14379 ;
    wire new_AGEMA_signal_14380 ;
    wire new_AGEMA_signal_14381 ;
    wire new_AGEMA_signal_14382 ;
    wire new_AGEMA_signal_14383 ;
    wire new_AGEMA_signal_14384 ;
    wire new_AGEMA_signal_14385 ;
    wire new_AGEMA_signal_14386 ;
    wire new_AGEMA_signal_14387 ;
    wire new_AGEMA_signal_14388 ;
    wire new_AGEMA_signal_14389 ;
    wire new_AGEMA_signal_14390 ;
    wire new_AGEMA_signal_14391 ;
    wire new_AGEMA_signal_14392 ;
    wire new_AGEMA_signal_14393 ;
    wire new_AGEMA_signal_14394 ;
    wire new_AGEMA_signal_14395 ;
    wire new_AGEMA_signal_14396 ;
    wire new_AGEMA_signal_14397 ;
    wire new_AGEMA_signal_14398 ;
    wire new_AGEMA_signal_14399 ;
    wire new_AGEMA_signal_14400 ;
    wire new_AGEMA_signal_14401 ;
    wire new_AGEMA_signal_14402 ;
    wire new_AGEMA_signal_14403 ;
    wire new_AGEMA_signal_14404 ;
    wire new_AGEMA_signal_14405 ;
    wire new_AGEMA_signal_14406 ;
    wire new_AGEMA_signal_14407 ;
    wire new_AGEMA_signal_14408 ;
    wire new_AGEMA_signal_14409 ;
    wire new_AGEMA_signal_14410 ;
    wire new_AGEMA_signal_14411 ;
    wire new_AGEMA_signal_14412 ;
    wire new_AGEMA_signal_14413 ;
    wire new_AGEMA_signal_14414 ;
    wire new_AGEMA_signal_14415 ;
    wire new_AGEMA_signal_14416 ;
    wire new_AGEMA_signal_14417 ;
    wire new_AGEMA_signal_14418 ;
    wire new_AGEMA_signal_14419 ;
    wire new_AGEMA_signal_14420 ;
    wire new_AGEMA_signal_14421 ;
    wire new_AGEMA_signal_14422 ;
    wire new_AGEMA_signal_14423 ;
    wire new_AGEMA_signal_14424 ;
    wire new_AGEMA_signal_14425 ;
    wire new_AGEMA_signal_14426 ;
    wire new_AGEMA_signal_14427 ;
    wire new_AGEMA_signal_14428 ;
    wire new_AGEMA_signal_14429 ;
    wire new_AGEMA_signal_14430 ;
    wire new_AGEMA_signal_14431 ;
    wire new_AGEMA_signal_14432 ;
    wire new_AGEMA_signal_14433 ;
    wire new_AGEMA_signal_14434 ;
    wire new_AGEMA_signal_14435 ;
    wire new_AGEMA_signal_14436 ;
    wire new_AGEMA_signal_14437 ;
    wire new_AGEMA_signal_14438 ;
    wire new_AGEMA_signal_14439 ;
    wire new_AGEMA_signal_14440 ;
    wire new_AGEMA_signal_14441 ;
    wire new_AGEMA_signal_14442 ;
    wire new_AGEMA_signal_14443 ;
    wire new_AGEMA_signal_14444 ;
    wire new_AGEMA_signal_14445 ;
    wire new_AGEMA_signal_14446 ;
    wire new_AGEMA_signal_14447 ;
    wire new_AGEMA_signal_14448 ;
    wire new_AGEMA_signal_14449 ;
    wire new_AGEMA_signal_14450 ;
    wire new_AGEMA_signal_14451 ;
    wire new_AGEMA_signal_14452 ;
    wire new_AGEMA_signal_14453 ;
    wire new_AGEMA_signal_14454 ;
    wire new_AGEMA_signal_14455 ;
    wire new_AGEMA_signal_14456 ;
    wire new_AGEMA_signal_14457 ;
    wire new_AGEMA_signal_14458 ;
    wire new_AGEMA_signal_14459 ;
    wire new_AGEMA_signal_14460 ;
    wire new_AGEMA_signal_14461 ;
    wire new_AGEMA_signal_14462 ;
    wire new_AGEMA_signal_14463 ;
    wire new_AGEMA_signal_14464 ;
    wire new_AGEMA_signal_14465 ;
    wire new_AGEMA_signal_14466 ;
    wire new_AGEMA_signal_14467 ;
    wire new_AGEMA_signal_14468 ;
    wire new_AGEMA_signal_14469 ;
    wire new_AGEMA_signal_14470 ;
    wire new_AGEMA_signal_14471 ;
    wire new_AGEMA_signal_14472 ;
    wire new_AGEMA_signal_14473 ;
    wire new_AGEMA_signal_14474 ;
    wire new_AGEMA_signal_14475 ;
    wire new_AGEMA_signal_14476 ;
    wire new_AGEMA_signal_14477 ;
    wire new_AGEMA_signal_14478 ;
    wire new_AGEMA_signal_14479 ;
    wire new_AGEMA_signal_14480 ;
    wire new_AGEMA_signal_14481 ;
    wire new_AGEMA_signal_14482 ;
    wire new_AGEMA_signal_14483 ;
    wire new_AGEMA_signal_14484 ;
    wire new_AGEMA_signal_14485 ;
    wire new_AGEMA_signal_14486 ;
    wire new_AGEMA_signal_14487 ;
    wire new_AGEMA_signal_14488 ;
    wire new_AGEMA_signal_14489 ;
    wire new_AGEMA_signal_14490 ;
    wire new_AGEMA_signal_14491 ;
    wire new_AGEMA_signal_14492 ;
    wire new_AGEMA_signal_14493 ;
    wire new_AGEMA_signal_14494 ;
    wire new_AGEMA_signal_14495 ;
    wire new_AGEMA_signal_14496 ;
    wire new_AGEMA_signal_14497 ;
    wire new_AGEMA_signal_14498 ;
    wire new_AGEMA_signal_14499 ;
    wire new_AGEMA_signal_14500 ;
    wire new_AGEMA_signal_14501 ;
    wire new_AGEMA_signal_14502 ;
    wire new_AGEMA_signal_14503 ;
    wire new_AGEMA_signal_14504 ;
    wire new_AGEMA_signal_14505 ;
    wire new_AGEMA_signal_14506 ;
    wire new_AGEMA_signal_14507 ;
    wire new_AGEMA_signal_14508 ;
    wire new_AGEMA_signal_14509 ;
    wire new_AGEMA_signal_14510 ;
    wire new_AGEMA_signal_14511 ;
    wire new_AGEMA_signal_14512 ;
    wire new_AGEMA_signal_14513 ;
    wire new_AGEMA_signal_14514 ;
    wire new_AGEMA_signal_14515 ;
    wire new_AGEMA_signal_14516 ;
    wire new_AGEMA_signal_14517 ;
    wire new_AGEMA_signal_14518 ;
    wire new_AGEMA_signal_14519 ;
    wire new_AGEMA_signal_14520 ;
    wire new_AGEMA_signal_14521 ;
    wire new_AGEMA_signal_14522 ;
    wire new_AGEMA_signal_14523 ;
    wire new_AGEMA_signal_14524 ;
    wire new_AGEMA_signal_14525 ;
    wire new_AGEMA_signal_14526 ;
    wire new_AGEMA_signal_14527 ;
    wire new_AGEMA_signal_14528 ;
    wire new_AGEMA_signal_14529 ;
    wire new_AGEMA_signal_14530 ;
    wire new_AGEMA_signal_14531 ;
    wire new_AGEMA_signal_14532 ;
    wire new_AGEMA_signal_14533 ;
    wire new_AGEMA_signal_14534 ;
    wire new_AGEMA_signal_14535 ;
    wire new_AGEMA_signal_14536 ;
    wire new_AGEMA_signal_14537 ;
    wire new_AGEMA_signal_14538 ;
    wire new_AGEMA_signal_14539 ;
    wire new_AGEMA_signal_14540 ;
    wire new_AGEMA_signal_14541 ;
    wire new_AGEMA_signal_14542 ;
    wire new_AGEMA_signal_14543 ;
    wire new_AGEMA_signal_14544 ;
    wire new_AGEMA_signal_14545 ;
    wire new_AGEMA_signal_14546 ;
    wire new_AGEMA_signal_14547 ;
    wire new_AGEMA_signal_14548 ;
    wire new_AGEMA_signal_14549 ;
    wire new_AGEMA_signal_14550 ;
    wire new_AGEMA_signal_14551 ;
    wire new_AGEMA_signal_14552 ;
    wire new_AGEMA_signal_14553 ;
    wire new_AGEMA_signal_14554 ;
    wire new_AGEMA_signal_14555 ;
    wire new_AGEMA_signal_14556 ;
    wire new_AGEMA_signal_14557 ;
    wire new_AGEMA_signal_14558 ;
    wire new_AGEMA_signal_14559 ;
    wire new_AGEMA_signal_14560 ;
    wire new_AGEMA_signal_14561 ;
    wire new_AGEMA_signal_14562 ;
    wire new_AGEMA_signal_14563 ;
    wire new_AGEMA_signal_14564 ;
    wire new_AGEMA_signal_14565 ;
    wire new_AGEMA_signal_14566 ;
    wire new_AGEMA_signal_14567 ;
    wire new_AGEMA_signal_14568 ;
    wire new_AGEMA_signal_14569 ;
    wire new_AGEMA_signal_14570 ;
    wire new_AGEMA_signal_14571 ;
    wire new_AGEMA_signal_14572 ;
    wire new_AGEMA_signal_14573 ;
    wire new_AGEMA_signal_14574 ;
    wire new_AGEMA_signal_14575 ;
    wire new_AGEMA_signal_14576 ;
    wire new_AGEMA_signal_14577 ;
    wire new_AGEMA_signal_14578 ;
    wire new_AGEMA_signal_14579 ;
    wire new_AGEMA_signal_14580 ;
    wire new_AGEMA_signal_14581 ;
    wire new_AGEMA_signal_14582 ;
    wire new_AGEMA_signal_14583 ;
    wire new_AGEMA_signal_14584 ;
    wire new_AGEMA_signal_14585 ;
    wire new_AGEMA_signal_14586 ;
    wire new_AGEMA_signal_14587 ;
    wire new_AGEMA_signal_14588 ;
    wire new_AGEMA_signal_14589 ;
    wire new_AGEMA_signal_14590 ;
    wire new_AGEMA_signal_14591 ;
    wire new_AGEMA_signal_14592 ;
    wire new_AGEMA_signal_14593 ;
    wire new_AGEMA_signal_14594 ;
    wire new_AGEMA_signal_14595 ;
    wire new_AGEMA_signal_14596 ;
    wire new_AGEMA_signal_14597 ;
    wire new_AGEMA_signal_14598 ;
    wire new_AGEMA_signal_14599 ;
    wire new_AGEMA_signal_14600 ;
    wire new_AGEMA_signal_14601 ;
    wire new_AGEMA_signal_14602 ;
    wire new_AGEMA_signal_14603 ;
    wire new_AGEMA_signal_14604 ;
    wire new_AGEMA_signal_14605 ;
    wire new_AGEMA_signal_14606 ;
    wire new_AGEMA_signal_14607 ;
    wire new_AGEMA_signal_14608 ;
    wire new_AGEMA_signal_14609 ;
    wire new_AGEMA_signal_14610 ;
    wire new_AGEMA_signal_14611 ;
    wire new_AGEMA_signal_14612 ;
    wire new_AGEMA_signal_14613 ;
    wire new_AGEMA_signal_14614 ;
    wire new_AGEMA_signal_14615 ;
    wire new_AGEMA_signal_14616 ;
    wire new_AGEMA_signal_14617 ;
    wire new_AGEMA_signal_14618 ;
    wire new_AGEMA_signal_14619 ;
    wire new_AGEMA_signal_14620 ;
    wire new_AGEMA_signal_14621 ;
    wire new_AGEMA_signal_14622 ;
    wire new_AGEMA_signal_14623 ;
    wire new_AGEMA_signal_14624 ;
    wire new_AGEMA_signal_14625 ;
    wire new_AGEMA_signal_14626 ;
    wire new_AGEMA_signal_14627 ;
    wire new_AGEMA_signal_14628 ;
    wire new_AGEMA_signal_14629 ;
    wire new_AGEMA_signal_14630 ;
    wire new_AGEMA_signal_14631 ;
    wire new_AGEMA_signal_14632 ;
    wire new_AGEMA_signal_14633 ;
    wire new_AGEMA_signal_14634 ;
    wire new_AGEMA_signal_14635 ;
    wire new_AGEMA_signal_14636 ;
    wire new_AGEMA_signal_14637 ;
    wire new_AGEMA_signal_14638 ;
    wire new_AGEMA_signal_14639 ;
    wire new_AGEMA_signal_14640 ;
    wire new_AGEMA_signal_14641 ;
    wire new_AGEMA_signal_14642 ;
    wire new_AGEMA_signal_14643 ;
    wire new_AGEMA_signal_14644 ;
    wire new_AGEMA_signal_14645 ;
    wire new_AGEMA_signal_14646 ;
    wire new_AGEMA_signal_14647 ;
    wire new_AGEMA_signal_14648 ;
    wire new_AGEMA_signal_14649 ;
    wire new_AGEMA_signal_14650 ;
    wire new_AGEMA_signal_14651 ;
    wire new_AGEMA_signal_14652 ;
    wire new_AGEMA_signal_14653 ;
    wire new_AGEMA_signal_14654 ;
    wire new_AGEMA_signal_14655 ;
    wire new_AGEMA_signal_14656 ;
    wire new_AGEMA_signal_14657 ;
    wire new_AGEMA_signal_14658 ;
    wire new_AGEMA_signal_14659 ;
    wire new_AGEMA_signal_14660 ;
    wire new_AGEMA_signal_14661 ;
    wire new_AGEMA_signal_14662 ;
    wire new_AGEMA_signal_14663 ;
    wire new_AGEMA_signal_14664 ;
    wire new_AGEMA_signal_14665 ;
    wire new_AGEMA_signal_14666 ;
    wire new_AGEMA_signal_14667 ;
    wire new_AGEMA_signal_14668 ;
    wire new_AGEMA_signal_14669 ;
    wire new_AGEMA_signal_14670 ;
    wire new_AGEMA_signal_14671 ;
    wire new_AGEMA_signal_14672 ;
    wire new_AGEMA_signal_14673 ;
    wire new_AGEMA_signal_14674 ;
    wire new_AGEMA_signal_14675 ;
    wire new_AGEMA_signal_14676 ;
    wire new_AGEMA_signal_14677 ;
    wire new_AGEMA_signal_14678 ;
    wire new_AGEMA_signal_14679 ;
    wire new_AGEMA_signal_14680 ;
    wire new_AGEMA_signal_14681 ;
    wire new_AGEMA_signal_14682 ;
    wire new_AGEMA_signal_14683 ;
    wire new_AGEMA_signal_14684 ;
    wire new_AGEMA_signal_14685 ;
    wire new_AGEMA_signal_14686 ;
    wire new_AGEMA_signal_14687 ;
    wire new_AGEMA_signal_14688 ;
    wire new_AGEMA_signal_14689 ;
    wire new_AGEMA_signal_14690 ;
    wire new_AGEMA_signal_14691 ;
    wire new_AGEMA_signal_14692 ;
    wire new_AGEMA_signal_14693 ;
    wire new_AGEMA_signal_14694 ;
    wire new_AGEMA_signal_14695 ;
    wire new_AGEMA_signal_14696 ;
    wire new_AGEMA_signal_14697 ;
    wire new_AGEMA_signal_14698 ;
    wire new_AGEMA_signal_14699 ;
    wire new_AGEMA_signal_14700 ;
    wire new_AGEMA_signal_14701 ;
    wire new_AGEMA_signal_14702 ;
    wire new_AGEMA_signal_14703 ;
    wire new_AGEMA_signal_14704 ;
    wire new_AGEMA_signal_14705 ;
    wire new_AGEMA_signal_14706 ;
    wire new_AGEMA_signal_14707 ;
    wire new_AGEMA_signal_14708 ;
    wire new_AGEMA_signal_14709 ;
    wire new_AGEMA_signal_14710 ;
    wire new_AGEMA_signal_14711 ;
    wire new_AGEMA_signal_14712 ;
    wire new_AGEMA_signal_14713 ;
    wire new_AGEMA_signal_14714 ;
    wire new_AGEMA_signal_14715 ;
    wire new_AGEMA_signal_14716 ;
    wire new_AGEMA_signal_14717 ;
    wire new_AGEMA_signal_14718 ;
    wire new_AGEMA_signal_14719 ;
    wire new_AGEMA_signal_14720 ;
    wire new_AGEMA_signal_14721 ;
    wire new_AGEMA_signal_14722 ;
    wire new_AGEMA_signal_14723 ;
    wire new_AGEMA_signal_14724 ;
    wire new_AGEMA_signal_14725 ;
    wire new_AGEMA_signal_14726 ;
    wire new_AGEMA_signal_14727 ;
    wire new_AGEMA_signal_14728 ;
    wire new_AGEMA_signal_14729 ;
    wire new_AGEMA_signal_14730 ;
    wire new_AGEMA_signal_14731 ;
    wire new_AGEMA_signal_14732 ;
    wire new_AGEMA_signal_14733 ;
    wire new_AGEMA_signal_14734 ;
    wire new_AGEMA_signal_14735 ;
    wire new_AGEMA_signal_14736 ;
    wire new_AGEMA_signal_14737 ;
    wire new_AGEMA_signal_14738 ;
    wire new_AGEMA_signal_14739 ;
    wire new_AGEMA_signal_14740 ;
    wire new_AGEMA_signal_14741 ;
    wire new_AGEMA_signal_14742 ;
    wire new_AGEMA_signal_14743 ;
    wire new_AGEMA_signal_14744 ;
    wire new_AGEMA_signal_14745 ;
    wire new_AGEMA_signal_14746 ;
    wire new_AGEMA_signal_14747 ;
    wire new_AGEMA_signal_14748 ;
    wire new_AGEMA_signal_14749 ;
    wire new_AGEMA_signal_14750 ;
    wire new_AGEMA_signal_14751 ;
    wire new_AGEMA_signal_14752 ;
    wire new_AGEMA_signal_14753 ;
    wire new_AGEMA_signal_14754 ;
    wire new_AGEMA_signal_14755 ;
    wire new_AGEMA_signal_14756 ;
    wire new_AGEMA_signal_14757 ;
    wire new_AGEMA_signal_14758 ;
    wire new_AGEMA_signal_14759 ;
    wire new_AGEMA_signal_14760 ;
    wire new_AGEMA_signal_14761 ;
    wire new_AGEMA_signal_14762 ;
    wire new_AGEMA_signal_14763 ;
    wire new_AGEMA_signal_14764 ;
    wire new_AGEMA_signal_14765 ;
    wire new_AGEMA_signal_14766 ;
    wire new_AGEMA_signal_14767 ;
    wire new_AGEMA_signal_14768 ;
    wire new_AGEMA_signal_14769 ;
    wire new_AGEMA_signal_14770 ;
    wire new_AGEMA_signal_14771 ;
    wire new_AGEMA_signal_14772 ;
    wire new_AGEMA_signal_14773 ;
    wire new_AGEMA_signal_14774 ;
    wire new_AGEMA_signal_14775 ;
    wire new_AGEMA_signal_14776 ;
    wire new_AGEMA_signal_14777 ;
    wire new_AGEMA_signal_14778 ;
    wire new_AGEMA_signal_14779 ;
    wire new_AGEMA_signal_14780 ;
    wire new_AGEMA_signal_14781 ;
    wire new_AGEMA_signal_14782 ;
    wire new_AGEMA_signal_14783 ;
    wire new_AGEMA_signal_14784 ;
    wire new_AGEMA_signal_14785 ;
    wire new_AGEMA_signal_14786 ;
    wire new_AGEMA_signal_14787 ;
    wire new_AGEMA_signal_14788 ;
    wire new_AGEMA_signal_14789 ;
    wire new_AGEMA_signal_14790 ;
    wire new_AGEMA_signal_14791 ;
    wire new_AGEMA_signal_14792 ;
    wire new_AGEMA_signal_14793 ;
    wire new_AGEMA_signal_14794 ;
    wire new_AGEMA_signal_14795 ;
    wire new_AGEMA_signal_14796 ;
    wire new_AGEMA_signal_14797 ;
    wire new_AGEMA_signal_14798 ;
    wire new_AGEMA_signal_14799 ;
    wire new_AGEMA_signal_14800 ;
    wire new_AGEMA_signal_14801 ;
    wire new_AGEMA_signal_14802 ;
    wire new_AGEMA_signal_14803 ;
    wire new_AGEMA_signal_14804 ;
    wire new_AGEMA_signal_14805 ;
    wire new_AGEMA_signal_14806 ;
    wire new_AGEMA_signal_14807 ;
    wire new_AGEMA_signal_14808 ;
    wire new_AGEMA_signal_14809 ;
    wire new_AGEMA_signal_14813 ;
    wire new_AGEMA_signal_14814 ;
    wire new_AGEMA_signal_14815 ;
    wire new_AGEMA_signal_14819 ;
    wire new_AGEMA_signal_14820 ;
    wire new_AGEMA_signal_14821 ;
    wire new_AGEMA_signal_14825 ;
    wire new_AGEMA_signal_14826 ;
    wire new_AGEMA_signal_14827 ;
    wire new_AGEMA_signal_14828 ;
    wire new_AGEMA_signal_14829 ;
    wire new_AGEMA_signal_14830 ;
    wire new_AGEMA_signal_14834 ;
    wire new_AGEMA_signal_14835 ;
    wire new_AGEMA_signal_14836 ;
    wire new_AGEMA_signal_14840 ;
    wire new_AGEMA_signal_14841 ;
    wire new_AGEMA_signal_14842 ;
    wire new_AGEMA_signal_14846 ;
    wire new_AGEMA_signal_14847 ;
    wire new_AGEMA_signal_14848 ;
    wire new_AGEMA_signal_14852 ;
    wire new_AGEMA_signal_14853 ;
    wire new_AGEMA_signal_14854 ;
    wire new_AGEMA_signal_14858 ;
    wire new_AGEMA_signal_14859 ;
    wire new_AGEMA_signal_14860 ;
    wire new_AGEMA_signal_14864 ;
    wire new_AGEMA_signal_14865 ;
    wire new_AGEMA_signal_14866 ;
    wire new_AGEMA_signal_14870 ;
    wire new_AGEMA_signal_14871 ;
    wire new_AGEMA_signal_14872 ;
    wire new_AGEMA_signal_14873 ;
    wire new_AGEMA_signal_14874 ;
    wire new_AGEMA_signal_14875 ;
    wire new_AGEMA_signal_14879 ;
    wire new_AGEMA_signal_14880 ;
    wire new_AGEMA_signal_14881 ;
    wire new_AGEMA_signal_14885 ;
    wire new_AGEMA_signal_14886 ;
    wire new_AGEMA_signal_14887 ;
    wire new_AGEMA_signal_14891 ;
    wire new_AGEMA_signal_14892 ;
    wire new_AGEMA_signal_14893 ;
    wire new_AGEMA_signal_14897 ;
    wire new_AGEMA_signal_14898 ;
    wire new_AGEMA_signal_14899 ;
    wire new_AGEMA_signal_14903 ;
    wire new_AGEMA_signal_14904 ;
    wire new_AGEMA_signal_14905 ;
    wire new_AGEMA_signal_14909 ;
    wire new_AGEMA_signal_14910 ;
    wire new_AGEMA_signal_14911 ;
    wire new_AGEMA_signal_14915 ;
    wire new_AGEMA_signal_14916 ;
    wire new_AGEMA_signal_14917 ;
    wire new_AGEMA_signal_14918 ;
    wire new_AGEMA_signal_14919 ;
    wire new_AGEMA_signal_14920 ;
    wire new_AGEMA_signal_14924 ;
    wire new_AGEMA_signal_14925 ;
    wire new_AGEMA_signal_14926 ;
    wire new_AGEMA_signal_14930 ;
    wire new_AGEMA_signal_14931 ;
    wire new_AGEMA_signal_14932 ;
    wire new_AGEMA_signal_14936 ;
    wire new_AGEMA_signal_14937 ;
    wire new_AGEMA_signal_14938 ;
    wire new_AGEMA_signal_14942 ;
    wire new_AGEMA_signal_14943 ;
    wire new_AGEMA_signal_14944 ;
    wire new_AGEMA_signal_14948 ;
    wire new_AGEMA_signal_14949 ;
    wire new_AGEMA_signal_14950 ;
    wire new_AGEMA_signal_14954 ;
    wire new_AGEMA_signal_14955 ;
    wire new_AGEMA_signal_14956 ;
    wire new_AGEMA_signal_14960 ;
    wire new_AGEMA_signal_14961 ;
    wire new_AGEMA_signal_14962 ;
    wire new_AGEMA_signal_14966 ;
    wire new_AGEMA_signal_14967 ;
    wire new_AGEMA_signal_14968 ;
    wire new_AGEMA_signal_14969 ;
    wire new_AGEMA_signal_14970 ;
    wire new_AGEMA_signal_14971 ;
    wire new_AGEMA_signal_14972 ;
    wire new_AGEMA_signal_14973 ;
    wire new_AGEMA_signal_14974 ;
    wire new_AGEMA_signal_14975 ;
    wire new_AGEMA_signal_14976 ;
    wire new_AGEMA_signal_14977 ;
    wire new_AGEMA_signal_14978 ;
    wire new_AGEMA_signal_14979 ;
    wire new_AGEMA_signal_14980 ;
    wire new_AGEMA_signal_14981 ;
    wire new_AGEMA_signal_14982 ;
    wire new_AGEMA_signal_14983 ;
    wire new_AGEMA_signal_14984 ;
    wire new_AGEMA_signal_14985 ;
    wire new_AGEMA_signal_14986 ;
    wire new_AGEMA_signal_14987 ;
    wire new_AGEMA_signal_14988 ;
    wire new_AGEMA_signal_14989 ;
    wire new_AGEMA_signal_14990 ;
    wire new_AGEMA_signal_14991 ;
    wire new_AGEMA_signal_14992 ;
    wire new_AGEMA_signal_14993 ;
    wire new_AGEMA_signal_14994 ;
    wire new_AGEMA_signal_14995 ;
    wire new_AGEMA_signal_14996 ;
    wire new_AGEMA_signal_14997 ;
    wire new_AGEMA_signal_14998 ;
    wire new_AGEMA_signal_14999 ;
    wire new_AGEMA_signal_15000 ;
    wire new_AGEMA_signal_15001 ;
    wire new_AGEMA_signal_15002 ;
    wire new_AGEMA_signal_15003 ;
    wire new_AGEMA_signal_15004 ;
    wire new_AGEMA_signal_15005 ;
    wire new_AGEMA_signal_15006 ;
    wire new_AGEMA_signal_15007 ;
    wire new_AGEMA_signal_15008 ;
    wire new_AGEMA_signal_15009 ;
    wire new_AGEMA_signal_15010 ;
    wire new_AGEMA_signal_15011 ;
    wire new_AGEMA_signal_15012 ;
    wire new_AGEMA_signal_15013 ;
    wire new_AGEMA_signal_15014 ;
    wire new_AGEMA_signal_15015 ;
    wire new_AGEMA_signal_15016 ;
    wire new_AGEMA_signal_15017 ;
    wire new_AGEMA_signal_15018 ;
    wire new_AGEMA_signal_15019 ;
    wire new_AGEMA_signal_15020 ;
    wire new_AGEMA_signal_15021 ;
    wire new_AGEMA_signal_15022 ;
    wire new_AGEMA_signal_15023 ;
    wire new_AGEMA_signal_15024 ;
    wire new_AGEMA_signal_15025 ;
    wire new_AGEMA_signal_15026 ;
    wire new_AGEMA_signal_15027 ;
    wire new_AGEMA_signal_15028 ;
    wire new_AGEMA_signal_15029 ;
    wire new_AGEMA_signal_15030 ;
    wire new_AGEMA_signal_15031 ;
    wire new_AGEMA_signal_15032 ;
    wire new_AGEMA_signal_15033 ;
    wire new_AGEMA_signal_15034 ;
    wire new_AGEMA_signal_15035 ;
    wire new_AGEMA_signal_15036 ;
    wire new_AGEMA_signal_15037 ;
    wire new_AGEMA_signal_15038 ;
    wire new_AGEMA_signal_15039 ;
    wire new_AGEMA_signal_15040 ;
    wire new_AGEMA_signal_15041 ;
    wire new_AGEMA_signal_15042 ;
    wire new_AGEMA_signal_15043 ;
    wire new_AGEMA_signal_15044 ;
    wire new_AGEMA_signal_15045 ;
    wire new_AGEMA_signal_15046 ;
    wire new_AGEMA_signal_15047 ;
    wire new_AGEMA_signal_15048 ;
    wire new_AGEMA_signal_15049 ;
    wire new_AGEMA_signal_15050 ;
    wire new_AGEMA_signal_15051 ;
    wire new_AGEMA_signal_15052 ;
    wire new_AGEMA_signal_15053 ;
    wire new_AGEMA_signal_15054 ;
    wire new_AGEMA_signal_15055 ;
    wire new_AGEMA_signal_15056 ;
    wire new_AGEMA_signal_15057 ;
    wire new_AGEMA_signal_15058 ;
    wire new_AGEMA_signal_15059 ;
    wire new_AGEMA_signal_15060 ;
    wire new_AGEMA_signal_15061 ;
    wire new_AGEMA_signal_15062 ;
    wire new_AGEMA_signal_15063 ;
    wire new_AGEMA_signal_15064 ;
    wire new_AGEMA_signal_15065 ;
    wire new_AGEMA_signal_15066 ;
    wire new_AGEMA_signal_15067 ;
    wire new_AGEMA_signal_15068 ;
    wire new_AGEMA_signal_15069 ;
    wire new_AGEMA_signal_15070 ;
    wire new_AGEMA_signal_15071 ;
    wire new_AGEMA_signal_15072 ;
    wire new_AGEMA_signal_15073 ;
    wire new_AGEMA_signal_15074 ;
    wire new_AGEMA_signal_15075 ;
    wire new_AGEMA_signal_15076 ;
    wire new_AGEMA_signal_15077 ;
    wire new_AGEMA_signal_15078 ;
    wire new_AGEMA_signal_15079 ;
    wire new_AGEMA_signal_15080 ;
    wire new_AGEMA_signal_15081 ;
    wire new_AGEMA_signal_15082 ;
    wire new_AGEMA_signal_15083 ;
    wire new_AGEMA_signal_15084 ;
    wire new_AGEMA_signal_15085 ;
    wire new_AGEMA_signal_15086 ;
    wire new_AGEMA_signal_15087 ;
    wire new_AGEMA_signal_15088 ;
    wire new_AGEMA_signal_15089 ;
    wire new_AGEMA_signal_15090 ;
    wire new_AGEMA_signal_15091 ;
    wire new_AGEMA_signal_15092 ;
    wire new_AGEMA_signal_15093 ;
    wire new_AGEMA_signal_15094 ;
    wire new_AGEMA_signal_15095 ;
    wire new_AGEMA_signal_15096 ;
    wire new_AGEMA_signal_15097 ;
    wire new_AGEMA_signal_15098 ;
    wire new_AGEMA_signal_15099 ;
    wire new_AGEMA_signal_15100 ;
    wire new_AGEMA_signal_15101 ;
    wire new_AGEMA_signal_15102 ;
    wire new_AGEMA_signal_15103 ;
    wire new_AGEMA_signal_15104 ;
    wire new_AGEMA_signal_15105 ;
    wire new_AGEMA_signal_15106 ;
    wire new_AGEMA_signal_15107 ;
    wire new_AGEMA_signal_15108 ;
    wire new_AGEMA_signal_15109 ;
    wire new_AGEMA_signal_15110 ;
    wire new_AGEMA_signal_15111 ;
    wire new_AGEMA_signal_15112 ;
    wire new_AGEMA_signal_15113 ;
    wire new_AGEMA_signal_15114 ;
    wire new_AGEMA_signal_15115 ;
    wire new_AGEMA_signal_15116 ;
    wire new_AGEMA_signal_15117 ;
    wire new_AGEMA_signal_15118 ;
    wire new_AGEMA_signal_15119 ;
    wire new_AGEMA_signal_15120 ;
    wire new_AGEMA_signal_15121 ;
    wire new_AGEMA_signal_15122 ;
    wire new_AGEMA_signal_15123 ;
    wire new_AGEMA_signal_15124 ;
    wire new_AGEMA_signal_15125 ;
    wire new_AGEMA_signal_15126 ;
    wire new_AGEMA_signal_15127 ;
    wire new_AGEMA_signal_15128 ;
    wire new_AGEMA_signal_15129 ;
    wire new_AGEMA_signal_15130 ;
    wire new_AGEMA_signal_15131 ;
    wire new_AGEMA_signal_15132 ;
    wire new_AGEMA_signal_15133 ;
    wire new_AGEMA_signal_15134 ;
    wire new_AGEMA_signal_15135 ;
    wire new_AGEMA_signal_15136 ;
    wire new_AGEMA_signal_15137 ;
    wire new_AGEMA_signal_15138 ;
    wire new_AGEMA_signal_15139 ;
    wire new_AGEMA_signal_15140 ;
    wire new_AGEMA_signal_15141 ;
    wire new_AGEMA_signal_15142 ;
    wire new_AGEMA_signal_15143 ;
    wire new_AGEMA_signal_15144 ;
    wire new_AGEMA_signal_15145 ;
    wire new_AGEMA_signal_15146 ;
    wire new_AGEMA_signal_15147 ;
    wire new_AGEMA_signal_15148 ;
    wire new_AGEMA_signal_15149 ;
    wire new_AGEMA_signal_15150 ;
    wire new_AGEMA_signal_15151 ;
    wire new_AGEMA_signal_15152 ;
    wire new_AGEMA_signal_15153 ;
    wire new_AGEMA_signal_15154 ;
    wire new_AGEMA_signal_15155 ;
    wire new_AGEMA_signal_15156 ;
    wire new_AGEMA_signal_15157 ;
    wire new_AGEMA_signal_15158 ;
    wire new_AGEMA_signal_15159 ;
    wire new_AGEMA_signal_15160 ;
    wire new_AGEMA_signal_15161 ;
    wire new_AGEMA_signal_15162 ;
    wire new_AGEMA_signal_15163 ;
    wire new_AGEMA_signal_15164 ;
    wire new_AGEMA_signal_15165 ;
    wire new_AGEMA_signal_15166 ;
    wire new_AGEMA_signal_15167 ;
    wire new_AGEMA_signal_15168 ;
    wire new_AGEMA_signal_15169 ;
    wire new_AGEMA_signal_15170 ;
    wire new_AGEMA_signal_15171 ;
    wire new_AGEMA_signal_15172 ;
    wire new_AGEMA_signal_15173 ;
    wire new_AGEMA_signal_15174 ;
    wire new_AGEMA_signal_15175 ;
    wire new_AGEMA_signal_15176 ;
    wire new_AGEMA_signal_15177 ;
    wire new_AGEMA_signal_15178 ;
    wire new_AGEMA_signal_15179 ;
    wire new_AGEMA_signal_15180 ;
    wire new_AGEMA_signal_15181 ;
    wire new_AGEMA_signal_15182 ;
    wire new_AGEMA_signal_15183 ;
    wire new_AGEMA_signal_15184 ;
    wire new_AGEMA_signal_15185 ;
    wire new_AGEMA_signal_15186 ;
    wire new_AGEMA_signal_15187 ;
    wire new_AGEMA_signal_15188 ;
    wire new_AGEMA_signal_15189 ;
    wire new_AGEMA_signal_15190 ;
    wire new_AGEMA_signal_15191 ;
    wire new_AGEMA_signal_15192 ;
    wire new_AGEMA_signal_15193 ;
    wire new_AGEMA_signal_15194 ;
    wire new_AGEMA_signal_15195 ;
    wire new_AGEMA_signal_15196 ;
    wire new_AGEMA_signal_15197 ;
    wire new_AGEMA_signal_15198 ;
    wire new_AGEMA_signal_15199 ;
    wire new_AGEMA_signal_15200 ;
    wire new_AGEMA_signal_15201 ;
    wire new_AGEMA_signal_15202 ;
    wire new_AGEMA_signal_15203 ;
    wire new_AGEMA_signal_15204 ;
    wire new_AGEMA_signal_15205 ;
    wire new_AGEMA_signal_15206 ;
    wire new_AGEMA_signal_15207 ;
    wire new_AGEMA_signal_15208 ;
    wire new_AGEMA_signal_15209 ;
    wire new_AGEMA_signal_15210 ;
    wire new_AGEMA_signal_15211 ;
    wire new_AGEMA_signal_15212 ;
    wire new_AGEMA_signal_15213 ;
    wire new_AGEMA_signal_15214 ;
    wire new_AGEMA_signal_15215 ;
    wire new_AGEMA_signal_15216 ;
    wire new_AGEMA_signal_15217 ;
    wire new_AGEMA_signal_15218 ;
    wire new_AGEMA_signal_15219 ;
    wire new_AGEMA_signal_15220 ;
    wire new_AGEMA_signal_15221 ;
    wire new_AGEMA_signal_15222 ;
    wire new_AGEMA_signal_15223 ;
    wire new_AGEMA_signal_15224 ;
    wire new_AGEMA_signal_15225 ;
    wire new_AGEMA_signal_15226 ;
    wire new_AGEMA_signal_15227 ;
    wire new_AGEMA_signal_15228 ;
    wire new_AGEMA_signal_15229 ;
    wire new_AGEMA_signal_15230 ;
    wire new_AGEMA_signal_15231 ;
    wire new_AGEMA_signal_15232 ;
    wire new_AGEMA_signal_15233 ;
    wire new_AGEMA_signal_15234 ;
    wire new_AGEMA_signal_15235 ;
    wire new_AGEMA_signal_15236 ;
    wire new_AGEMA_signal_15237 ;
    wire new_AGEMA_signal_15238 ;
    wire new_AGEMA_signal_15239 ;
    wire new_AGEMA_signal_15240 ;
    wire new_AGEMA_signal_15241 ;
    wire new_AGEMA_signal_15242 ;
    wire new_AGEMA_signal_15243 ;
    wire new_AGEMA_signal_15244 ;
    wire new_AGEMA_signal_15245 ;
    wire new_AGEMA_signal_15246 ;
    wire new_AGEMA_signal_15247 ;
    wire new_AGEMA_signal_15248 ;
    wire new_AGEMA_signal_15249 ;
    wire new_AGEMA_signal_15250 ;
    wire new_AGEMA_signal_15251 ;
    wire new_AGEMA_signal_15252 ;
    wire new_AGEMA_signal_15253 ;
    wire new_AGEMA_signal_15254 ;
    wire new_AGEMA_signal_15255 ;
    wire new_AGEMA_signal_15256 ;
    wire new_AGEMA_signal_15257 ;
    wire new_AGEMA_signal_15258 ;
    wire new_AGEMA_signal_15259 ;
    wire new_AGEMA_signal_15260 ;
    wire new_AGEMA_signal_15261 ;
    wire new_AGEMA_signal_15262 ;
    wire new_AGEMA_signal_15263 ;
    wire new_AGEMA_signal_15264 ;
    wire new_AGEMA_signal_15265 ;
    wire new_AGEMA_signal_15266 ;
    wire new_AGEMA_signal_15267 ;
    wire new_AGEMA_signal_15268 ;
    wire new_AGEMA_signal_15269 ;
    wire new_AGEMA_signal_15270 ;
    wire new_AGEMA_signal_15271 ;
    wire new_AGEMA_signal_15272 ;
    wire new_AGEMA_signal_15273 ;
    wire new_AGEMA_signal_15274 ;
    wire new_AGEMA_signal_15275 ;
    wire new_AGEMA_signal_15276 ;
    wire new_AGEMA_signal_15277 ;
    wire new_AGEMA_signal_15278 ;
    wire new_AGEMA_signal_15279 ;
    wire new_AGEMA_signal_15280 ;
    wire new_AGEMA_signal_15281 ;
    wire new_AGEMA_signal_15282 ;
    wire new_AGEMA_signal_15283 ;
    wire new_AGEMA_signal_15284 ;
    wire new_AGEMA_signal_15285 ;
    wire new_AGEMA_signal_15286 ;
    wire new_AGEMA_signal_15287 ;
    wire new_AGEMA_signal_15288 ;
    wire new_AGEMA_signal_15289 ;
    wire new_AGEMA_signal_15290 ;
    wire new_AGEMA_signal_15291 ;
    wire new_AGEMA_signal_15292 ;
    wire new_AGEMA_signal_15293 ;
    wire new_AGEMA_signal_15294 ;
    wire new_AGEMA_signal_15295 ;
    wire new_AGEMA_signal_15296 ;
    wire new_AGEMA_signal_15297 ;
    wire new_AGEMA_signal_15298 ;
    wire new_AGEMA_signal_15299 ;
    wire new_AGEMA_signal_15300 ;
    wire new_AGEMA_signal_15301 ;
    wire new_AGEMA_signal_15302 ;
    wire new_AGEMA_signal_15303 ;
    wire new_AGEMA_signal_15304 ;
    wire new_AGEMA_signal_15305 ;
    wire new_AGEMA_signal_15306 ;
    wire new_AGEMA_signal_15307 ;
    wire new_AGEMA_signal_15308 ;
    wire new_AGEMA_signal_15309 ;
    wire new_AGEMA_signal_15310 ;
    wire new_AGEMA_signal_15311 ;
    wire new_AGEMA_signal_15312 ;
    wire new_AGEMA_signal_15313 ;
    wire new_AGEMA_signal_15314 ;
    wire new_AGEMA_signal_15315 ;
    wire new_AGEMA_signal_15316 ;
    wire new_AGEMA_signal_15317 ;
    wire new_AGEMA_signal_15318 ;
    wire new_AGEMA_signal_15319 ;
    wire new_AGEMA_signal_15320 ;
    wire new_AGEMA_signal_15321 ;
    wire new_AGEMA_signal_15322 ;
    wire new_AGEMA_signal_15323 ;
    wire new_AGEMA_signal_15324 ;
    wire new_AGEMA_signal_15325 ;
    wire new_AGEMA_signal_15326 ;
    wire new_AGEMA_signal_15327 ;
    wire new_AGEMA_signal_15328 ;
    wire new_AGEMA_signal_15329 ;
    wire new_AGEMA_signal_15330 ;
    wire new_AGEMA_signal_15331 ;
    wire new_AGEMA_signal_15332 ;
    wire new_AGEMA_signal_15333 ;
    wire new_AGEMA_signal_15334 ;
    wire new_AGEMA_signal_15335 ;
    wire new_AGEMA_signal_15336 ;
    wire new_AGEMA_signal_15337 ;
    wire new_AGEMA_signal_15338 ;
    wire new_AGEMA_signal_15339 ;
    wire new_AGEMA_signal_15340 ;
    wire new_AGEMA_signal_15341 ;
    wire new_AGEMA_signal_15342 ;
    wire new_AGEMA_signal_15343 ;
    wire new_AGEMA_signal_15344 ;
    wire new_AGEMA_signal_15345 ;
    wire new_AGEMA_signal_15346 ;
    wire new_AGEMA_signal_15347 ;
    wire new_AGEMA_signal_15348 ;
    wire new_AGEMA_signal_15349 ;
    wire new_AGEMA_signal_15350 ;
    wire new_AGEMA_signal_15351 ;
    wire new_AGEMA_signal_15352 ;
    wire new_AGEMA_signal_15353 ;
    wire new_AGEMA_signal_15354 ;
    wire new_AGEMA_signal_15355 ;
    wire new_AGEMA_signal_15356 ;
    wire new_AGEMA_signal_15357 ;
    wire new_AGEMA_signal_15358 ;
    wire new_AGEMA_signal_15359 ;
    wire new_AGEMA_signal_15360 ;
    wire new_AGEMA_signal_15361 ;
    wire new_AGEMA_signal_15362 ;
    wire new_AGEMA_signal_15363 ;
    wire new_AGEMA_signal_15364 ;
    wire new_AGEMA_signal_15365 ;
    wire new_AGEMA_signal_15366 ;
    wire new_AGEMA_signal_15367 ;
    wire new_AGEMA_signal_15368 ;
    wire new_AGEMA_signal_15369 ;
    wire new_AGEMA_signal_15370 ;
    wire new_AGEMA_signal_15371 ;
    wire new_AGEMA_signal_15372 ;
    wire new_AGEMA_signal_15373 ;
    wire new_AGEMA_signal_15374 ;
    wire new_AGEMA_signal_15375 ;
    wire new_AGEMA_signal_15376 ;
    wire new_AGEMA_signal_15377 ;
    wire new_AGEMA_signal_15378 ;
    wire new_AGEMA_signal_15379 ;
    wire new_AGEMA_signal_15380 ;
    wire new_AGEMA_signal_15381 ;
    wire new_AGEMA_signal_15382 ;
    wire new_AGEMA_signal_15383 ;
    wire new_AGEMA_signal_15384 ;
    wire new_AGEMA_signal_15385 ;
    wire new_AGEMA_signal_15386 ;
    wire new_AGEMA_signal_15387 ;
    wire new_AGEMA_signal_15388 ;
    wire new_AGEMA_signal_15389 ;
    wire new_AGEMA_signal_15390 ;
    wire new_AGEMA_signal_15391 ;
    wire new_AGEMA_signal_15392 ;
    wire new_AGEMA_signal_15393 ;
    wire new_AGEMA_signal_15394 ;
    wire new_AGEMA_signal_15395 ;
    wire new_AGEMA_signal_15396 ;
    wire new_AGEMA_signal_15397 ;
    wire new_AGEMA_signal_15398 ;
    wire new_AGEMA_signal_15399 ;
    wire new_AGEMA_signal_15400 ;
    wire new_AGEMA_signal_15401 ;
    wire new_AGEMA_signal_15402 ;
    wire new_AGEMA_signal_15403 ;
    wire new_AGEMA_signal_15404 ;
    wire new_AGEMA_signal_15405 ;
    wire new_AGEMA_signal_15406 ;
    wire new_AGEMA_signal_15407 ;
    wire new_AGEMA_signal_15408 ;
    wire new_AGEMA_signal_15409 ;
    wire new_AGEMA_signal_15410 ;
    wire new_AGEMA_signal_15411 ;
    wire new_AGEMA_signal_15412 ;
    wire new_AGEMA_signal_15413 ;
    wire new_AGEMA_signal_15414 ;
    wire new_AGEMA_signal_15415 ;
    wire new_AGEMA_signal_15416 ;
    wire new_AGEMA_signal_15417 ;
    wire new_AGEMA_signal_15418 ;
    wire new_AGEMA_signal_15419 ;
    wire new_AGEMA_signal_15420 ;
    wire new_AGEMA_signal_15421 ;
    wire new_AGEMA_signal_15422 ;
    wire new_AGEMA_signal_15423 ;
    wire new_AGEMA_signal_15424 ;
    wire new_AGEMA_signal_15425 ;
    wire new_AGEMA_signal_15426 ;
    wire new_AGEMA_signal_15427 ;
    wire new_AGEMA_signal_15428 ;
    wire new_AGEMA_signal_15429 ;
    wire new_AGEMA_signal_15430 ;
    wire new_AGEMA_signal_15431 ;
    wire new_AGEMA_signal_15432 ;
    wire new_AGEMA_signal_15433 ;
    wire new_AGEMA_signal_15434 ;
    wire new_AGEMA_signal_15435 ;
    wire new_AGEMA_signal_15436 ;
    wire new_AGEMA_signal_15437 ;
    wire new_AGEMA_signal_15438 ;
    wire new_AGEMA_signal_15439 ;
    wire new_AGEMA_signal_15440 ;
    wire new_AGEMA_signal_15441 ;
    wire new_AGEMA_signal_15442 ;
    wire new_AGEMA_signal_15443 ;
    wire new_AGEMA_signal_15444 ;
    wire new_AGEMA_signal_15445 ;
    wire new_AGEMA_signal_15446 ;
    wire new_AGEMA_signal_15447 ;
    wire new_AGEMA_signal_15448 ;
    wire new_AGEMA_signal_15452 ;
    wire new_AGEMA_signal_15453 ;
    wire new_AGEMA_signal_15454 ;
    wire new_AGEMA_signal_15458 ;
    wire new_AGEMA_signal_15459 ;
    wire new_AGEMA_signal_15460 ;
    wire new_AGEMA_signal_15464 ;
    wire new_AGEMA_signal_15465 ;
    wire new_AGEMA_signal_15466 ;
    wire new_AGEMA_signal_15467 ;
    wire new_AGEMA_signal_15468 ;
    wire new_AGEMA_signal_15469 ;
    wire new_AGEMA_signal_15473 ;
    wire new_AGEMA_signal_15474 ;
    wire new_AGEMA_signal_15475 ;
    wire new_AGEMA_signal_15479 ;
    wire new_AGEMA_signal_15480 ;
    wire new_AGEMA_signal_15481 ;
    wire new_AGEMA_signal_15485 ;
    wire new_AGEMA_signal_15486 ;
    wire new_AGEMA_signal_15487 ;
    wire new_AGEMA_signal_15491 ;
    wire new_AGEMA_signal_15492 ;
    wire new_AGEMA_signal_15493 ;
    wire new_AGEMA_signal_15497 ;
    wire new_AGEMA_signal_15498 ;
    wire new_AGEMA_signal_15499 ;
    wire new_AGEMA_signal_15503 ;
    wire new_AGEMA_signal_15504 ;
    wire new_AGEMA_signal_15505 ;
    wire new_AGEMA_signal_15509 ;
    wire new_AGEMA_signal_15510 ;
    wire new_AGEMA_signal_15511 ;
    wire new_AGEMA_signal_15512 ;
    wire new_AGEMA_signal_15513 ;
    wire new_AGEMA_signal_15514 ;
    wire new_AGEMA_signal_15518 ;
    wire new_AGEMA_signal_15519 ;
    wire new_AGEMA_signal_15520 ;
    wire new_AGEMA_signal_15524 ;
    wire new_AGEMA_signal_15525 ;
    wire new_AGEMA_signal_15526 ;
    wire new_AGEMA_signal_15530 ;
    wire new_AGEMA_signal_15531 ;
    wire new_AGEMA_signal_15532 ;
    wire new_AGEMA_signal_15536 ;
    wire new_AGEMA_signal_15537 ;
    wire new_AGEMA_signal_15538 ;
    wire new_AGEMA_signal_15542 ;
    wire new_AGEMA_signal_15543 ;
    wire new_AGEMA_signal_15544 ;
    wire new_AGEMA_signal_15548 ;
    wire new_AGEMA_signal_15549 ;
    wire new_AGEMA_signal_15550 ;
    wire new_AGEMA_signal_15554 ;
    wire new_AGEMA_signal_15555 ;
    wire new_AGEMA_signal_15556 ;
    wire new_AGEMA_signal_15557 ;
    wire new_AGEMA_signal_15558 ;
    wire new_AGEMA_signal_15559 ;
    wire new_AGEMA_signal_15563 ;
    wire new_AGEMA_signal_15564 ;
    wire new_AGEMA_signal_15565 ;
    wire new_AGEMA_signal_15569 ;
    wire new_AGEMA_signal_15570 ;
    wire new_AGEMA_signal_15571 ;
    wire new_AGEMA_signal_15575 ;
    wire new_AGEMA_signal_15576 ;
    wire new_AGEMA_signal_15577 ;
    wire new_AGEMA_signal_15581 ;
    wire new_AGEMA_signal_15582 ;
    wire new_AGEMA_signal_15583 ;
    wire new_AGEMA_signal_15587 ;
    wire new_AGEMA_signal_15588 ;
    wire new_AGEMA_signal_15589 ;
    wire new_AGEMA_signal_15593 ;
    wire new_AGEMA_signal_15594 ;
    wire new_AGEMA_signal_15595 ;
    wire new_AGEMA_signal_15599 ;
    wire new_AGEMA_signal_15600 ;
    wire new_AGEMA_signal_15601 ;
    wire new_AGEMA_signal_15605 ;
    wire new_AGEMA_signal_15606 ;
    wire new_AGEMA_signal_15607 ;
    wire new_AGEMA_signal_15608 ;
    wire new_AGEMA_signal_15609 ;
    wire new_AGEMA_signal_15610 ;
    wire new_AGEMA_signal_15611 ;
    wire new_AGEMA_signal_15612 ;
    wire new_AGEMA_signal_15613 ;
    wire new_AGEMA_signal_15614 ;
    wire new_AGEMA_signal_15615 ;
    wire new_AGEMA_signal_15616 ;
    wire new_AGEMA_signal_15617 ;
    wire new_AGEMA_signal_15618 ;
    wire new_AGEMA_signal_15619 ;
    wire new_AGEMA_signal_15620 ;
    wire new_AGEMA_signal_15621 ;
    wire new_AGEMA_signal_15622 ;
    wire new_AGEMA_signal_15623 ;
    wire new_AGEMA_signal_15624 ;
    wire new_AGEMA_signal_15625 ;
    wire new_AGEMA_signal_15626 ;
    wire new_AGEMA_signal_15627 ;
    wire new_AGEMA_signal_15628 ;
    wire new_AGEMA_signal_15629 ;
    wire new_AGEMA_signal_15630 ;
    wire new_AGEMA_signal_15631 ;
    wire new_AGEMA_signal_15632 ;
    wire new_AGEMA_signal_15633 ;
    wire new_AGEMA_signal_15634 ;
    wire new_AGEMA_signal_15635 ;
    wire new_AGEMA_signal_15636 ;
    wire new_AGEMA_signal_15637 ;
    wire new_AGEMA_signal_15638 ;
    wire new_AGEMA_signal_15639 ;
    wire new_AGEMA_signal_15640 ;
    wire new_AGEMA_signal_15641 ;
    wire new_AGEMA_signal_15642 ;
    wire new_AGEMA_signal_15643 ;
    wire new_AGEMA_signal_15644 ;
    wire new_AGEMA_signal_15645 ;
    wire new_AGEMA_signal_15646 ;
    wire new_AGEMA_signal_15647 ;
    wire new_AGEMA_signal_15648 ;
    wire new_AGEMA_signal_15649 ;
    wire new_AGEMA_signal_15650 ;
    wire new_AGEMA_signal_15651 ;
    wire new_AGEMA_signal_15652 ;
    wire new_AGEMA_signal_15653 ;
    wire new_AGEMA_signal_15654 ;
    wire new_AGEMA_signal_15655 ;
    wire new_AGEMA_signal_15656 ;
    wire new_AGEMA_signal_15657 ;
    wire new_AGEMA_signal_15658 ;
    wire new_AGEMA_signal_15659 ;
    wire new_AGEMA_signal_15660 ;
    wire new_AGEMA_signal_15661 ;
    wire new_AGEMA_signal_15662 ;
    wire new_AGEMA_signal_15663 ;
    wire new_AGEMA_signal_15664 ;
    wire new_AGEMA_signal_15665 ;
    wire new_AGEMA_signal_15666 ;
    wire new_AGEMA_signal_15667 ;
    wire new_AGEMA_signal_15668 ;
    wire new_AGEMA_signal_15669 ;
    wire new_AGEMA_signal_15670 ;
    wire new_AGEMA_signal_15671 ;
    wire new_AGEMA_signal_15672 ;
    wire new_AGEMA_signal_15673 ;
    wire new_AGEMA_signal_15677 ;
    wire new_AGEMA_signal_15678 ;
    wire new_AGEMA_signal_15679 ;
    wire new_AGEMA_signal_15683 ;
    wire new_AGEMA_signal_15684 ;
    wire new_AGEMA_signal_15685 ;
    wire new_AGEMA_signal_15689 ;
    wire new_AGEMA_signal_15690 ;
    wire new_AGEMA_signal_15691 ;
    wire new_AGEMA_signal_15695 ;
    wire new_AGEMA_signal_15696 ;
    wire new_AGEMA_signal_15697 ;
    wire new_AGEMA_signal_15701 ;
    wire new_AGEMA_signal_15702 ;
    wire new_AGEMA_signal_15703 ;
    wire new_AGEMA_signal_15707 ;
    wire new_AGEMA_signal_15708 ;
    wire new_AGEMA_signal_15709 ;
    wire new_AGEMA_signal_15713 ;
    wire new_AGEMA_signal_15714 ;
    wire new_AGEMA_signal_15715 ;
    wire new_AGEMA_signal_15716 ;
    wire new_AGEMA_signal_15717 ;
    wire new_AGEMA_signal_15718 ;
    wire new_AGEMA_signal_15719 ;
    wire new_AGEMA_signal_15720 ;
    wire new_AGEMA_signal_15721 ;
    wire new_AGEMA_signal_15722 ;
    wire new_AGEMA_signal_15723 ;
    wire new_AGEMA_signal_15724 ;
    wire new_AGEMA_signal_15725 ;
    wire new_AGEMA_signal_15726 ;
    wire new_AGEMA_signal_15727 ;
    wire new_AGEMA_signal_15728 ;
    wire new_AGEMA_signal_15729 ;
    wire new_AGEMA_signal_15730 ;
    wire new_AGEMA_signal_15731 ;
    wire new_AGEMA_signal_15732 ;
    wire new_AGEMA_signal_15733 ;
    wire new_AGEMA_signal_15734 ;
    wire new_AGEMA_signal_15735 ;
    wire new_AGEMA_signal_15736 ;
    wire new_AGEMA_signal_15737 ;
    wire new_AGEMA_signal_15738 ;
    wire new_AGEMA_signal_15739 ;
    wire new_AGEMA_signal_15740 ;
    wire new_AGEMA_signal_15741 ;
    wire new_AGEMA_signal_15742 ;
    wire new_AGEMA_signal_15743 ;
    wire new_AGEMA_signal_15744 ;
    wire new_AGEMA_signal_15745 ;
    wire new_AGEMA_signal_15746 ;
    wire new_AGEMA_signal_15747 ;
    wire new_AGEMA_signal_15748 ;
    wire new_AGEMA_signal_15749 ;
    wire new_AGEMA_signal_15750 ;
    wire new_AGEMA_signal_15751 ;
    wire new_AGEMA_signal_15752 ;
    wire new_AGEMA_signal_15753 ;
    wire new_AGEMA_signal_15754 ;
    wire new_AGEMA_signal_15755 ;
    wire new_AGEMA_signal_15756 ;
    wire new_AGEMA_signal_15757 ;
    wire new_AGEMA_signal_15758 ;
    wire new_AGEMA_signal_15759 ;
    wire new_AGEMA_signal_15760 ;
    wire new_AGEMA_signal_15761 ;
    wire new_AGEMA_signal_15762 ;
    wire new_AGEMA_signal_15763 ;
    wire new_AGEMA_signal_15764 ;
    wire new_AGEMA_signal_15765 ;
    wire new_AGEMA_signal_15766 ;
    wire new_AGEMA_signal_15767 ;
    wire new_AGEMA_signal_15768 ;
    wire new_AGEMA_signal_15769 ;
    wire new_AGEMA_signal_15770 ;
    wire new_AGEMA_signal_15771 ;
    wire new_AGEMA_signal_15772 ;
    wire new_AGEMA_signal_15773 ;
    wire new_AGEMA_signal_15774 ;
    wire new_AGEMA_signal_15775 ;
    wire new_AGEMA_signal_15776 ;
    wire new_AGEMA_signal_15777 ;
    wire new_AGEMA_signal_15778 ;
    wire new_AGEMA_signal_15779 ;
    wire new_AGEMA_signal_15780 ;
    wire new_AGEMA_signal_15781 ;
    wire new_AGEMA_signal_15782 ;
    wire new_AGEMA_signal_15783 ;
    wire new_AGEMA_signal_15784 ;
    wire new_AGEMA_signal_15785 ;
    wire new_AGEMA_signal_15786 ;
    wire new_AGEMA_signal_15787 ;
    wire new_AGEMA_signal_15788 ;
    wire new_AGEMA_signal_15789 ;
    wire new_AGEMA_signal_15790 ;
    wire new_AGEMA_signal_15791 ;
    wire new_AGEMA_signal_15792 ;
    wire new_AGEMA_signal_15793 ;
    wire new_AGEMA_signal_15794 ;
    wire new_AGEMA_signal_15795 ;
    wire new_AGEMA_signal_15796 ;
    wire new_AGEMA_signal_15797 ;
    wire new_AGEMA_signal_15798 ;
    wire new_AGEMA_signal_15799 ;
    wire new_AGEMA_signal_15800 ;
    wire new_AGEMA_signal_15801 ;
    wire new_AGEMA_signal_15802 ;
    wire new_AGEMA_signal_15803 ;
    wire new_AGEMA_signal_15804 ;
    wire new_AGEMA_signal_15805 ;
    wire new_AGEMA_signal_15806 ;
    wire new_AGEMA_signal_15807 ;
    wire new_AGEMA_signal_15808 ;
    wire new_AGEMA_signal_15809 ;
    wire new_AGEMA_signal_15810 ;
    wire new_AGEMA_signal_15811 ;
    wire new_AGEMA_signal_15812 ;
    wire new_AGEMA_signal_15813 ;
    wire new_AGEMA_signal_15814 ;
    wire new_AGEMA_signal_15815 ;
    wire new_AGEMA_signal_15816 ;
    wire new_AGEMA_signal_15817 ;
    wire new_AGEMA_signal_15818 ;
    wire new_AGEMA_signal_15819 ;
    wire new_AGEMA_signal_15820 ;
    wire new_AGEMA_signal_15821 ;
    wire new_AGEMA_signal_15822 ;
    wire new_AGEMA_signal_15823 ;
    wire new_AGEMA_signal_15824 ;
    wire new_AGEMA_signal_15825 ;
    wire new_AGEMA_signal_15826 ;
    wire new_AGEMA_signal_15827 ;
    wire new_AGEMA_signal_15828 ;
    wire new_AGEMA_signal_15829 ;
    wire new_AGEMA_signal_15830 ;
    wire new_AGEMA_signal_15831 ;
    wire new_AGEMA_signal_15832 ;
    wire new_AGEMA_signal_15833 ;
    wire new_AGEMA_signal_15834 ;
    wire new_AGEMA_signal_15835 ;
    wire new_AGEMA_signal_15836 ;
    wire new_AGEMA_signal_15837 ;
    wire new_AGEMA_signal_15838 ;
    wire new_AGEMA_signal_15839 ;
    wire new_AGEMA_signal_15840 ;
    wire new_AGEMA_signal_15841 ;
    wire new_AGEMA_signal_15842 ;
    wire new_AGEMA_signal_15843 ;
    wire new_AGEMA_signal_15844 ;
    wire new_AGEMA_signal_15845 ;
    wire new_AGEMA_signal_15846 ;
    wire new_AGEMA_signal_15847 ;
    wire new_AGEMA_signal_15848 ;
    wire new_AGEMA_signal_15849 ;
    wire new_AGEMA_signal_15850 ;
    wire new_AGEMA_signal_15851 ;
    wire new_AGEMA_signal_15852 ;
    wire new_AGEMA_signal_15853 ;
    wire new_AGEMA_signal_15854 ;
    wire new_AGEMA_signal_15855 ;
    wire new_AGEMA_signal_15856 ;
    wire new_AGEMA_signal_15857 ;
    wire new_AGEMA_signal_15858 ;
    wire new_AGEMA_signal_15859 ;
    wire new_AGEMA_signal_15860 ;
    wire new_AGEMA_signal_15861 ;
    wire new_AGEMA_signal_15862 ;
    wire new_AGEMA_signal_15863 ;
    wire new_AGEMA_signal_15864 ;
    wire new_AGEMA_signal_15865 ;
    wire new_AGEMA_signal_15866 ;
    wire new_AGEMA_signal_15867 ;
    wire new_AGEMA_signal_15868 ;
    wire new_AGEMA_signal_15869 ;
    wire new_AGEMA_signal_15870 ;
    wire new_AGEMA_signal_15871 ;
    wire new_AGEMA_signal_15872 ;
    wire new_AGEMA_signal_15873 ;
    wire new_AGEMA_signal_15874 ;
    wire new_AGEMA_signal_15875 ;
    wire new_AGEMA_signal_15876 ;
    wire new_AGEMA_signal_15877 ;
    wire new_AGEMA_signal_15878 ;
    wire new_AGEMA_signal_15879 ;
    wire new_AGEMA_signal_15880 ;
    wire new_AGEMA_signal_15881 ;
    wire new_AGEMA_signal_15882 ;
    wire new_AGEMA_signal_15883 ;
    wire new_AGEMA_signal_15884 ;
    wire new_AGEMA_signal_15885 ;
    wire new_AGEMA_signal_15886 ;
    wire new_AGEMA_signal_15887 ;
    wire new_AGEMA_signal_15888 ;
    wire new_AGEMA_signal_15889 ;
    wire new_AGEMA_signal_15890 ;
    wire new_AGEMA_signal_15891 ;
    wire new_AGEMA_signal_15892 ;
    wire new_AGEMA_signal_15893 ;
    wire new_AGEMA_signal_15894 ;
    wire new_AGEMA_signal_15895 ;
    wire new_AGEMA_signal_15896 ;
    wire new_AGEMA_signal_15897 ;
    wire new_AGEMA_signal_15898 ;
    wire new_AGEMA_signal_15899 ;
    wire new_AGEMA_signal_15900 ;
    wire new_AGEMA_signal_15901 ;
    wire new_AGEMA_signal_15902 ;
    wire new_AGEMA_signal_15903 ;
    wire new_AGEMA_signal_15904 ;
    wire new_AGEMA_signal_15905 ;
    wire new_AGEMA_signal_15906 ;
    wire new_AGEMA_signal_15907 ;
    wire new_AGEMA_signal_15908 ;
    wire new_AGEMA_signal_15909 ;
    wire new_AGEMA_signal_15910 ;
    wire new_AGEMA_signal_15911 ;
    wire new_AGEMA_signal_15912 ;
    wire new_AGEMA_signal_15913 ;
    wire new_AGEMA_signal_15914 ;
    wire new_AGEMA_signal_15915 ;
    wire new_AGEMA_signal_15916 ;
    wire new_AGEMA_signal_15917 ;
    wire new_AGEMA_signal_15918 ;
    wire new_AGEMA_signal_15919 ;
    wire new_AGEMA_signal_15920 ;
    wire new_AGEMA_signal_15921 ;
    wire new_AGEMA_signal_15922 ;
    wire new_AGEMA_signal_15923 ;
    wire new_AGEMA_signal_15924 ;
    wire new_AGEMA_signal_15925 ;
    wire new_AGEMA_signal_15926 ;
    wire new_AGEMA_signal_15927 ;
    wire new_AGEMA_signal_15928 ;
    wire new_AGEMA_signal_15929 ;
    wire new_AGEMA_signal_15930 ;
    wire new_AGEMA_signal_15931 ;
    wire new_AGEMA_signal_15932 ;
    wire new_AGEMA_signal_15933 ;
    wire new_AGEMA_signal_15934 ;
    wire new_AGEMA_signal_15935 ;
    wire new_AGEMA_signal_15936 ;
    wire new_AGEMA_signal_15937 ;
    wire new_AGEMA_signal_15938 ;
    wire new_AGEMA_signal_15939 ;
    wire new_AGEMA_signal_15940 ;
    wire new_AGEMA_signal_15941 ;
    wire new_AGEMA_signal_15942 ;
    wire new_AGEMA_signal_15943 ;
    wire new_AGEMA_signal_15944 ;
    wire new_AGEMA_signal_15945 ;
    wire new_AGEMA_signal_15946 ;
    wire new_AGEMA_signal_15947 ;
    wire new_AGEMA_signal_15948 ;
    wire new_AGEMA_signal_15949 ;
    wire new_AGEMA_signal_15950 ;
    wire new_AGEMA_signal_15951 ;
    wire new_AGEMA_signal_15952 ;
    wire new_AGEMA_signal_15953 ;
    wire new_AGEMA_signal_15954 ;
    wire new_AGEMA_signal_15955 ;
    wire new_AGEMA_signal_15956 ;
    wire new_AGEMA_signal_15957 ;
    wire new_AGEMA_signal_15958 ;
    wire new_AGEMA_signal_15959 ;
    wire new_AGEMA_signal_15960 ;
    wire new_AGEMA_signal_15961 ;
    wire new_AGEMA_signal_15962 ;
    wire new_AGEMA_signal_15963 ;
    wire new_AGEMA_signal_15964 ;
    wire new_AGEMA_signal_15965 ;
    wire new_AGEMA_signal_15966 ;
    wire new_AGEMA_signal_15967 ;
    wire new_AGEMA_signal_15968 ;
    wire new_AGEMA_signal_15969 ;
    wire new_AGEMA_signal_15970 ;
    wire new_AGEMA_signal_15971 ;
    wire new_AGEMA_signal_15972 ;
    wire new_AGEMA_signal_15973 ;
    wire new_AGEMA_signal_15974 ;
    wire new_AGEMA_signal_15975 ;
    wire new_AGEMA_signal_15976 ;
    wire new_AGEMA_signal_15977 ;
    wire new_AGEMA_signal_15978 ;
    wire new_AGEMA_signal_15979 ;
    wire new_AGEMA_signal_15980 ;
    wire new_AGEMA_signal_15981 ;
    wire new_AGEMA_signal_15982 ;
    wire new_AGEMA_signal_15983 ;
    wire new_AGEMA_signal_15984 ;
    wire new_AGEMA_signal_15985 ;
    wire new_AGEMA_signal_15986 ;
    wire new_AGEMA_signal_15987 ;
    wire new_AGEMA_signal_15988 ;
    wire new_AGEMA_signal_15989 ;
    wire new_AGEMA_signal_15990 ;
    wire new_AGEMA_signal_15991 ;
    wire new_AGEMA_signal_15992 ;
    wire new_AGEMA_signal_15993 ;
    wire new_AGEMA_signal_15994 ;
    wire new_AGEMA_signal_15995 ;
    wire new_AGEMA_signal_15996 ;
    wire new_AGEMA_signal_15997 ;
    wire new_AGEMA_signal_15998 ;
    wire new_AGEMA_signal_15999 ;
    wire new_AGEMA_signal_16000 ;
    wire new_AGEMA_signal_16001 ;
    wire new_AGEMA_signal_16002 ;
    wire new_AGEMA_signal_16003 ;
    wire new_AGEMA_signal_16004 ;
    wire new_AGEMA_signal_16005 ;
    wire new_AGEMA_signal_16006 ;
    wire new_AGEMA_signal_16007 ;
    wire new_AGEMA_signal_16008 ;
    wire new_AGEMA_signal_16009 ;
    wire new_AGEMA_signal_16010 ;
    wire new_AGEMA_signal_16011 ;
    wire new_AGEMA_signal_16012 ;
    wire new_AGEMA_signal_16013 ;
    wire new_AGEMA_signal_16014 ;
    wire new_AGEMA_signal_16015 ;
    wire new_AGEMA_signal_16016 ;
    wire new_AGEMA_signal_16017 ;
    wire new_AGEMA_signal_16018 ;
    wire new_AGEMA_signal_16019 ;
    wire new_AGEMA_signal_16020 ;
    wire new_AGEMA_signal_16021 ;
    wire new_AGEMA_signal_16022 ;
    wire new_AGEMA_signal_16023 ;
    wire new_AGEMA_signal_16024 ;
    wire new_AGEMA_signal_16025 ;
    wire new_AGEMA_signal_16026 ;
    wire new_AGEMA_signal_16027 ;
    wire new_AGEMA_signal_16028 ;
    wire new_AGEMA_signal_16029 ;
    wire new_AGEMA_signal_16030 ;
    wire new_AGEMA_signal_16031 ;
    wire new_AGEMA_signal_16032 ;
    wire new_AGEMA_signal_16033 ;
    wire new_AGEMA_signal_16034 ;
    wire new_AGEMA_signal_16035 ;
    wire new_AGEMA_signal_16036 ;
    wire new_AGEMA_signal_16037 ;
    wire new_AGEMA_signal_16038 ;
    wire new_AGEMA_signal_16039 ;
    wire new_AGEMA_signal_16040 ;
    wire new_AGEMA_signal_16041 ;
    wire new_AGEMA_signal_16042 ;
    wire new_AGEMA_signal_16043 ;
    wire new_AGEMA_signal_16044 ;
    wire new_AGEMA_signal_16045 ;
    wire new_AGEMA_signal_16046 ;
    wire new_AGEMA_signal_16047 ;
    wire new_AGEMA_signal_16048 ;
    wire new_AGEMA_signal_16049 ;
    wire new_AGEMA_signal_16050 ;
    wire new_AGEMA_signal_16051 ;
    wire new_AGEMA_signal_16052 ;
    wire new_AGEMA_signal_16053 ;
    wire new_AGEMA_signal_16054 ;
    wire new_AGEMA_signal_16055 ;
    wire new_AGEMA_signal_16056 ;
    wire new_AGEMA_signal_16057 ;
    wire new_AGEMA_signal_16058 ;
    wire new_AGEMA_signal_16059 ;
    wire new_AGEMA_signal_16060 ;
    wire new_AGEMA_signal_16061 ;
    wire new_AGEMA_signal_16062 ;
    wire new_AGEMA_signal_16063 ;
    wire new_AGEMA_signal_16064 ;
    wire new_AGEMA_signal_16065 ;
    wire new_AGEMA_signal_16066 ;
    wire new_AGEMA_signal_16067 ;
    wire new_AGEMA_signal_16068 ;
    wire new_AGEMA_signal_16069 ;
    wire new_AGEMA_signal_16070 ;
    wire new_AGEMA_signal_16071 ;
    wire new_AGEMA_signal_16072 ;
    wire new_AGEMA_signal_16073 ;
    wire new_AGEMA_signal_16074 ;
    wire new_AGEMA_signal_16075 ;
    wire new_AGEMA_signal_16076 ;
    wire new_AGEMA_signal_16077 ;
    wire new_AGEMA_signal_16078 ;
    wire new_AGEMA_signal_16079 ;
    wire new_AGEMA_signal_16080 ;
    wire new_AGEMA_signal_16081 ;
    wire new_AGEMA_signal_16082 ;
    wire new_AGEMA_signal_16083 ;
    wire new_AGEMA_signal_16084 ;
    wire new_AGEMA_signal_16085 ;
    wire new_AGEMA_signal_16086 ;
    wire new_AGEMA_signal_16087 ;
    wire new_AGEMA_signal_16088 ;
    wire new_AGEMA_signal_16089 ;
    wire new_AGEMA_signal_16090 ;
    wire new_AGEMA_signal_16091 ;
    wire new_AGEMA_signal_16092 ;
    wire new_AGEMA_signal_16093 ;
    wire new_AGEMA_signal_16094 ;
    wire new_AGEMA_signal_16095 ;
    wire new_AGEMA_signal_16096 ;
    wire new_AGEMA_signal_16097 ;
    wire new_AGEMA_signal_16098 ;
    wire new_AGEMA_signal_16099 ;
    wire new_AGEMA_signal_16100 ;
    wire new_AGEMA_signal_16101 ;
    wire new_AGEMA_signal_16102 ;
    wire new_AGEMA_signal_16103 ;
    wire new_AGEMA_signal_16104 ;
    wire new_AGEMA_signal_16105 ;
    wire new_AGEMA_signal_16106 ;
    wire new_AGEMA_signal_16107 ;
    wire new_AGEMA_signal_16108 ;
    wire new_AGEMA_signal_16109 ;
    wire new_AGEMA_signal_16110 ;
    wire new_AGEMA_signal_16111 ;
    wire new_AGEMA_signal_16112 ;
    wire new_AGEMA_signal_16113 ;
    wire new_AGEMA_signal_16114 ;
    wire new_AGEMA_signal_16115 ;
    wire new_AGEMA_signal_16116 ;
    wire new_AGEMA_signal_16117 ;
    wire new_AGEMA_signal_16118 ;
    wire new_AGEMA_signal_16119 ;
    wire new_AGEMA_signal_16120 ;
    wire new_AGEMA_signal_16121 ;
    wire new_AGEMA_signal_16122 ;
    wire new_AGEMA_signal_16123 ;
    wire new_AGEMA_signal_16124 ;
    wire new_AGEMA_signal_16125 ;
    wire new_AGEMA_signal_16126 ;
    wire new_AGEMA_signal_16127 ;
    wire new_AGEMA_signal_16128 ;
    wire new_AGEMA_signal_16129 ;
    wire new_AGEMA_signal_16130 ;
    wire new_AGEMA_signal_16131 ;
    wire new_AGEMA_signal_16132 ;
    wire new_AGEMA_signal_16133 ;
    wire new_AGEMA_signal_16134 ;
    wire new_AGEMA_signal_16135 ;
    wire new_AGEMA_signal_16136 ;
    wire new_AGEMA_signal_16137 ;
    wire new_AGEMA_signal_16138 ;
    wire new_AGEMA_signal_16139 ;
    wire new_AGEMA_signal_16140 ;
    wire new_AGEMA_signal_16141 ;
    wire new_AGEMA_signal_16142 ;
    wire new_AGEMA_signal_16143 ;
    wire new_AGEMA_signal_16144 ;
    wire new_AGEMA_signal_16145 ;
    wire new_AGEMA_signal_16146 ;
    wire new_AGEMA_signal_16147 ;
    wire new_AGEMA_signal_16148 ;
    wire new_AGEMA_signal_16149 ;
    wire new_AGEMA_signal_16150 ;
    wire new_AGEMA_signal_16151 ;
    wire new_AGEMA_signal_16152 ;
    wire new_AGEMA_signal_16153 ;
    wire new_AGEMA_signal_16154 ;
    wire new_AGEMA_signal_16155 ;
    wire new_AGEMA_signal_16156 ;
    wire new_AGEMA_signal_16157 ;
    wire new_AGEMA_signal_16158 ;
    wire new_AGEMA_signal_16159 ;
    wire new_AGEMA_signal_16160 ;
    wire new_AGEMA_signal_16161 ;
    wire new_AGEMA_signal_16162 ;
    wire new_AGEMA_signal_16163 ;
    wire new_AGEMA_signal_16164 ;
    wire new_AGEMA_signal_16165 ;
    wire new_AGEMA_signal_16166 ;
    wire new_AGEMA_signal_16167 ;
    wire new_AGEMA_signal_16168 ;
    wire new_AGEMA_signal_16169 ;
    wire new_AGEMA_signal_16170 ;
    wire new_AGEMA_signal_16171 ;
    wire new_AGEMA_signal_16172 ;
    wire new_AGEMA_signal_16173 ;
    wire new_AGEMA_signal_16174 ;
    wire new_AGEMA_signal_16175 ;
    wire new_AGEMA_signal_16176 ;
    wire new_AGEMA_signal_16177 ;
    wire new_AGEMA_signal_16178 ;
    wire new_AGEMA_signal_16179 ;
    wire new_AGEMA_signal_16180 ;
    wire new_AGEMA_signal_16181 ;
    wire new_AGEMA_signal_16182 ;
    wire new_AGEMA_signal_16183 ;
    wire new_AGEMA_signal_16184 ;
    wire new_AGEMA_signal_16185 ;
    wire new_AGEMA_signal_16186 ;
    wire new_AGEMA_signal_16187 ;
    wire new_AGEMA_signal_16188 ;
    wire new_AGEMA_signal_16189 ;
    wire new_AGEMA_signal_16190 ;
    wire new_AGEMA_signal_16191 ;
    wire new_AGEMA_signal_16192 ;
    wire new_AGEMA_signal_16193 ;
    wire new_AGEMA_signal_16194 ;
    wire new_AGEMA_signal_16195 ;
    wire new_AGEMA_signal_16199 ;
    wire new_AGEMA_signal_16200 ;
    wire new_AGEMA_signal_16201 ;
    wire new_AGEMA_signal_16205 ;
    wire new_AGEMA_signal_16206 ;
    wire new_AGEMA_signal_16207 ;
    wire new_AGEMA_signal_16211 ;
    wire new_AGEMA_signal_16212 ;
    wire new_AGEMA_signal_16213 ;
    wire new_AGEMA_signal_16214 ;
    wire new_AGEMA_signal_16215 ;
    wire new_AGEMA_signal_16216 ;
    wire new_AGEMA_signal_16220 ;
    wire new_AGEMA_signal_16221 ;
    wire new_AGEMA_signal_16222 ;
    wire new_AGEMA_signal_16226 ;
    wire new_AGEMA_signal_16227 ;
    wire new_AGEMA_signal_16228 ;
    wire new_AGEMA_signal_16232 ;
    wire new_AGEMA_signal_16233 ;
    wire new_AGEMA_signal_16234 ;
    wire new_AGEMA_signal_16238 ;
    wire new_AGEMA_signal_16239 ;
    wire new_AGEMA_signal_16240 ;
    wire new_AGEMA_signal_16244 ;
    wire new_AGEMA_signal_16245 ;
    wire new_AGEMA_signal_16246 ;
    wire new_AGEMA_signal_16250 ;
    wire new_AGEMA_signal_16251 ;
    wire new_AGEMA_signal_16252 ;
    wire new_AGEMA_signal_16256 ;
    wire new_AGEMA_signal_16257 ;
    wire new_AGEMA_signal_16258 ;
    wire new_AGEMA_signal_16259 ;
    wire new_AGEMA_signal_16260 ;
    wire new_AGEMA_signal_16261 ;
    wire new_AGEMA_signal_16265 ;
    wire new_AGEMA_signal_16266 ;
    wire new_AGEMA_signal_16267 ;
    wire new_AGEMA_signal_16271 ;
    wire new_AGEMA_signal_16272 ;
    wire new_AGEMA_signal_16273 ;
    wire new_AGEMA_signal_16277 ;
    wire new_AGEMA_signal_16278 ;
    wire new_AGEMA_signal_16279 ;
    wire new_AGEMA_signal_16283 ;
    wire new_AGEMA_signal_16284 ;
    wire new_AGEMA_signal_16285 ;
    wire new_AGEMA_signal_16289 ;
    wire new_AGEMA_signal_16290 ;
    wire new_AGEMA_signal_16291 ;
    wire new_AGEMA_signal_16295 ;
    wire new_AGEMA_signal_16296 ;
    wire new_AGEMA_signal_16297 ;
    wire new_AGEMA_signal_16301 ;
    wire new_AGEMA_signal_16302 ;
    wire new_AGEMA_signal_16303 ;
    wire new_AGEMA_signal_16304 ;
    wire new_AGEMA_signal_16305 ;
    wire new_AGEMA_signal_16306 ;
    wire new_AGEMA_signal_16310 ;
    wire new_AGEMA_signal_16311 ;
    wire new_AGEMA_signal_16312 ;
    wire new_AGEMA_signal_16316 ;
    wire new_AGEMA_signal_16317 ;
    wire new_AGEMA_signal_16318 ;
    wire new_AGEMA_signal_16322 ;
    wire new_AGEMA_signal_16323 ;
    wire new_AGEMA_signal_16324 ;
    wire new_AGEMA_signal_16328 ;
    wire new_AGEMA_signal_16329 ;
    wire new_AGEMA_signal_16330 ;
    wire new_AGEMA_signal_16334 ;
    wire new_AGEMA_signal_16335 ;
    wire new_AGEMA_signal_16336 ;
    wire new_AGEMA_signal_16340 ;
    wire new_AGEMA_signal_16341 ;
    wire new_AGEMA_signal_16342 ;
    wire new_AGEMA_signal_16346 ;
    wire new_AGEMA_signal_16347 ;
    wire new_AGEMA_signal_16348 ;
    wire new_AGEMA_signal_16352 ;
    wire new_AGEMA_signal_16353 ;
    wire new_AGEMA_signal_16354 ;
    wire new_AGEMA_signal_16355 ;
    wire new_AGEMA_signal_16356 ;
    wire new_AGEMA_signal_16357 ;
    wire new_AGEMA_signal_16358 ;
    wire new_AGEMA_signal_16359 ;
    wire new_AGEMA_signal_16360 ;
    wire new_AGEMA_signal_16361 ;
    wire new_AGEMA_signal_16362 ;
    wire new_AGEMA_signal_16363 ;
    wire new_AGEMA_signal_16364 ;
    wire new_AGEMA_signal_16365 ;
    wire new_AGEMA_signal_16366 ;
    wire new_AGEMA_signal_16367 ;
    wire new_AGEMA_signal_16368 ;
    wire new_AGEMA_signal_16369 ;
    wire new_AGEMA_signal_16370 ;
    wire new_AGEMA_signal_16371 ;
    wire new_AGEMA_signal_16372 ;
    wire new_AGEMA_signal_16373 ;
    wire new_AGEMA_signal_16374 ;
    wire new_AGEMA_signal_16375 ;
    wire new_AGEMA_signal_16376 ;
    wire new_AGEMA_signal_16377 ;
    wire new_AGEMA_signal_16378 ;
    wire new_AGEMA_signal_16379 ;
    wire new_AGEMA_signal_16380 ;
    wire new_AGEMA_signal_16381 ;
    wire new_AGEMA_signal_16382 ;
    wire new_AGEMA_signal_16383 ;
    wire new_AGEMA_signal_16384 ;
    wire new_AGEMA_signal_16385 ;
    wire new_AGEMA_signal_16386 ;
    wire new_AGEMA_signal_16387 ;
    wire new_AGEMA_signal_16388 ;
    wire new_AGEMA_signal_16389 ;
    wire new_AGEMA_signal_16390 ;
    wire new_AGEMA_signal_16391 ;
    wire new_AGEMA_signal_16392 ;
    wire new_AGEMA_signal_16393 ;
    wire new_AGEMA_signal_16394 ;
    wire new_AGEMA_signal_16395 ;
    wire new_AGEMA_signal_16396 ;
    wire new_AGEMA_signal_16397 ;
    wire new_AGEMA_signal_16398 ;
    wire new_AGEMA_signal_16399 ;
    wire new_AGEMA_signal_16400 ;
    wire new_AGEMA_signal_16401 ;
    wire new_AGEMA_signal_16402 ;
    wire new_AGEMA_signal_16403 ;
    wire new_AGEMA_signal_16404 ;
    wire new_AGEMA_signal_16405 ;
    wire new_AGEMA_signal_16406 ;
    wire new_AGEMA_signal_16407 ;
    wire new_AGEMA_signal_16408 ;
    wire new_AGEMA_signal_16409 ;
    wire new_AGEMA_signal_16410 ;
    wire new_AGEMA_signal_16411 ;
    wire new_AGEMA_signal_16412 ;
    wire new_AGEMA_signal_16413 ;
    wire new_AGEMA_signal_16414 ;
    wire new_AGEMA_signal_16415 ;
    wire new_AGEMA_signal_16416 ;
    wire new_AGEMA_signal_16417 ;
    wire new_AGEMA_signal_16418 ;
    wire new_AGEMA_signal_16419 ;
    wire new_AGEMA_signal_16420 ;
    wire new_AGEMA_signal_16424 ;
    wire new_AGEMA_signal_16425 ;
    wire new_AGEMA_signal_16426 ;
    wire new_AGEMA_signal_16430 ;
    wire new_AGEMA_signal_16431 ;
    wire new_AGEMA_signal_16432 ;
    wire new_AGEMA_signal_16436 ;
    wire new_AGEMA_signal_16437 ;
    wire new_AGEMA_signal_16438 ;
    wire new_AGEMA_signal_16442 ;
    wire new_AGEMA_signal_16443 ;
    wire new_AGEMA_signal_16444 ;
    wire new_AGEMA_signal_16448 ;
    wire new_AGEMA_signal_16449 ;
    wire new_AGEMA_signal_16450 ;
    wire new_AGEMA_signal_16454 ;
    wire new_AGEMA_signal_16455 ;
    wire new_AGEMA_signal_16456 ;
    wire new_AGEMA_signal_16460 ;
    wire new_AGEMA_signal_16461 ;
    wire new_AGEMA_signal_16462 ;
    wire new_AGEMA_signal_16463 ;
    wire new_AGEMA_signal_16464 ;
    wire new_AGEMA_signal_16465 ;
    wire new_AGEMA_signal_16466 ;
    wire new_AGEMA_signal_16467 ;
    wire new_AGEMA_signal_16468 ;
    wire new_AGEMA_signal_16469 ;
    wire new_AGEMA_signal_16470 ;
    wire new_AGEMA_signal_16471 ;
    wire new_AGEMA_signal_16472 ;
    wire new_AGEMA_signal_16473 ;
    wire new_AGEMA_signal_16474 ;
    wire new_AGEMA_signal_16475 ;
    wire new_AGEMA_signal_16476 ;
    wire new_AGEMA_signal_16477 ;
    wire new_AGEMA_signal_16478 ;
    wire new_AGEMA_signal_16479 ;
    wire new_AGEMA_signal_16480 ;
    wire new_AGEMA_signal_16481 ;
    wire new_AGEMA_signal_16482 ;
    wire new_AGEMA_signal_16483 ;
    wire new_AGEMA_signal_16484 ;
    wire new_AGEMA_signal_16485 ;
    wire new_AGEMA_signal_16486 ;
    wire new_AGEMA_signal_16487 ;
    wire new_AGEMA_signal_16488 ;
    wire new_AGEMA_signal_16489 ;
    wire new_AGEMA_signal_16490 ;
    wire new_AGEMA_signal_16491 ;
    wire new_AGEMA_signal_16492 ;
    wire new_AGEMA_signal_16493 ;
    wire new_AGEMA_signal_16494 ;
    wire new_AGEMA_signal_16495 ;
    wire new_AGEMA_signal_16496 ;
    wire new_AGEMA_signal_16497 ;
    wire new_AGEMA_signal_16498 ;
    wire new_AGEMA_signal_16499 ;
    wire new_AGEMA_signal_16500 ;
    wire new_AGEMA_signal_16501 ;
    wire new_AGEMA_signal_16502 ;
    wire new_AGEMA_signal_16503 ;
    wire new_AGEMA_signal_16504 ;
    wire new_AGEMA_signal_16505 ;
    wire new_AGEMA_signal_16506 ;
    wire new_AGEMA_signal_16507 ;
    wire new_AGEMA_signal_16508 ;
    wire new_AGEMA_signal_16509 ;
    wire new_AGEMA_signal_16510 ;
    wire new_AGEMA_signal_16511 ;
    wire new_AGEMA_signal_16512 ;
    wire new_AGEMA_signal_16513 ;
    wire new_AGEMA_signal_16514 ;
    wire new_AGEMA_signal_16515 ;
    wire new_AGEMA_signal_16516 ;
    wire new_AGEMA_signal_16517 ;
    wire new_AGEMA_signal_16518 ;
    wire new_AGEMA_signal_16519 ;
    wire new_AGEMA_signal_16520 ;
    wire new_AGEMA_signal_16521 ;
    wire new_AGEMA_signal_16522 ;
    wire new_AGEMA_signal_16523 ;
    wire new_AGEMA_signal_16524 ;
    wire new_AGEMA_signal_16525 ;
    wire new_AGEMA_signal_16526 ;
    wire new_AGEMA_signal_16527 ;
    wire new_AGEMA_signal_16528 ;
    wire new_AGEMA_signal_16529 ;
    wire new_AGEMA_signal_16530 ;
    wire new_AGEMA_signal_16531 ;
    wire new_AGEMA_signal_16532 ;
    wire new_AGEMA_signal_16533 ;
    wire new_AGEMA_signal_16534 ;
    wire new_AGEMA_signal_16535 ;
    wire new_AGEMA_signal_16536 ;
    wire new_AGEMA_signal_16537 ;
    wire new_AGEMA_signal_16538 ;
    wire new_AGEMA_signal_16539 ;
    wire new_AGEMA_signal_16540 ;
    wire new_AGEMA_signal_16541 ;
    wire new_AGEMA_signal_16542 ;
    wire new_AGEMA_signal_16543 ;
    wire new_AGEMA_signal_16544 ;
    wire new_AGEMA_signal_16545 ;
    wire new_AGEMA_signal_16546 ;
    wire new_AGEMA_signal_16547 ;
    wire new_AGEMA_signal_16548 ;
    wire new_AGEMA_signal_16549 ;
    wire new_AGEMA_signal_16550 ;
    wire new_AGEMA_signal_16551 ;
    wire new_AGEMA_signal_16552 ;
    wire new_AGEMA_signal_16553 ;
    wire new_AGEMA_signal_16554 ;
    wire new_AGEMA_signal_16555 ;
    wire new_AGEMA_signal_16556 ;
    wire new_AGEMA_signal_16557 ;
    wire new_AGEMA_signal_16558 ;
    wire new_AGEMA_signal_16559 ;
    wire new_AGEMA_signal_16560 ;
    wire new_AGEMA_signal_16561 ;
    wire new_AGEMA_signal_16562 ;
    wire new_AGEMA_signal_16563 ;
    wire new_AGEMA_signal_16564 ;
    wire new_AGEMA_signal_16565 ;
    wire new_AGEMA_signal_16566 ;
    wire new_AGEMA_signal_16567 ;
    wire new_AGEMA_signal_16568 ;
    wire new_AGEMA_signal_16569 ;
    wire new_AGEMA_signal_16570 ;
    wire new_AGEMA_signal_16571 ;
    wire new_AGEMA_signal_16572 ;
    wire new_AGEMA_signal_16573 ;
    wire new_AGEMA_signal_16574 ;
    wire new_AGEMA_signal_16575 ;
    wire new_AGEMA_signal_16576 ;
    wire new_AGEMA_signal_16577 ;
    wire new_AGEMA_signal_16578 ;
    wire new_AGEMA_signal_16579 ;
    wire new_AGEMA_signal_16580 ;
    wire new_AGEMA_signal_16581 ;
    wire new_AGEMA_signal_16582 ;
    wire new_AGEMA_signal_16583 ;
    wire new_AGEMA_signal_16584 ;
    wire new_AGEMA_signal_16585 ;
    wire new_AGEMA_signal_16586 ;
    wire new_AGEMA_signal_16587 ;
    wire new_AGEMA_signal_16588 ;
    wire new_AGEMA_signal_16589 ;
    wire new_AGEMA_signal_16590 ;
    wire new_AGEMA_signal_16591 ;
    wire new_AGEMA_signal_16592 ;
    wire new_AGEMA_signal_16593 ;
    wire new_AGEMA_signal_16594 ;
    wire new_AGEMA_signal_16595 ;
    wire new_AGEMA_signal_16596 ;
    wire new_AGEMA_signal_16597 ;
    wire new_AGEMA_signal_16598 ;
    wire new_AGEMA_signal_16599 ;
    wire new_AGEMA_signal_16600 ;
    wire new_AGEMA_signal_16601 ;
    wire new_AGEMA_signal_16602 ;
    wire new_AGEMA_signal_16603 ;
    wire new_AGEMA_signal_16604 ;
    wire new_AGEMA_signal_16605 ;
    wire new_AGEMA_signal_16606 ;
    wire new_AGEMA_signal_16607 ;
    wire new_AGEMA_signal_16608 ;
    wire new_AGEMA_signal_16609 ;
    wire new_AGEMA_signal_16610 ;
    wire new_AGEMA_signal_16611 ;
    wire new_AGEMA_signal_16612 ;
    wire new_AGEMA_signal_16613 ;
    wire new_AGEMA_signal_16614 ;
    wire new_AGEMA_signal_16615 ;
    wire new_AGEMA_signal_16616 ;
    wire new_AGEMA_signal_16617 ;
    wire new_AGEMA_signal_16618 ;
    wire new_AGEMA_signal_16619 ;
    wire new_AGEMA_signal_16620 ;
    wire new_AGEMA_signal_16621 ;
    wire new_AGEMA_signal_16622 ;
    wire new_AGEMA_signal_16623 ;
    wire new_AGEMA_signal_16624 ;
    wire new_AGEMA_signal_16625 ;
    wire new_AGEMA_signal_16626 ;
    wire new_AGEMA_signal_16627 ;
    wire new_AGEMA_signal_16628 ;
    wire new_AGEMA_signal_16629 ;
    wire new_AGEMA_signal_16630 ;
    wire new_AGEMA_signal_16631 ;
    wire new_AGEMA_signal_16632 ;
    wire new_AGEMA_signal_16633 ;
    wire new_AGEMA_signal_16634 ;
    wire new_AGEMA_signal_16635 ;
    wire new_AGEMA_signal_16636 ;
    wire new_AGEMA_signal_16637 ;
    wire new_AGEMA_signal_16638 ;
    wire new_AGEMA_signal_16639 ;
    wire new_AGEMA_signal_16640 ;
    wire new_AGEMA_signal_16641 ;
    wire new_AGEMA_signal_16642 ;
    wire new_AGEMA_signal_16643 ;
    wire new_AGEMA_signal_16644 ;
    wire new_AGEMA_signal_16645 ;
    wire new_AGEMA_signal_16646 ;
    wire new_AGEMA_signal_16647 ;
    wire new_AGEMA_signal_16648 ;
    wire new_AGEMA_signal_16649 ;
    wire new_AGEMA_signal_16650 ;
    wire new_AGEMA_signal_16651 ;
    wire new_AGEMA_signal_16652 ;
    wire new_AGEMA_signal_16653 ;
    wire new_AGEMA_signal_16654 ;
    wire new_AGEMA_signal_16655 ;
    wire new_AGEMA_signal_16656 ;
    wire new_AGEMA_signal_16657 ;
    wire new_AGEMA_signal_16658 ;
    wire new_AGEMA_signal_16659 ;
    wire new_AGEMA_signal_16660 ;
    wire new_AGEMA_signal_16661 ;
    wire new_AGEMA_signal_16662 ;
    wire new_AGEMA_signal_16663 ;
    wire new_AGEMA_signal_16664 ;
    wire new_AGEMA_signal_16665 ;
    wire new_AGEMA_signal_16666 ;
    wire new_AGEMA_signal_16667 ;
    wire new_AGEMA_signal_16668 ;
    wire new_AGEMA_signal_16669 ;
    wire new_AGEMA_signal_16670 ;
    wire new_AGEMA_signal_16671 ;
    wire new_AGEMA_signal_16672 ;
    wire new_AGEMA_signal_16673 ;
    wire new_AGEMA_signal_16674 ;
    wire new_AGEMA_signal_16675 ;
    wire new_AGEMA_signal_16676 ;
    wire new_AGEMA_signal_16677 ;
    wire new_AGEMA_signal_16678 ;
    wire new_AGEMA_signal_16679 ;
    wire new_AGEMA_signal_16680 ;
    wire new_AGEMA_signal_16681 ;
    wire new_AGEMA_signal_16682 ;
    wire new_AGEMA_signal_16683 ;
    wire new_AGEMA_signal_16684 ;
    wire new_AGEMA_signal_16685 ;
    wire new_AGEMA_signal_16686 ;
    wire new_AGEMA_signal_16687 ;
    wire new_AGEMA_signal_16688 ;
    wire new_AGEMA_signal_16689 ;
    wire new_AGEMA_signal_16690 ;
    wire new_AGEMA_signal_16691 ;
    wire new_AGEMA_signal_16692 ;
    wire new_AGEMA_signal_16693 ;
    wire new_AGEMA_signal_16694 ;
    wire new_AGEMA_signal_16695 ;
    wire new_AGEMA_signal_16696 ;
    wire new_AGEMA_signal_16697 ;
    wire new_AGEMA_signal_16698 ;
    wire new_AGEMA_signal_16699 ;
    wire new_AGEMA_signal_16700 ;
    wire new_AGEMA_signal_16701 ;
    wire new_AGEMA_signal_16702 ;
    wire new_AGEMA_signal_16703 ;
    wire new_AGEMA_signal_16704 ;
    wire new_AGEMA_signal_16705 ;
    wire new_AGEMA_signal_16706 ;
    wire new_AGEMA_signal_16707 ;
    wire new_AGEMA_signal_16708 ;
    wire new_AGEMA_signal_16709 ;
    wire new_AGEMA_signal_16710 ;
    wire new_AGEMA_signal_16711 ;
    wire new_AGEMA_signal_16712 ;
    wire new_AGEMA_signal_16713 ;
    wire new_AGEMA_signal_16714 ;
    wire new_AGEMA_signal_16715 ;
    wire new_AGEMA_signal_16716 ;
    wire new_AGEMA_signal_16717 ;
    wire new_AGEMA_signal_16718 ;
    wire new_AGEMA_signal_16719 ;
    wire new_AGEMA_signal_16720 ;
    wire new_AGEMA_signal_16721 ;
    wire new_AGEMA_signal_16722 ;
    wire new_AGEMA_signal_16723 ;
    wire new_AGEMA_signal_16724 ;
    wire new_AGEMA_signal_16725 ;
    wire new_AGEMA_signal_16726 ;
    wire new_AGEMA_signal_16727 ;
    wire new_AGEMA_signal_16728 ;
    wire new_AGEMA_signal_16729 ;
    wire new_AGEMA_signal_16730 ;
    wire new_AGEMA_signal_16731 ;
    wire new_AGEMA_signal_16732 ;
    wire new_AGEMA_signal_16733 ;
    wire new_AGEMA_signal_16734 ;
    wire new_AGEMA_signal_16735 ;
    wire new_AGEMA_signal_16736 ;
    wire new_AGEMA_signal_16737 ;
    wire new_AGEMA_signal_16738 ;
    wire new_AGEMA_signal_16739 ;
    wire new_AGEMA_signal_16740 ;
    wire new_AGEMA_signal_16741 ;
    wire new_AGEMA_signal_16742 ;
    wire new_AGEMA_signal_16743 ;
    wire new_AGEMA_signal_16744 ;
    wire new_AGEMA_signal_16745 ;
    wire new_AGEMA_signal_16746 ;
    wire new_AGEMA_signal_16747 ;
    wire new_AGEMA_signal_16748 ;
    wire new_AGEMA_signal_16749 ;
    wire new_AGEMA_signal_16750 ;
    wire new_AGEMA_signal_16751 ;
    wire new_AGEMA_signal_16752 ;
    wire new_AGEMA_signal_16753 ;
    wire new_AGEMA_signal_16754 ;
    wire new_AGEMA_signal_16755 ;
    wire new_AGEMA_signal_16756 ;
    wire new_AGEMA_signal_16757 ;
    wire new_AGEMA_signal_16758 ;
    wire new_AGEMA_signal_16759 ;
    wire new_AGEMA_signal_16760 ;
    wire new_AGEMA_signal_16761 ;
    wire new_AGEMA_signal_16762 ;
    wire new_AGEMA_signal_16763 ;
    wire new_AGEMA_signal_16764 ;
    wire new_AGEMA_signal_16765 ;
    wire new_AGEMA_signal_16766 ;
    wire new_AGEMA_signal_16767 ;
    wire new_AGEMA_signal_16768 ;
    wire new_AGEMA_signal_16769 ;
    wire new_AGEMA_signal_16770 ;
    wire new_AGEMA_signal_16771 ;
    wire new_AGEMA_signal_16772 ;
    wire new_AGEMA_signal_16773 ;
    wire new_AGEMA_signal_16774 ;
    wire new_AGEMA_signal_16775 ;
    wire new_AGEMA_signal_16776 ;
    wire new_AGEMA_signal_16777 ;
    wire new_AGEMA_signal_16778 ;
    wire new_AGEMA_signal_16779 ;
    wire new_AGEMA_signal_16780 ;
    wire new_AGEMA_signal_16781 ;
    wire new_AGEMA_signal_16782 ;
    wire new_AGEMA_signal_16783 ;
    wire new_AGEMA_signal_16784 ;
    wire new_AGEMA_signal_16785 ;
    wire new_AGEMA_signal_16786 ;
    wire new_AGEMA_signal_16787 ;
    wire new_AGEMA_signal_16788 ;
    wire new_AGEMA_signal_16789 ;
    wire new_AGEMA_signal_16790 ;
    wire new_AGEMA_signal_16791 ;
    wire new_AGEMA_signal_16792 ;
    wire new_AGEMA_signal_16793 ;
    wire new_AGEMA_signal_16794 ;
    wire new_AGEMA_signal_16795 ;
    wire new_AGEMA_signal_16796 ;
    wire new_AGEMA_signal_16797 ;
    wire new_AGEMA_signal_16798 ;
    wire new_AGEMA_signal_16799 ;
    wire new_AGEMA_signal_16800 ;
    wire new_AGEMA_signal_16801 ;
    wire new_AGEMA_signal_16802 ;
    wire new_AGEMA_signal_16803 ;
    wire new_AGEMA_signal_16804 ;
    wire new_AGEMA_signal_16805 ;
    wire new_AGEMA_signal_16806 ;
    wire new_AGEMA_signal_16807 ;
    wire new_AGEMA_signal_16808 ;
    wire new_AGEMA_signal_16809 ;
    wire new_AGEMA_signal_16810 ;
    wire new_AGEMA_signal_16811 ;
    wire new_AGEMA_signal_16812 ;
    wire new_AGEMA_signal_16813 ;
    wire new_AGEMA_signal_16814 ;
    wire new_AGEMA_signal_16815 ;
    wire new_AGEMA_signal_16816 ;
    wire new_AGEMA_signal_16817 ;
    wire new_AGEMA_signal_16818 ;
    wire new_AGEMA_signal_16819 ;
    wire new_AGEMA_signal_16820 ;
    wire new_AGEMA_signal_16821 ;
    wire new_AGEMA_signal_16822 ;
    wire new_AGEMA_signal_16823 ;
    wire new_AGEMA_signal_16824 ;
    wire new_AGEMA_signal_16825 ;
    wire new_AGEMA_signal_16826 ;
    wire new_AGEMA_signal_16827 ;
    wire new_AGEMA_signal_16828 ;
    wire new_AGEMA_signal_16829 ;
    wire new_AGEMA_signal_16830 ;
    wire new_AGEMA_signal_16831 ;
    wire new_AGEMA_signal_16832 ;
    wire new_AGEMA_signal_16833 ;
    wire new_AGEMA_signal_16834 ;
    wire new_AGEMA_signal_16835 ;
    wire new_AGEMA_signal_16836 ;
    wire new_AGEMA_signal_16837 ;
    wire new_AGEMA_signal_16838 ;
    wire new_AGEMA_signal_16839 ;
    wire new_AGEMA_signal_16840 ;
    wire new_AGEMA_signal_16841 ;
    wire new_AGEMA_signal_16842 ;
    wire new_AGEMA_signal_16843 ;
    wire new_AGEMA_signal_16844 ;
    wire new_AGEMA_signal_16845 ;
    wire new_AGEMA_signal_16846 ;
    wire new_AGEMA_signal_16847 ;
    wire new_AGEMA_signal_16848 ;
    wire new_AGEMA_signal_16849 ;
    wire new_AGEMA_signal_16850 ;
    wire new_AGEMA_signal_16851 ;
    wire new_AGEMA_signal_16852 ;
    wire new_AGEMA_signal_16853 ;
    wire new_AGEMA_signal_16854 ;
    wire new_AGEMA_signal_16855 ;
    wire new_AGEMA_signal_16856 ;
    wire new_AGEMA_signal_16857 ;
    wire new_AGEMA_signal_16858 ;
    wire new_AGEMA_signal_16859 ;
    wire new_AGEMA_signal_16860 ;
    wire new_AGEMA_signal_16861 ;
    wire new_AGEMA_signal_16862 ;
    wire new_AGEMA_signal_16863 ;
    wire new_AGEMA_signal_16864 ;
    wire new_AGEMA_signal_16865 ;
    wire new_AGEMA_signal_16866 ;
    wire new_AGEMA_signal_16867 ;
    wire new_AGEMA_signal_16868 ;
    wire new_AGEMA_signal_16869 ;
    wire new_AGEMA_signal_16870 ;
    wire new_AGEMA_signal_16871 ;
    wire new_AGEMA_signal_16872 ;
    wire new_AGEMA_signal_16873 ;
    wire new_AGEMA_signal_16874 ;
    wire new_AGEMA_signal_16875 ;
    wire new_AGEMA_signal_16876 ;
    wire new_AGEMA_signal_16877 ;
    wire new_AGEMA_signal_16878 ;
    wire new_AGEMA_signal_16879 ;
    wire new_AGEMA_signal_16880 ;
    wire new_AGEMA_signal_16881 ;
    wire new_AGEMA_signal_16882 ;
    wire new_AGEMA_signal_16883 ;
    wire new_AGEMA_signal_16884 ;
    wire new_AGEMA_signal_16885 ;
    wire new_AGEMA_signal_16886 ;
    wire new_AGEMA_signal_16887 ;
    wire new_AGEMA_signal_16888 ;
    wire new_AGEMA_signal_16889 ;
    wire new_AGEMA_signal_16890 ;
    wire new_AGEMA_signal_16891 ;
    wire new_AGEMA_signal_16892 ;
    wire new_AGEMA_signal_16893 ;
    wire new_AGEMA_signal_16894 ;
    wire new_AGEMA_signal_16895 ;
    wire new_AGEMA_signal_16896 ;
    wire new_AGEMA_signal_16897 ;
    wire new_AGEMA_signal_16898 ;
    wire new_AGEMA_signal_16899 ;
    wire new_AGEMA_signal_16900 ;
    wire new_AGEMA_signal_16901 ;
    wire new_AGEMA_signal_16902 ;
    wire new_AGEMA_signal_16903 ;
    wire new_AGEMA_signal_16904 ;
    wire new_AGEMA_signal_16905 ;
    wire new_AGEMA_signal_16906 ;
    wire new_AGEMA_signal_16907 ;
    wire new_AGEMA_signal_16908 ;
    wire new_AGEMA_signal_16909 ;
    wire new_AGEMA_signal_16910 ;
    wire new_AGEMA_signal_16911 ;
    wire new_AGEMA_signal_16912 ;
    wire new_AGEMA_signal_16913 ;
    wire new_AGEMA_signal_16914 ;
    wire new_AGEMA_signal_16915 ;
    wire new_AGEMA_signal_16916 ;
    wire new_AGEMA_signal_16917 ;
    wire new_AGEMA_signal_16918 ;
    wire new_AGEMA_signal_16919 ;
    wire new_AGEMA_signal_16920 ;
    wire new_AGEMA_signal_16921 ;
    wire new_AGEMA_signal_16922 ;
    wire new_AGEMA_signal_16923 ;
    wire new_AGEMA_signal_16924 ;
    wire new_AGEMA_signal_16925 ;
    wire new_AGEMA_signal_16926 ;
    wire new_AGEMA_signal_16927 ;
    wire new_AGEMA_signal_16928 ;
    wire new_AGEMA_signal_16929 ;
    wire new_AGEMA_signal_16930 ;
    wire new_AGEMA_signal_16931 ;
    wire new_AGEMA_signal_16932 ;
    wire new_AGEMA_signal_16933 ;
    wire new_AGEMA_signal_16934 ;
    wire new_AGEMA_signal_16935 ;
    wire new_AGEMA_signal_16936 ;
    wire new_AGEMA_signal_16937 ;
    wire new_AGEMA_signal_16938 ;
    wire new_AGEMA_signal_16939 ;
    wire new_AGEMA_signal_16940 ;
    wire new_AGEMA_signal_16941 ;
    wire new_AGEMA_signal_16942 ;
    wire new_AGEMA_signal_16943 ;
    wire new_AGEMA_signal_16944 ;
    wire new_AGEMA_signal_16945 ;
    wire new_AGEMA_signal_16946 ;
    wire new_AGEMA_signal_16947 ;
    wire new_AGEMA_signal_16948 ;
    wire new_AGEMA_signal_16949 ;
    wire new_AGEMA_signal_16950 ;
    wire new_AGEMA_signal_16951 ;
    wire new_AGEMA_signal_16952 ;
    wire new_AGEMA_signal_16953 ;
    wire new_AGEMA_signal_16954 ;
    wire new_AGEMA_signal_16955 ;
    wire new_AGEMA_signal_16956 ;
    wire new_AGEMA_signal_16957 ;
    wire new_AGEMA_signal_16961 ;
    wire new_AGEMA_signal_16962 ;
    wire new_AGEMA_signal_16963 ;
    wire new_AGEMA_signal_16967 ;
    wire new_AGEMA_signal_16968 ;
    wire new_AGEMA_signal_16969 ;
    wire new_AGEMA_signal_16973 ;
    wire new_AGEMA_signal_16974 ;
    wire new_AGEMA_signal_16975 ;
    wire new_AGEMA_signal_16979 ;
    wire new_AGEMA_signal_16980 ;
    wire new_AGEMA_signal_16981 ;
    wire new_AGEMA_signal_16985 ;
    wire new_AGEMA_signal_16986 ;
    wire new_AGEMA_signal_16987 ;
    wire new_AGEMA_signal_16991 ;
    wire new_AGEMA_signal_16992 ;
    wire new_AGEMA_signal_16993 ;
    wire new_AGEMA_signal_16997 ;
    wire new_AGEMA_signal_16998 ;
    wire new_AGEMA_signal_16999 ;
    wire new_AGEMA_signal_17000 ;
    wire new_AGEMA_signal_17001 ;
    wire new_AGEMA_signal_17002 ;
    wire new_AGEMA_signal_17006 ;
    wire new_AGEMA_signal_17007 ;
    wire new_AGEMA_signal_17008 ;
    wire new_AGEMA_signal_17012 ;
    wire new_AGEMA_signal_17013 ;
    wire new_AGEMA_signal_17014 ;
    wire new_AGEMA_signal_17018 ;
    wire new_AGEMA_signal_17019 ;
    wire new_AGEMA_signal_17020 ;
    wire new_AGEMA_signal_17024 ;
    wire new_AGEMA_signal_17025 ;
    wire new_AGEMA_signal_17026 ;
    wire new_AGEMA_signal_17030 ;
    wire new_AGEMA_signal_17031 ;
    wire new_AGEMA_signal_17032 ;
    wire new_AGEMA_signal_17036 ;
    wire new_AGEMA_signal_17037 ;
    wire new_AGEMA_signal_17038 ;
    wire new_AGEMA_signal_17042 ;
    wire new_AGEMA_signal_17043 ;
    wire new_AGEMA_signal_17044 ;
    wire new_AGEMA_signal_17045 ;
    wire new_AGEMA_signal_17046 ;
    wire new_AGEMA_signal_17047 ;
    wire new_AGEMA_signal_17051 ;
    wire new_AGEMA_signal_17052 ;
    wire new_AGEMA_signal_17053 ;
    wire new_AGEMA_signal_17057 ;
    wire new_AGEMA_signal_17058 ;
    wire new_AGEMA_signal_17059 ;
    wire new_AGEMA_signal_17063 ;
    wire new_AGEMA_signal_17064 ;
    wire new_AGEMA_signal_17065 ;
    wire new_AGEMA_signal_17069 ;
    wire new_AGEMA_signal_17070 ;
    wire new_AGEMA_signal_17071 ;
    wire new_AGEMA_signal_17075 ;
    wire new_AGEMA_signal_17076 ;
    wire new_AGEMA_signal_17077 ;
    wire new_AGEMA_signal_17081 ;
    wire new_AGEMA_signal_17082 ;
    wire new_AGEMA_signal_17083 ;
    wire new_AGEMA_signal_17087 ;
    wire new_AGEMA_signal_17088 ;
    wire new_AGEMA_signal_17089 ;
    wire new_AGEMA_signal_17093 ;
    wire new_AGEMA_signal_17094 ;
    wire new_AGEMA_signal_17095 ;
    wire new_AGEMA_signal_17096 ;
    wire new_AGEMA_signal_17097 ;
    wire new_AGEMA_signal_17098 ;
    wire new_AGEMA_signal_17099 ;
    wire new_AGEMA_signal_17100 ;
    wire new_AGEMA_signal_17101 ;
    wire new_AGEMA_signal_17102 ;
    wire new_AGEMA_signal_17103 ;
    wire new_AGEMA_signal_17104 ;
    wire new_AGEMA_signal_17105 ;
    wire new_AGEMA_signal_17106 ;
    wire new_AGEMA_signal_17107 ;
    wire new_AGEMA_signal_17108 ;
    wire new_AGEMA_signal_17109 ;
    wire new_AGEMA_signal_17110 ;
    wire new_AGEMA_signal_17111 ;
    wire new_AGEMA_signal_17112 ;
    wire new_AGEMA_signal_17113 ;
    wire new_AGEMA_signal_17114 ;
    wire new_AGEMA_signal_17115 ;
    wire new_AGEMA_signal_17116 ;
    wire new_AGEMA_signal_17117 ;
    wire new_AGEMA_signal_17118 ;
    wire new_AGEMA_signal_17119 ;
    wire new_AGEMA_signal_17120 ;
    wire new_AGEMA_signal_17121 ;
    wire new_AGEMA_signal_17122 ;
    wire new_AGEMA_signal_17123 ;
    wire new_AGEMA_signal_17124 ;
    wire new_AGEMA_signal_17125 ;
    wire new_AGEMA_signal_17126 ;
    wire new_AGEMA_signal_17127 ;
    wire new_AGEMA_signal_17128 ;
    wire new_AGEMA_signal_17129 ;
    wire new_AGEMA_signal_17130 ;
    wire new_AGEMA_signal_17131 ;
    wire new_AGEMA_signal_17132 ;
    wire new_AGEMA_signal_17133 ;
    wire new_AGEMA_signal_17134 ;
    wire new_AGEMA_signal_17135 ;
    wire new_AGEMA_signal_17136 ;
    wire new_AGEMA_signal_17137 ;
    wire new_AGEMA_signal_17138 ;
    wire new_AGEMA_signal_17139 ;
    wire new_AGEMA_signal_17140 ;
    wire new_AGEMA_signal_17141 ;
    wire new_AGEMA_signal_17142 ;
    wire new_AGEMA_signal_17143 ;
    wire new_AGEMA_signal_17144 ;
    wire new_AGEMA_signal_17145 ;
    wire new_AGEMA_signal_17146 ;
    wire new_AGEMA_signal_17147 ;
    wire new_AGEMA_signal_17148 ;
    wire new_AGEMA_signal_17149 ;
    wire new_AGEMA_signal_17150 ;
    wire new_AGEMA_signal_17151 ;
    wire new_AGEMA_signal_17152 ;
    wire new_AGEMA_signal_17153 ;
    wire new_AGEMA_signal_17154 ;
    wire new_AGEMA_signal_17155 ;
    wire new_AGEMA_signal_17156 ;
    wire new_AGEMA_signal_17157 ;
    wire new_AGEMA_signal_17158 ;
    wire new_AGEMA_signal_17159 ;
    wire new_AGEMA_signal_17160 ;
    wire new_AGEMA_signal_17161 ;
    wire new_AGEMA_signal_17165 ;
    wire new_AGEMA_signal_17166 ;
    wire new_AGEMA_signal_17167 ;
    wire new_AGEMA_signal_17171 ;
    wire new_AGEMA_signal_17172 ;
    wire new_AGEMA_signal_17173 ;
    wire new_AGEMA_signal_17177 ;
    wire new_AGEMA_signal_17178 ;
    wire new_AGEMA_signal_17179 ;
    wire new_AGEMA_signal_17183 ;
    wire new_AGEMA_signal_17184 ;
    wire new_AGEMA_signal_17185 ;
    wire new_AGEMA_signal_17189 ;
    wire new_AGEMA_signal_17190 ;
    wire new_AGEMA_signal_17191 ;
    wire new_AGEMA_signal_17195 ;
    wire new_AGEMA_signal_17196 ;
    wire new_AGEMA_signal_17197 ;
    wire new_AGEMA_signal_17201 ;
    wire new_AGEMA_signal_17202 ;
    wire new_AGEMA_signal_17203 ;
    wire new_AGEMA_signal_17204 ;
    wire new_AGEMA_signal_17205 ;
    wire new_AGEMA_signal_17206 ;
    wire new_AGEMA_signal_17207 ;
    wire new_AGEMA_signal_17208 ;
    wire new_AGEMA_signal_17209 ;
    wire new_AGEMA_signal_17210 ;
    wire new_AGEMA_signal_17211 ;
    wire new_AGEMA_signal_17212 ;
    wire new_AGEMA_signal_17213 ;
    wire new_AGEMA_signal_17214 ;
    wire new_AGEMA_signal_17215 ;
    wire new_AGEMA_signal_17216 ;
    wire new_AGEMA_signal_17217 ;
    wire new_AGEMA_signal_17218 ;
    wire new_AGEMA_signal_17219 ;
    wire new_AGEMA_signal_17220 ;
    wire new_AGEMA_signal_17221 ;
    wire new_AGEMA_signal_17222 ;
    wire new_AGEMA_signal_17223 ;
    wire new_AGEMA_signal_17224 ;
    wire new_AGEMA_signal_17225 ;
    wire new_AGEMA_signal_17226 ;
    wire new_AGEMA_signal_17227 ;
    wire new_AGEMA_signal_17228 ;
    wire new_AGEMA_signal_17229 ;
    wire new_AGEMA_signal_17230 ;
    wire new_AGEMA_signal_17231 ;
    wire new_AGEMA_signal_17232 ;
    wire new_AGEMA_signal_17233 ;
    wire new_AGEMA_signal_17234 ;
    wire new_AGEMA_signal_17235 ;
    wire new_AGEMA_signal_17236 ;
    wire new_AGEMA_signal_17237 ;
    wire new_AGEMA_signal_17238 ;
    wire new_AGEMA_signal_17239 ;
    wire new_AGEMA_signal_17240 ;
    wire new_AGEMA_signal_17241 ;
    wire new_AGEMA_signal_17242 ;
    wire new_AGEMA_signal_17243 ;
    wire new_AGEMA_signal_17244 ;
    wire new_AGEMA_signal_17245 ;
    wire new_AGEMA_signal_17246 ;
    wire new_AGEMA_signal_17247 ;
    wire new_AGEMA_signal_17248 ;
    wire new_AGEMA_signal_17249 ;
    wire new_AGEMA_signal_17250 ;
    wire new_AGEMA_signal_17251 ;
    wire new_AGEMA_signal_17252 ;
    wire new_AGEMA_signal_17253 ;
    wire new_AGEMA_signal_17254 ;
    wire new_AGEMA_signal_17255 ;
    wire new_AGEMA_signal_17256 ;
    wire new_AGEMA_signal_17257 ;
    wire new_AGEMA_signal_17258 ;
    wire new_AGEMA_signal_17259 ;
    wire new_AGEMA_signal_17260 ;
    wire new_AGEMA_signal_17261 ;
    wire new_AGEMA_signal_17262 ;
    wire new_AGEMA_signal_17263 ;
    wire new_AGEMA_signal_17264 ;
    wire new_AGEMA_signal_17265 ;
    wire new_AGEMA_signal_17266 ;
    wire new_AGEMA_signal_17267 ;
    wire new_AGEMA_signal_17268 ;
    wire new_AGEMA_signal_17269 ;
    wire new_AGEMA_signal_17270 ;
    wire new_AGEMA_signal_17271 ;
    wire new_AGEMA_signal_17272 ;
    wire new_AGEMA_signal_17273 ;
    wire new_AGEMA_signal_17274 ;
    wire new_AGEMA_signal_17275 ;
    wire new_AGEMA_signal_17276 ;
    wire new_AGEMA_signal_17277 ;
    wire new_AGEMA_signal_17278 ;
    wire new_AGEMA_signal_17279 ;
    wire new_AGEMA_signal_17280 ;
    wire new_AGEMA_signal_17281 ;
    wire new_AGEMA_signal_17282 ;
    wire new_AGEMA_signal_17283 ;
    wire new_AGEMA_signal_17284 ;
    wire new_AGEMA_signal_17285 ;
    wire new_AGEMA_signal_17286 ;
    wire new_AGEMA_signal_17287 ;
    wire new_AGEMA_signal_17288 ;
    wire new_AGEMA_signal_17289 ;
    wire new_AGEMA_signal_17290 ;
    wire new_AGEMA_signal_17291 ;
    wire new_AGEMA_signal_17292 ;
    wire new_AGEMA_signal_17293 ;
    wire new_AGEMA_signal_17294 ;
    wire new_AGEMA_signal_17295 ;
    wire new_AGEMA_signal_17296 ;
    wire new_AGEMA_signal_17297 ;
    wire new_AGEMA_signal_17298 ;
    wire new_AGEMA_signal_17299 ;
    wire new_AGEMA_signal_17300 ;
    wire new_AGEMA_signal_17301 ;
    wire new_AGEMA_signal_17302 ;
    wire new_AGEMA_signal_17303 ;
    wire new_AGEMA_signal_17304 ;
    wire new_AGEMA_signal_17305 ;
    wire new_AGEMA_signal_17306 ;
    wire new_AGEMA_signal_17307 ;
    wire new_AGEMA_signal_17308 ;
    wire new_AGEMA_signal_17309 ;
    wire new_AGEMA_signal_17310 ;
    wire new_AGEMA_signal_17311 ;
    wire new_AGEMA_signal_17312 ;
    wire new_AGEMA_signal_17313 ;
    wire new_AGEMA_signal_17314 ;
    wire new_AGEMA_signal_17315 ;
    wire new_AGEMA_signal_17316 ;
    wire new_AGEMA_signal_17317 ;
    wire new_AGEMA_signal_17318 ;
    wire new_AGEMA_signal_17319 ;
    wire new_AGEMA_signal_17320 ;
    wire new_AGEMA_signal_17321 ;
    wire new_AGEMA_signal_17322 ;
    wire new_AGEMA_signal_17323 ;
    wire new_AGEMA_signal_17324 ;
    wire new_AGEMA_signal_17325 ;
    wire new_AGEMA_signal_17326 ;
    wire new_AGEMA_signal_17327 ;
    wire new_AGEMA_signal_17328 ;
    wire new_AGEMA_signal_17329 ;
    wire new_AGEMA_signal_17330 ;
    wire new_AGEMA_signal_17331 ;
    wire new_AGEMA_signal_17332 ;
    wire new_AGEMA_signal_17333 ;
    wire new_AGEMA_signal_17334 ;
    wire new_AGEMA_signal_17335 ;
    wire new_AGEMA_signal_17336 ;
    wire new_AGEMA_signal_17337 ;
    wire new_AGEMA_signal_17338 ;
    wire new_AGEMA_signal_17339 ;
    wire new_AGEMA_signal_17340 ;
    wire new_AGEMA_signal_17341 ;
    wire new_AGEMA_signal_17342 ;
    wire new_AGEMA_signal_17343 ;
    wire new_AGEMA_signal_17344 ;
    wire new_AGEMA_signal_17345 ;
    wire new_AGEMA_signal_17346 ;
    wire new_AGEMA_signal_17347 ;
    wire new_AGEMA_signal_17348 ;
    wire new_AGEMA_signal_17349 ;
    wire new_AGEMA_signal_17350 ;
    wire new_AGEMA_signal_17351 ;
    wire new_AGEMA_signal_17352 ;
    wire new_AGEMA_signal_17353 ;
    wire new_AGEMA_signal_17354 ;
    wire new_AGEMA_signal_17355 ;
    wire new_AGEMA_signal_17356 ;
    wire new_AGEMA_signal_17357 ;
    wire new_AGEMA_signal_17358 ;
    wire new_AGEMA_signal_17359 ;
    wire new_AGEMA_signal_17360 ;
    wire new_AGEMA_signal_17361 ;
    wire new_AGEMA_signal_17362 ;
    wire new_AGEMA_signal_17363 ;
    wire new_AGEMA_signal_17364 ;
    wire new_AGEMA_signal_17365 ;
    wire new_AGEMA_signal_17366 ;
    wire new_AGEMA_signal_17367 ;
    wire new_AGEMA_signal_17368 ;
    wire new_AGEMA_signal_17369 ;
    wire new_AGEMA_signal_17370 ;
    wire new_AGEMA_signal_17371 ;
    wire new_AGEMA_signal_17372 ;
    wire new_AGEMA_signal_17373 ;
    wire new_AGEMA_signal_17374 ;
    wire new_AGEMA_signal_17375 ;
    wire new_AGEMA_signal_17376 ;
    wire new_AGEMA_signal_17377 ;
    wire new_AGEMA_signal_17378 ;
    wire new_AGEMA_signal_17379 ;
    wire new_AGEMA_signal_17380 ;
    wire new_AGEMA_signal_17381 ;
    wire new_AGEMA_signal_17382 ;
    wire new_AGEMA_signal_17383 ;
    wire new_AGEMA_signal_17384 ;
    wire new_AGEMA_signal_17385 ;
    wire new_AGEMA_signal_17386 ;
    wire new_AGEMA_signal_17387 ;
    wire new_AGEMA_signal_17388 ;
    wire new_AGEMA_signal_17389 ;
    wire new_AGEMA_signal_17390 ;
    wire new_AGEMA_signal_17391 ;
    wire new_AGEMA_signal_17392 ;
    wire new_AGEMA_signal_17393 ;
    wire new_AGEMA_signal_17394 ;
    wire new_AGEMA_signal_17395 ;
    wire new_AGEMA_signal_17396 ;
    wire new_AGEMA_signal_17397 ;
    wire new_AGEMA_signal_17398 ;
    wire new_AGEMA_signal_17399 ;
    wire new_AGEMA_signal_17400 ;
    wire new_AGEMA_signal_17401 ;
    wire new_AGEMA_signal_17402 ;
    wire new_AGEMA_signal_17403 ;
    wire new_AGEMA_signal_17404 ;
    wire new_AGEMA_signal_17405 ;
    wire new_AGEMA_signal_17406 ;
    wire new_AGEMA_signal_17407 ;
    wire new_AGEMA_signal_17408 ;
    wire new_AGEMA_signal_17409 ;
    wire new_AGEMA_signal_17410 ;
    wire new_AGEMA_signal_17411 ;
    wire new_AGEMA_signal_17412 ;
    wire new_AGEMA_signal_17413 ;
    wire new_AGEMA_signal_17414 ;
    wire new_AGEMA_signal_17415 ;
    wire new_AGEMA_signal_17416 ;
    wire new_AGEMA_signal_17417 ;
    wire new_AGEMA_signal_17418 ;
    wire new_AGEMA_signal_17419 ;
    wire new_AGEMA_signal_17420 ;
    wire new_AGEMA_signal_17421 ;
    wire new_AGEMA_signal_17422 ;
    wire new_AGEMA_signal_17423 ;
    wire new_AGEMA_signal_17424 ;
    wire new_AGEMA_signal_17425 ;
    wire new_AGEMA_signal_17426 ;
    wire new_AGEMA_signal_17427 ;
    wire new_AGEMA_signal_17428 ;
    wire new_AGEMA_signal_17429 ;
    wire new_AGEMA_signal_17430 ;
    wire new_AGEMA_signal_17431 ;
    wire new_AGEMA_signal_17432 ;
    wire new_AGEMA_signal_17433 ;
    wire new_AGEMA_signal_17434 ;
    wire new_AGEMA_signal_17435 ;
    wire new_AGEMA_signal_17436 ;
    wire new_AGEMA_signal_17437 ;
    wire new_AGEMA_signal_17438 ;
    wire new_AGEMA_signal_17439 ;
    wire new_AGEMA_signal_17440 ;
    wire new_AGEMA_signal_17441 ;
    wire new_AGEMA_signal_17442 ;
    wire new_AGEMA_signal_17443 ;
    wire new_AGEMA_signal_17444 ;
    wire new_AGEMA_signal_17445 ;
    wire new_AGEMA_signal_17446 ;
    wire new_AGEMA_signal_17447 ;
    wire new_AGEMA_signal_17448 ;
    wire new_AGEMA_signal_17449 ;
    wire new_AGEMA_signal_17450 ;
    wire new_AGEMA_signal_17451 ;
    wire new_AGEMA_signal_17452 ;
    wire new_AGEMA_signal_17453 ;
    wire new_AGEMA_signal_17454 ;
    wire new_AGEMA_signal_17455 ;
    wire new_AGEMA_signal_17456 ;
    wire new_AGEMA_signal_17457 ;
    wire new_AGEMA_signal_17458 ;
    wire new_AGEMA_signal_17459 ;
    wire new_AGEMA_signal_17460 ;
    wire new_AGEMA_signal_17461 ;
    wire new_AGEMA_signal_17462 ;
    wire new_AGEMA_signal_17463 ;
    wire new_AGEMA_signal_17464 ;
    wire new_AGEMA_signal_17465 ;
    wire new_AGEMA_signal_17466 ;
    wire new_AGEMA_signal_17467 ;
    wire new_AGEMA_signal_17468 ;
    wire new_AGEMA_signal_17469 ;
    wire new_AGEMA_signal_17470 ;
    wire new_AGEMA_signal_17471 ;
    wire new_AGEMA_signal_17472 ;
    wire new_AGEMA_signal_17473 ;
    wire new_AGEMA_signal_17474 ;
    wire new_AGEMA_signal_17475 ;
    wire new_AGEMA_signal_17476 ;
    wire new_AGEMA_signal_17477 ;
    wire new_AGEMA_signal_17478 ;
    wire new_AGEMA_signal_17479 ;
    wire new_AGEMA_signal_17480 ;
    wire new_AGEMA_signal_17481 ;
    wire new_AGEMA_signal_17482 ;
    wire new_AGEMA_signal_17483 ;
    wire new_AGEMA_signal_17484 ;
    wire new_AGEMA_signal_17485 ;
    wire new_AGEMA_signal_17486 ;
    wire new_AGEMA_signal_17487 ;
    wire new_AGEMA_signal_17488 ;
    wire new_AGEMA_signal_17489 ;
    wire new_AGEMA_signal_17490 ;
    wire new_AGEMA_signal_17491 ;
    wire new_AGEMA_signal_17492 ;
    wire new_AGEMA_signal_17493 ;
    wire new_AGEMA_signal_17494 ;
    wire new_AGEMA_signal_17495 ;
    wire new_AGEMA_signal_17496 ;
    wire new_AGEMA_signal_17497 ;
    wire new_AGEMA_signal_17498 ;
    wire new_AGEMA_signal_17499 ;
    wire new_AGEMA_signal_17500 ;
    wire new_AGEMA_signal_17501 ;
    wire new_AGEMA_signal_17502 ;
    wire new_AGEMA_signal_17503 ;
    wire new_AGEMA_signal_17504 ;
    wire new_AGEMA_signal_17505 ;
    wire new_AGEMA_signal_17506 ;
    wire new_AGEMA_signal_17507 ;
    wire new_AGEMA_signal_17508 ;
    wire new_AGEMA_signal_17509 ;
    wire new_AGEMA_signal_17510 ;
    wire new_AGEMA_signal_17511 ;
    wire new_AGEMA_signal_17512 ;
    wire new_AGEMA_signal_17513 ;
    wire new_AGEMA_signal_17514 ;
    wire new_AGEMA_signal_17515 ;
    wire new_AGEMA_signal_17516 ;
    wire new_AGEMA_signal_17517 ;
    wire new_AGEMA_signal_17518 ;
    wire new_AGEMA_signal_17519 ;
    wire new_AGEMA_signal_17520 ;
    wire new_AGEMA_signal_17521 ;
    wire new_AGEMA_signal_17522 ;
    wire new_AGEMA_signal_17523 ;
    wire new_AGEMA_signal_17524 ;
    wire new_AGEMA_signal_17525 ;
    wire new_AGEMA_signal_17526 ;
    wire new_AGEMA_signal_17527 ;
    wire new_AGEMA_signal_17528 ;
    wire new_AGEMA_signal_17529 ;
    wire new_AGEMA_signal_17530 ;
    wire new_AGEMA_signal_17531 ;
    wire new_AGEMA_signal_17532 ;
    wire new_AGEMA_signal_17533 ;
    wire new_AGEMA_signal_17534 ;
    wire new_AGEMA_signal_17535 ;
    wire new_AGEMA_signal_17536 ;
    wire new_AGEMA_signal_17537 ;
    wire new_AGEMA_signal_17538 ;
    wire new_AGEMA_signal_17539 ;
    wire new_AGEMA_signal_17540 ;
    wire new_AGEMA_signal_17541 ;
    wire new_AGEMA_signal_17542 ;
    wire new_AGEMA_signal_17543 ;
    wire new_AGEMA_signal_17544 ;
    wire new_AGEMA_signal_17545 ;
    wire new_AGEMA_signal_17546 ;
    wire new_AGEMA_signal_17547 ;
    wire new_AGEMA_signal_17548 ;
    wire new_AGEMA_signal_17549 ;
    wire new_AGEMA_signal_17550 ;
    wire new_AGEMA_signal_17551 ;
    wire new_AGEMA_signal_17552 ;
    wire new_AGEMA_signal_17553 ;
    wire new_AGEMA_signal_17554 ;
    wire new_AGEMA_signal_17555 ;
    wire new_AGEMA_signal_17556 ;
    wire new_AGEMA_signal_17557 ;
    wire new_AGEMA_signal_17558 ;
    wire new_AGEMA_signal_17559 ;
    wire new_AGEMA_signal_17560 ;
    wire new_AGEMA_signal_17561 ;
    wire new_AGEMA_signal_17562 ;
    wire new_AGEMA_signal_17563 ;
    wire new_AGEMA_signal_17564 ;
    wire new_AGEMA_signal_17565 ;
    wire new_AGEMA_signal_17566 ;
    wire new_AGEMA_signal_17567 ;
    wire new_AGEMA_signal_17568 ;
    wire new_AGEMA_signal_17569 ;
    wire new_AGEMA_signal_17570 ;
    wire new_AGEMA_signal_17571 ;
    wire new_AGEMA_signal_17572 ;
    wire new_AGEMA_signal_17573 ;
    wire new_AGEMA_signal_17574 ;
    wire new_AGEMA_signal_17575 ;
    wire new_AGEMA_signal_17576 ;
    wire new_AGEMA_signal_17577 ;
    wire new_AGEMA_signal_17578 ;
    wire new_AGEMA_signal_17579 ;
    wire new_AGEMA_signal_17580 ;
    wire new_AGEMA_signal_17581 ;
    wire new_AGEMA_signal_17582 ;
    wire new_AGEMA_signal_17583 ;
    wire new_AGEMA_signal_17584 ;
    wire new_AGEMA_signal_17585 ;
    wire new_AGEMA_signal_17586 ;
    wire new_AGEMA_signal_17587 ;
    wire new_AGEMA_signal_17588 ;
    wire new_AGEMA_signal_17589 ;
    wire new_AGEMA_signal_17590 ;
    wire new_AGEMA_signal_17591 ;
    wire new_AGEMA_signal_17592 ;
    wire new_AGEMA_signal_17593 ;
    wire new_AGEMA_signal_17594 ;
    wire new_AGEMA_signal_17595 ;
    wire new_AGEMA_signal_17596 ;
    wire new_AGEMA_signal_17597 ;
    wire new_AGEMA_signal_17598 ;
    wire new_AGEMA_signal_17599 ;
    wire new_AGEMA_signal_17600 ;
    wire new_AGEMA_signal_17601 ;
    wire new_AGEMA_signal_17602 ;
    wire new_AGEMA_signal_17603 ;
    wire new_AGEMA_signal_17604 ;
    wire new_AGEMA_signal_17605 ;
    wire new_AGEMA_signal_17606 ;
    wire new_AGEMA_signal_17607 ;
    wire new_AGEMA_signal_17608 ;
    wire new_AGEMA_signal_17609 ;
    wire new_AGEMA_signal_17610 ;
    wire new_AGEMA_signal_17611 ;
    wire new_AGEMA_signal_17612 ;
    wire new_AGEMA_signal_17613 ;
    wire new_AGEMA_signal_17614 ;
    wire new_AGEMA_signal_17615 ;
    wire new_AGEMA_signal_17616 ;
    wire new_AGEMA_signal_17617 ;
    wire new_AGEMA_signal_17618 ;
    wire new_AGEMA_signal_17619 ;
    wire new_AGEMA_signal_17620 ;
    wire new_AGEMA_signal_17621 ;
    wire new_AGEMA_signal_17622 ;
    wire new_AGEMA_signal_17623 ;
    wire new_AGEMA_signal_17624 ;
    wire new_AGEMA_signal_17625 ;
    wire new_AGEMA_signal_17626 ;
    wire new_AGEMA_signal_17627 ;
    wire new_AGEMA_signal_17628 ;
    wire new_AGEMA_signal_17629 ;
    wire new_AGEMA_signal_17630 ;
    wire new_AGEMA_signal_17631 ;
    wire new_AGEMA_signal_17632 ;
    wire new_AGEMA_signal_17633 ;
    wire new_AGEMA_signal_17634 ;
    wire new_AGEMA_signal_17635 ;
    wire new_AGEMA_signal_17636 ;
    wire new_AGEMA_signal_17637 ;
    wire new_AGEMA_signal_17638 ;
    wire new_AGEMA_signal_17639 ;
    wire new_AGEMA_signal_17640 ;
    wire new_AGEMA_signal_17641 ;
    wire new_AGEMA_signal_17642 ;
    wire new_AGEMA_signal_17643 ;
    wire new_AGEMA_signal_17644 ;
    wire new_AGEMA_signal_17645 ;
    wire new_AGEMA_signal_17646 ;
    wire new_AGEMA_signal_17647 ;
    wire new_AGEMA_signal_17648 ;
    wire new_AGEMA_signal_17649 ;
    wire new_AGEMA_signal_17650 ;
    wire new_AGEMA_signal_17651 ;
    wire new_AGEMA_signal_17652 ;
    wire new_AGEMA_signal_17653 ;
    wire new_AGEMA_signal_17654 ;
    wire new_AGEMA_signal_17655 ;
    wire new_AGEMA_signal_17656 ;
    wire new_AGEMA_signal_17657 ;
    wire new_AGEMA_signal_17658 ;
    wire new_AGEMA_signal_17659 ;
    wire new_AGEMA_signal_17660 ;
    wire new_AGEMA_signal_17661 ;
    wire new_AGEMA_signal_17662 ;
    wire new_AGEMA_signal_17663 ;
    wire new_AGEMA_signal_17664 ;
    wire new_AGEMA_signal_17665 ;
    wire new_AGEMA_signal_17666 ;
    wire new_AGEMA_signal_17667 ;
    wire new_AGEMA_signal_17668 ;
    wire new_AGEMA_signal_17669 ;
    wire new_AGEMA_signal_17670 ;
    wire new_AGEMA_signal_17671 ;
    wire new_AGEMA_signal_17672 ;
    wire new_AGEMA_signal_17673 ;
    wire new_AGEMA_signal_17674 ;
    wire new_AGEMA_signal_17675 ;
    wire new_AGEMA_signal_17676 ;
    wire new_AGEMA_signal_17677 ;
    wire new_AGEMA_signal_17678 ;
    wire new_AGEMA_signal_17679 ;
    wire new_AGEMA_signal_17680 ;
    wire new_AGEMA_signal_17681 ;
    wire new_AGEMA_signal_17682 ;
    wire new_AGEMA_signal_17683 ;
    wire new_AGEMA_signal_17684 ;
    wire new_AGEMA_signal_17685 ;
    wire new_AGEMA_signal_17686 ;
    wire new_AGEMA_signal_17687 ;
    wire new_AGEMA_signal_17688 ;
    wire new_AGEMA_signal_17689 ;
    wire new_AGEMA_signal_17690 ;
    wire new_AGEMA_signal_17691 ;
    wire new_AGEMA_signal_17692 ;
    wire new_AGEMA_signal_17693 ;
    wire new_AGEMA_signal_17694 ;
    wire new_AGEMA_signal_17695 ;
    wire new_AGEMA_signal_17699 ;
    wire new_AGEMA_signal_17700 ;
    wire new_AGEMA_signal_17701 ;
    wire new_AGEMA_signal_17705 ;
    wire new_AGEMA_signal_17706 ;
    wire new_AGEMA_signal_17707 ;
    wire new_AGEMA_signal_17711 ;
    wire new_AGEMA_signal_17712 ;
    wire new_AGEMA_signal_17713 ;
    wire new_AGEMA_signal_17717 ;
    wire new_AGEMA_signal_17718 ;
    wire new_AGEMA_signal_17719 ;
    wire new_AGEMA_signal_17723 ;
    wire new_AGEMA_signal_17724 ;
    wire new_AGEMA_signal_17725 ;
    wire new_AGEMA_signal_17729 ;
    wire new_AGEMA_signal_17730 ;
    wire new_AGEMA_signal_17731 ;
    wire new_AGEMA_signal_17735 ;
    wire new_AGEMA_signal_17736 ;
    wire new_AGEMA_signal_17737 ;
    wire new_AGEMA_signal_17738 ;
    wire new_AGEMA_signal_17739 ;
    wire new_AGEMA_signal_17740 ;
    wire new_AGEMA_signal_17741 ;
    wire new_AGEMA_signal_17742 ;
    wire new_AGEMA_signal_17743 ;
    wire new_AGEMA_signal_17744 ;
    wire new_AGEMA_signal_17745 ;
    wire new_AGEMA_signal_17746 ;
    wire new_AGEMA_signal_17747 ;
    wire new_AGEMA_signal_17748 ;
    wire new_AGEMA_signal_17749 ;
    wire new_AGEMA_signal_17750 ;
    wire new_AGEMA_signal_17751 ;
    wire new_AGEMA_signal_17752 ;
    wire new_AGEMA_signal_17753 ;
    wire new_AGEMA_signal_17754 ;
    wire new_AGEMA_signal_17755 ;
    wire new_AGEMA_signal_17756 ;
    wire new_AGEMA_signal_17757 ;
    wire new_AGEMA_signal_17758 ;
    wire new_AGEMA_signal_17759 ;
    wire new_AGEMA_signal_17760 ;
    wire new_AGEMA_signal_17761 ;
    wire new_AGEMA_signal_17762 ;
    wire new_AGEMA_signal_17763 ;
    wire new_AGEMA_signal_17764 ;
    wire new_AGEMA_signal_17765 ;
    wire new_AGEMA_signal_17766 ;
    wire new_AGEMA_signal_17767 ;
    wire new_AGEMA_signal_17768 ;
    wire new_AGEMA_signal_17769 ;
    wire new_AGEMA_signal_17770 ;
    wire new_AGEMA_signal_17771 ;
    wire new_AGEMA_signal_17772 ;
    wire new_AGEMA_signal_17773 ;
    wire new_AGEMA_signal_17774 ;
    wire new_AGEMA_signal_17775 ;
    wire new_AGEMA_signal_17776 ;
    wire new_AGEMA_signal_17777 ;
    wire new_AGEMA_signal_17778 ;
    wire new_AGEMA_signal_17779 ;
    wire new_AGEMA_signal_17780 ;
    wire new_AGEMA_signal_17781 ;
    wire new_AGEMA_signal_17782 ;
    wire new_AGEMA_signal_17783 ;
    wire new_AGEMA_signal_17784 ;
    wire new_AGEMA_signal_17785 ;
    wire new_AGEMA_signal_17786 ;
    wire new_AGEMA_signal_17787 ;
    wire new_AGEMA_signal_17788 ;
    wire new_AGEMA_signal_17789 ;
    wire new_AGEMA_signal_17790 ;
    wire new_AGEMA_signal_17791 ;
    wire new_AGEMA_signal_17792 ;
    wire new_AGEMA_signal_17793 ;
    wire new_AGEMA_signal_17794 ;
    wire new_AGEMA_signal_17795 ;
    wire new_AGEMA_signal_17796 ;
    wire new_AGEMA_signal_17797 ;
    wire new_AGEMA_signal_17798 ;
    wire new_AGEMA_signal_17799 ;
    wire new_AGEMA_signal_17800 ;
    wire new_AGEMA_signal_17801 ;
    wire new_AGEMA_signal_17802 ;
    wire new_AGEMA_signal_17803 ;
    wire new_AGEMA_signal_17804 ;
    wire new_AGEMA_signal_17805 ;
    wire new_AGEMA_signal_17806 ;
    wire new_AGEMA_signal_17807 ;
    wire new_AGEMA_signal_17808 ;
    wire new_AGEMA_signal_17809 ;
    wire new_AGEMA_signal_17810 ;
    wire new_AGEMA_signal_17811 ;
    wire new_AGEMA_signal_17812 ;
    wire new_AGEMA_signal_17813 ;
    wire new_AGEMA_signal_17814 ;
    wire new_AGEMA_signal_17815 ;
    wire new_AGEMA_signal_17816 ;
    wire new_AGEMA_signal_17817 ;
    wire new_AGEMA_signal_17818 ;
    wire new_AGEMA_signal_17819 ;
    wire new_AGEMA_signal_17820 ;
    wire new_AGEMA_signal_17821 ;
    wire new_AGEMA_signal_17822 ;
    wire new_AGEMA_signal_17823 ;
    wire new_AGEMA_signal_17824 ;
    wire new_AGEMA_signal_17825 ;
    wire new_AGEMA_signal_17826 ;
    wire new_AGEMA_signal_17827 ;
    wire new_AGEMA_signal_17828 ;
    wire new_AGEMA_signal_17829 ;
    wire new_AGEMA_signal_17830 ;
    wire new_AGEMA_signal_17831 ;
    wire new_AGEMA_signal_17832 ;
    wire new_AGEMA_signal_17833 ;
    wire new_AGEMA_signal_17834 ;
    wire new_AGEMA_signal_17835 ;
    wire new_AGEMA_signal_17836 ;
    wire new_AGEMA_signal_17837 ;
    wire new_AGEMA_signal_17838 ;
    wire new_AGEMA_signal_17839 ;
    wire new_AGEMA_signal_17840 ;
    wire new_AGEMA_signal_17841 ;
    wire new_AGEMA_signal_17842 ;
    wire new_AGEMA_signal_17843 ;
    wire new_AGEMA_signal_17844 ;
    wire new_AGEMA_signal_17845 ;
    wire new_AGEMA_signal_17846 ;
    wire new_AGEMA_signal_17847 ;
    wire new_AGEMA_signal_17848 ;
    wire new_AGEMA_signal_17849 ;
    wire new_AGEMA_signal_17850 ;
    wire new_AGEMA_signal_17851 ;
    wire new_AGEMA_signal_17852 ;
    wire new_AGEMA_signal_17853 ;
    wire new_AGEMA_signal_17854 ;
    wire new_AGEMA_signal_17855 ;
    wire new_AGEMA_signal_17856 ;
    wire new_AGEMA_signal_17857 ;
    wire new_AGEMA_signal_17858 ;
    wire new_AGEMA_signal_17859 ;
    wire new_AGEMA_signal_17860 ;
    wire new_AGEMA_signal_17861 ;
    wire new_AGEMA_signal_17862 ;
    wire new_AGEMA_signal_17863 ;
    wire new_AGEMA_signal_17864 ;
    wire new_AGEMA_signal_17865 ;
    wire new_AGEMA_signal_17866 ;
    wire new_AGEMA_signal_17867 ;
    wire new_AGEMA_signal_17868 ;
    wire new_AGEMA_signal_17869 ;
    wire new_AGEMA_signal_17870 ;
    wire new_AGEMA_signal_17871 ;
    wire new_AGEMA_signal_17872 ;
    wire new_AGEMA_signal_17873 ;
    wire new_AGEMA_signal_17874 ;
    wire new_AGEMA_signal_17875 ;
    wire new_AGEMA_signal_17876 ;
    wire new_AGEMA_signal_17877 ;
    wire new_AGEMA_signal_17878 ;
    wire new_AGEMA_signal_17879 ;
    wire new_AGEMA_signal_17880 ;
    wire new_AGEMA_signal_17881 ;
    wire new_AGEMA_signal_17882 ;
    wire new_AGEMA_signal_17883 ;
    wire new_AGEMA_signal_17884 ;
    wire new_AGEMA_signal_17885 ;
    wire new_AGEMA_signal_17886 ;
    wire new_AGEMA_signal_17887 ;
    wire new_AGEMA_signal_17888 ;
    wire new_AGEMA_signal_17889 ;
    wire new_AGEMA_signal_17890 ;
    wire new_AGEMA_signal_17891 ;
    wire new_AGEMA_signal_17892 ;
    wire new_AGEMA_signal_17893 ;
    wire new_AGEMA_signal_17894 ;
    wire new_AGEMA_signal_17895 ;
    wire new_AGEMA_signal_17896 ;
    wire new_AGEMA_signal_17897 ;
    wire new_AGEMA_signal_17898 ;
    wire new_AGEMA_signal_17899 ;
    wire new_AGEMA_signal_17900 ;
    wire new_AGEMA_signal_17901 ;
    wire new_AGEMA_signal_17902 ;
    wire new_AGEMA_signal_17906 ;
    wire new_AGEMA_signal_17907 ;
    wire new_AGEMA_signal_17908 ;
    wire new_AGEMA_signal_17912 ;
    wire new_AGEMA_signal_17913 ;
    wire new_AGEMA_signal_17914 ;
    wire new_AGEMA_signal_17918 ;
    wire new_AGEMA_signal_17919 ;
    wire new_AGEMA_signal_17920 ;
    wire new_AGEMA_signal_17924 ;
    wire new_AGEMA_signal_17925 ;
    wire new_AGEMA_signal_17926 ;
    wire new_AGEMA_signal_17930 ;
    wire new_AGEMA_signal_17931 ;
    wire new_AGEMA_signal_17932 ;
    wire new_AGEMA_signal_17936 ;
    wire new_AGEMA_signal_17937 ;
    wire new_AGEMA_signal_17938 ;
    wire new_AGEMA_signal_17942 ;
    wire new_AGEMA_signal_17943 ;
    wire new_AGEMA_signal_17944 ;
    wire new_AGEMA_signal_17948 ;
    wire new_AGEMA_signal_17949 ;
    wire new_AGEMA_signal_17950 ;
    wire new_AGEMA_signal_17954 ;
    wire new_AGEMA_signal_17955 ;
    wire new_AGEMA_signal_17956 ;
    wire new_AGEMA_signal_17960 ;
    wire new_AGEMA_signal_17961 ;
    wire new_AGEMA_signal_17962 ;
    wire new_AGEMA_signal_17966 ;
    wire new_AGEMA_signal_17967 ;
    wire new_AGEMA_signal_17968 ;
    wire new_AGEMA_signal_17972 ;
    wire new_AGEMA_signal_17973 ;
    wire new_AGEMA_signal_17974 ;
    wire new_AGEMA_signal_17978 ;
    wire new_AGEMA_signal_17979 ;
    wire new_AGEMA_signal_17980 ;
    wire new_AGEMA_signal_17984 ;
    wire new_AGEMA_signal_17985 ;
    wire new_AGEMA_signal_17986 ;
    wire new_AGEMA_signal_17990 ;
    wire new_AGEMA_signal_17991 ;
    wire new_AGEMA_signal_17992 ;
    wire new_AGEMA_signal_17996 ;
    wire new_AGEMA_signal_17997 ;
    wire new_AGEMA_signal_17998 ;
    wire new_AGEMA_signal_18002 ;
    wire new_AGEMA_signal_18003 ;
    wire new_AGEMA_signal_18004 ;
    wire new_AGEMA_signal_18008 ;
    wire new_AGEMA_signal_18009 ;
    wire new_AGEMA_signal_18010 ;
    wire new_AGEMA_signal_18014 ;
    wire new_AGEMA_signal_18015 ;
    wire new_AGEMA_signal_18016 ;
    wire new_AGEMA_signal_18020 ;
    wire new_AGEMA_signal_18021 ;
    wire new_AGEMA_signal_18022 ;
    wire new_AGEMA_signal_18026 ;
    wire new_AGEMA_signal_18027 ;
    wire new_AGEMA_signal_18028 ;
    wire new_AGEMA_signal_18032 ;
    wire new_AGEMA_signal_18033 ;
    wire new_AGEMA_signal_18034 ;
    wire new_AGEMA_signal_18038 ;
    wire new_AGEMA_signal_18039 ;
    wire new_AGEMA_signal_18040 ;
    wire new_AGEMA_signal_18044 ;
    wire new_AGEMA_signal_18045 ;
    wire new_AGEMA_signal_18046 ;
    wire new_AGEMA_signal_18050 ;
    wire new_AGEMA_signal_18051 ;
    wire new_AGEMA_signal_18052 ;
    wire new_AGEMA_signal_18056 ;
    wire new_AGEMA_signal_18057 ;
    wire new_AGEMA_signal_18058 ;
    wire new_AGEMA_signal_18062 ;
    wire new_AGEMA_signal_18063 ;
    wire new_AGEMA_signal_18064 ;
    wire new_AGEMA_signal_18068 ;
    wire new_AGEMA_signal_18069 ;
    wire new_AGEMA_signal_18070 ;
    wire new_AGEMA_signal_18074 ;
    wire new_AGEMA_signal_18075 ;
    wire new_AGEMA_signal_18076 ;
    wire new_AGEMA_signal_18080 ;
    wire new_AGEMA_signal_18081 ;
    wire new_AGEMA_signal_18082 ;
    wire new_AGEMA_signal_18086 ;
    wire new_AGEMA_signal_18087 ;
    wire new_AGEMA_signal_18088 ;
    wire new_AGEMA_signal_18092 ;
    wire new_AGEMA_signal_18093 ;
    wire new_AGEMA_signal_18094 ;
    wire new_AGEMA_signal_18098 ;
    wire new_AGEMA_signal_18099 ;
    wire new_AGEMA_signal_18100 ;
    wire new_AGEMA_signal_18104 ;
    wire new_AGEMA_signal_18105 ;
    wire new_AGEMA_signal_18106 ;
    wire new_AGEMA_signal_18110 ;
    wire new_AGEMA_signal_18111 ;
    wire new_AGEMA_signal_18112 ;
    wire new_AGEMA_signal_18116 ;
    wire new_AGEMA_signal_18117 ;
    wire new_AGEMA_signal_18118 ;
    wire new_AGEMA_signal_18122 ;
    wire new_AGEMA_signal_18123 ;
    wire new_AGEMA_signal_18124 ;
    wire new_AGEMA_signal_18128 ;
    wire new_AGEMA_signal_18129 ;
    wire new_AGEMA_signal_18130 ;
    wire new_AGEMA_signal_18134 ;
    wire new_AGEMA_signal_18135 ;
    wire new_AGEMA_signal_18136 ;
    wire new_AGEMA_signal_18140 ;
    wire new_AGEMA_signal_18141 ;
    wire new_AGEMA_signal_18142 ;
    wire new_AGEMA_signal_18146 ;
    wire new_AGEMA_signal_18147 ;
    wire new_AGEMA_signal_18148 ;
    wire new_AGEMA_signal_18152 ;
    wire new_AGEMA_signal_18153 ;
    wire new_AGEMA_signal_18154 ;
    wire new_AGEMA_signal_18158 ;
    wire new_AGEMA_signal_18159 ;
    wire new_AGEMA_signal_18160 ;
    wire new_AGEMA_signal_18164 ;
    wire new_AGEMA_signal_18165 ;
    wire new_AGEMA_signal_18166 ;
    wire new_AGEMA_signal_18170 ;
    wire new_AGEMA_signal_18171 ;
    wire new_AGEMA_signal_18172 ;
    wire new_AGEMA_signal_18176 ;
    wire new_AGEMA_signal_18177 ;
    wire new_AGEMA_signal_18178 ;
    wire new_AGEMA_signal_18182 ;
    wire new_AGEMA_signal_18183 ;
    wire new_AGEMA_signal_18184 ;
    wire new_AGEMA_signal_18188 ;
    wire new_AGEMA_signal_18189 ;
    wire new_AGEMA_signal_18190 ;
    wire new_AGEMA_signal_18194 ;
    wire new_AGEMA_signal_18195 ;
    wire new_AGEMA_signal_18196 ;
    wire new_AGEMA_signal_18200 ;
    wire new_AGEMA_signal_18201 ;
    wire new_AGEMA_signal_18202 ;
    wire new_AGEMA_signal_18206 ;
    wire new_AGEMA_signal_18207 ;
    wire new_AGEMA_signal_18208 ;
    wire new_AGEMA_signal_18212 ;
    wire new_AGEMA_signal_18213 ;
    wire new_AGEMA_signal_18214 ;
    wire new_AGEMA_signal_18218 ;
    wire new_AGEMA_signal_18219 ;
    wire new_AGEMA_signal_18220 ;
    wire new_AGEMA_signal_18224 ;
    wire new_AGEMA_signal_18225 ;
    wire new_AGEMA_signal_18226 ;
    wire new_AGEMA_signal_18230 ;
    wire new_AGEMA_signal_18231 ;
    wire new_AGEMA_signal_18232 ;
    wire new_AGEMA_signal_18236 ;
    wire new_AGEMA_signal_18237 ;
    wire new_AGEMA_signal_18238 ;
    wire new_AGEMA_signal_18242 ;
    wire new_AGEMA_signal_18243 ;
    wire new_AGEMA_signal_18244 ;
    wire new_AGEMA_signal_18248 ;
    wire new_AGEMA_signal_18249 ;
    wire new_AGEMA_signal_18250 ;
    wire new_AGEMA_signal_18254 ;
    wire new_AGEMA_signal_18255 ;
    wire new_AGEMA_signal_18256 ;
    wire new_AGEMA_signal_18260 ;
    wire new_AGEMA_signal_18261 ;
    wire new_AGEMA_signal_18262 ;
    wire new_AGEMA_signal_18266 ;
    wire new_AGEMA_signal_18267 ;
    wire new_AGEMA_signal_18268 ;
    wire new_AGEMA_signal_18272 ;
    wire new_AGEMA_signal_18273 ;
    wire new_AGEMA_signal_18274 ;
    wire new_AGEMA_signal_18278 ;
    wire new_AGEMA_signal_18279 ;
    wire new_AGEMA_signal_18280 ;
    wire new_AGEMA_signal_18284 ;
    wire new_AGEMA_signal_18285 ;
    wire new_AGEMA_signal_18286 ;
    wire new_AGEMA_signal_18290 ;
    wire new_AGEMA_signal_18291 ;
    wire new_AGEMA_signal_18292 ;
    wire new_AGEMA_signal_18296 ;
    wire new_AGEMA_signal_18297 ;
    wire new_AGEMA_signal_18298 ;
    wire new_AGEMA_signal_18302 ;
    wire new_AGEMA_signal_18303 ;
    wire new_AGEMA_signal_18304 ;
    wire new_AGEMA_signal_18308 ;
    wire new_AGEMA_signal_18309 ;
    wire new_AGEMA_signal_18310 ;
    wire new_AGEMA_signal_18314 ;
    wire new_AGEMA_signal_18315 ;
    wire new_AGEMA_signal_18316 ;
    wire new_AGEMA_signal_18320 ;
    wire new_AGEMA_signal_18321 ;
    wire new_AGEMA_signal_18322 ;
    wire new_AGEMA_signal_18326 ;
    wire new_AGEMA_signal_18327 ;
    wire new_AGEMA_signal_18328 ;
    wire new_AGEMA_signal_18332 ;
    wire new_AGEMA_signal_18333 ;
    wire new_AGEMA_signal_18334 ;
    wire new_AGEMA_signal_18338 ;
    wire new_AGEMA_signal_18339 ;
    wire new_AGEMA_signal_18340 ;
    wire new_AGEMA_signal_18344 ;
    wire new_AGEMA_signal_18345 ;
    wire new_AGEMA_signal_18346 ;
    wire new_AGEMA_signal_18350 ;
    wire new_AGEMA_signal_18351 ;
    wire new_AGEMA_signal_18352 ;
    wire new_AGEMA_signal_18356 ;
    wire new_AGEMA_signal_18357 ;
    wire new_AGEMA_signal_18358 ;
    wire new_AGEMA_signal_18362 ;
    wire new_AGEMA_signal_18363 ;
    wire new_AGEMA_signal_18364 ;
    wire new_AGEMA_signal_18368 ;
    wire new_AGEMA_signal_18369 ;
    wire new_AGEMA_signal_18370 ;
    wire new_AGEMA_signal_18374 ;
    wire new_AGEMA_signal_18375 ;
    wire new_AGEMA_signal_18376 ;
    wire new_AGEMA_signal_18380 ;
    wire new_AGEMA_signal_18381 ;
    wire new_AGEMA_signal_18382 ;
    wire new_AGEMA_signal_18383 ;
    wire new_AGEMA_signal_18384 ;
    wire new_AGEMA_signal_18385 ;
    wire new_AGEMA_signal_18386 ;
    wire new_AGEMA_signal_18387 ;
    wire new_AGEMA_signal_18388 ;
    wire new_AGEMA_signal_18389 ;
    wire new_AGEMA_signal_18390 ;
    wire new_AGEMA_signal_18391 ;
    wire new_AGEMA_signal_18392 ;
    wire new_AGEMA_signal_18393 ;
    wire new_AGEMA_signal_18394 ;
    wire new_AGEMA_signal_18395 ;
    wire new_AGEMA_signal_18396 ;
    wire new_AGEMA_signal_18397 ;
    wire new_AGEMA_signal_18398 ;
    wire new_AGEMA_signal_18399 ;
    wire new_AGEMA_signal_18400 ;
    wire new_AGEMA_signal_18401 ;
    wire new_AGEMA_signal_18402 ;
    wire new_AGEMA_signal_18403 ;
    wire new_AGEMA_signal_18404 ;
    wire new_AGEMA_signal_18405 ;
    wire new_AGEMA_signal_18406 ;
    wire new_AGEMA_signal_18410 ;
    wire new_AGEMA_signal_18411 ;
    wire new_AGEMA_signal_18412 ;
    wire new_AGEMA_signal_18413 ;
    wire new_AGEMA_signal_18414 ;
    wire new_AGEMA_signal_18415 ;
    wire new_AGEMA_signal_18419 ;
    wire new_AGEMA_signal_18420 ;
    wire new_AGEMA_signal_18421 ;
    wire new_AGEMA_signal_18425 ;
    wire new_AGEMA_signal_18426 ;
    wire new_AGEMA_signal_18427 ;
    wire new_AGEMA_signal_18428 ;
    wire new_AGEMA_signal_18429 ;
    wire new_AGEMA_signal_18430 ;
    wire new_AGEMA_signal_18431 ;
    wire new_AGEMA_signal_18432 ;
    wire new_AGEMA_signal_18433 ;
    wire new_AGEMA_signal_18434 ;
    wire new_AGEMA_signal_18435 ;
    wire new_AGEMA_signal_18436 ;
    wire new_AGEMA_signal_18437 ;
    wire new_AGEMA_signal_18438 ;
    wire new_AGEMA_signal_18439 ;
    wire new_AGEMA_signal_18443 ;
    wire new_AGEMA_signal_18444 ;
    wire new_AGEMA_signal_18445 ;
    wire new_AGEMA_signal_18446 ;
    wire new_AGEMA_signal_18447 ;
    wire new_AGEMA_signal_18448 ;
    wire new_AGEMA_signal_18452 ;
    wire new_AGEMA_signal_18453 ;
    wire new_AGEMA_signal_18454 ;
    wire new_AGEMA_signal_18458 ;
    wire new_AGEMA_signal_18459 ;
    wire new_AGEMA_signal_18460 ;
    wire new_AGEMA_signal_18461 ;
    wire new_AGEMA_signal_18462 ;
    wire new_AGEMA_signal_18463 ;
    wire new_AGEMA_signal_18464 ;
    wire new_AGEMA_signal_18465 ;
    wire new_AGEMA_signal_18466 ;
    wire new_AGEMA_signal_18467 ;
    wire new_AGEMA_signal_18468 ;
    wire new_AGEMA_signal_18469 ;
    wire new_AGEMA_signal_18470 ;
    wire new_AGEMA_signal_18471 ;
    wire new_AGEMA_signal_18472 ;
    wire new_AGEMA_signal_18476 ;
    wire new_AGEMA_signal_18477 ;
    wire new_AGEMA_signal_18478 ;
    wire new_AGEMA_signal_18479 ;
    wire new_AGEMA_signal_18480 ;
    wire new_AGEMA_signal_18481 ;
    wire new_AGEMA_signal_18485 ;
    wire new_AGEMA_signal_18486 ;
    wire new_AGEMA_signal_18487 ;
    wire new_AGEMA_signal_18491 ;
    wire new_AGEMA_signal_18492 ;
    wire new_AGEMA_signal_18493 ;
    wire new_AGEMA_signal_18494 ;
    wire new_AGEMA_signal_18495 ;
    wire new_AGEMA_signal_18496 ;
    wire new_AGEMA_signal_18497 ;
    wire new_AGEMA_signal_18498 ;
    wire new_AGEMA_signal_18499 ;
    wire new_AGEMA_signal_18500 ;
    wire new_AGEMA_signal_18501 ;
    wire new_AGEMA_signal_18502 ;
    wire new_AGEMA_signal_18503 ;
    wire new_AGEMA_signal_18504 ;
    wire new_AGEMA_signal_18505 ;
    wire new_AGEMA_signal_18509 ;
    wire new_AGEMA_signal_18510 ;
    wire new_AGEMA_signal_18511 ;
    wire new_AGEMA_signal_18512 ;
    wire new_AGEMA_signal_18513 ;
    wire new_AGEMA_signal_18514 ;
    wire new_AGEMA_signal_18518 ;
    wire new_AGEMA_signal_18519 ;
    wire new_AGEMA_signal_18520 ;
    wire new_AGEMA_signal_18524 ;
    wire new_AGEMA_signal_18525 ;
    wire new_AGEMA_signal_18526 ;
    wire new_AGEMA_signal_18527 ;
    wire new_AGEMA_signal_18528 ;
    wire new_AGEMA_signal_18529 ;
    wire new_AGEMA_signal_18530 ;
    wire new_AGEMA_signal_18531 ;
    wire new_AGEMA_signal_18532 ;
    wire new_AGEMA_signal_18533 ;
    wire new_AGEMA_signal_18534 ;
    wire new_AGEMA_signal_18535 ;
    wire new_AGEMA_signal_18536 ;
    wire new_AGEMA_signal_18537 ;
    wire new_AGEMA_signal_18538 ;
    wire new_AGEMA_signal_18542 ;
    wire new_AGEMA_signal_18543 ;
    wire new_AGEMA_signal_18544 ;
    wire new_AGEMA_signal_18545 ;
    wire new_AGEMA_signal_18546 ;
    wire new_AGEMA_signal_18547 ;
    wire new_AGEMA_signal_18551 ;
    wire new_AGEMA_signal_18552 ;
    wire new_AGEMA_signal_18553 ;
    wire new_AGEMA_signal_18557 ;
    wire new_AGEMA_signal_18558 ;
    wire new_AGEMA_signal_18559 ;
    wire new_AGEMA_signal_18560 ;
    wire new_AGEMA_signal_18561 ;
    wire new_AGEMA_signal_18562 ;
    wire new_AGEMA_signal_18563 ;
    wire new_AGEMA_signal_18564 ;
    wire new_AGEMA_signal_18565 ;
    wire new_AGEMA_signal_18566 ;
    wire new_AGEMA_signal_18567 ;
    wire new_AGEMA_signal_18568 ;
    wire new_AGEMA_signal_18569 ;
    wire new_AGEMA_signal_18570 ;
    wire new_AGEMA_signal_18571 ;
    wire new_AGEMA_signal_18575 ;
    wire new_AGEMA_signal_18576 ;
    wire new_AGEMA_signal_18577 ;
    wire new_AGEMA_signal_18578 ;
    wire new_AGEMA_signal_18579 ;
    wire new_AGEMA_signal_18580 ;
    wire new_AGEMA_signal_18584 ;
    wire new_AGEMA_signal_18585 ;
    wire new_AGEMA_signal_18586 ;
    wire new_AGEMA_signal_18590 ;
    wire new_AGEMA_signal_18591 ;
    wire new_AGEMA_signal_18592 ;
    wire new_AGEMA_signal_18593 ;
    wire new_AGEMA_signal_18594 ;
    wire new_AGEMA_signal_18595 ;
    wire new_AGEMA_signal_18596 ;
    wire new_AGEMA_signal_18597 ;
    wire new_AGEMA_signal_18598 ;
    wire new_AGEMA_signal_18599 ;
    wire new_AGEMA_signal_18600 ;
    wire new_AGEMA_signal_18601 ;
    wire new_AGEMA_signal_18602 ;
    wire new_AGEMA_signal_18603 ;
    wire new_AGEMA_signal_18604 ;
    wire new_AGEMA_signal_18608 ;
    wire new_AGEMA_signal_18609 ;
    wire new_AGEMA_signal_18610 ;
    wire new_AGEMA_signal_18611 ;
    wire new_AGEMA_signal_18612 ;
    wire new_AGEMA_signal_18613 ;
    wire new_AGEMA_signal_18617 ;
    wire new_AGEMA_signal_18618 ;
    wire new_AGEMA_signal_18619 ;
    wire new_AGEMA_signal_18623 ;
    wire new_AGEMA_signal_18624 ;
    wire new_AGEMA_signal_18625 ;
    wire new_AGEMA_signal_18626 ;
    wire new_AGEMA_signal_18627 ;
    wire new_AGEMA_signal_18628 ;
    wire new_AGEMA_signal_18629 ;
    wire new_AGEMA_signal_18630 ;
    wire new_AGEMA_signal_18631 ;
    wire new_AGEMA_signal_18632 ;
    wire new_AGEMA_signal_18633 ;
    wire new_AGEMA_signal_18634 ;
    wire new_AGEMA_signal_18635 ;
    wire new_AGEMA_signal_18636 ;
    wire new_AGEMA_signal_18637 ;
    wire new_AGEMA_signal_18641 ;
    wire new_AGEMA_signal_18642 ;
    wire new_AGEMA_signal_18643 ;
    wire new_AGEMA_signal_18644 ;
    wire new_AGEMA_signal_18645 ;
    wire new_AGEMA_signal_18646 ;
    wire new_AGEMA_signal_18650 ;
    wire new_AGEMA_signal_18651 ;
    wire new_AGEMA_signal_18652 ;
    wire new_AGEMA_signal_18656 ;
    wire new_AGEMA_signal_18657 ;
    wire new_AGEMA_signal_18658 ;
    wire new_AGEMA_signal_18659 ;
    wire new_AGEMA_signal_18660 ;
    wire new_AGEMA_signal_18661 ;
    wire new_AGEMA_signal_18662 ;
    wire new_AGEMA_signal_18663 ;
    wire new_AGEMA_signal_18664 ;
    wire new_AGEMA_signal_18665 ;
    wire new_AGEMA_signal_18666 ;
    wire new_AGEMA_signal_18667 ;
    wire new_AGEMA_signal_18668 ;
    wire new_AGEMA_signal_18669 ;
    wire new_AGEMA_signal_18670 ;
    wire new_AGEMA_signal_18674 ;
    wire new_AGEMA_signal_18675 ;
    wire new_AGEMA_signal_18676 ;
    wire new_AGEMA_signal_18677 ;
    wire new_AGEMA_signal_18678 ;
    wire new_AGEMA_signal_18679 ;
    wire new_AGEMA_signal_18683 ;
    wire new_AGEMA_signal_18684 ;
    wire new_AGEMA_signal_18685 ;
    wire new_AGEMA_signal_18689 ;
    wire new_AGEMA_signal_18690 ;
    wire new_AGEMA_signal_18691 ;
    wire new_AGEMA_signal_18692 ;
    wire new_AGEMA_signal_18693 ;
    wire new_AGEMA_signal_18694 ;
    wire new_AGEMA_signal_18695 ;
    wire new_AGEMA_signal_18696 ;
    wire new_AGEMA_signal_18697 ;
    wire new_AGEMA_signal_18698 ;
    wire new_AGEMA_signal_18699 ;
    wire new_AGEMA_signal_18700 ;
    wire new_AGEMA_signal_18701 ;
    wire new_AGEMA_signal_18702 ;
    wire new_AGEMA_signal_18703 ;
    wire new_AGEMA_signal_18707 ;
    wire new_AGEMA_signal_18708 ;
    wire new_AGEMA_signal_18709 ;
    wire new_AGEMA_signal_18710 ;
    wire new_AGEMA_signal_18711 ;
    wire new_AGEMA_signal_18712 ;
    wire new_AGEMA_signal_18716 ;
    wire new_AGEMA_signal_18717 ;
    wire new_AGEMA_signal_18718 ;
    wire new_AGEMA_signal_18722 ;
    wire new_AGEMA_signal_18723 ;
    wire new_AGEMA_signal_18724 ;
    wire new_AGEMA_signal_18725 ;
    wire new_AGEMA_signal_18726 ;
    wire new_AGEMA_signal_18727 ;
    wire new_AGEMA_signal_18728 ;
    wire new_AGEMA_signal_18729 ;
    wire new_AGEMA_signal_18730 ;
    wire new_AGEMA_signal_18731 ;
    wire new_AGEMA_signal_18732 ;
    wire new_AGEMA_signal_18733 ;
    wire new_AGEMA_signal_18734 ;
    wire new_AGEMA_signal_18735 ;
    wire new_AGEMA_signal_18736 ;
    wire new_AGEMA_signal_18740 ;
    wire new_AGEMA_signal_18741 ;
    wire new_AGEMA_signal_18742 ;
    wire new_AGEMA_signal_18743 ;
    wire new_AGEMA_signal_18744 ;
    wire new_AGEMA_signal_18745 ;
    wire new_AGEMA_signal_18749 ;
    wire new_AGEMA_signal_18750 ;
    wire new_AGEMA_signal_18751 ;
    wire new_AGEMA_signal_18755 ;
    wire new_AGEMA_signal_18756 ;
    wire new_AGEMA_signal_18757 ;
    wire new_AGEMA_signal_18758 ;
    wire new_AGEMA_signal_18759 ;
    wire new_AGEMA_signal_18760 ;
    wire new_AGEMA_signal_18761 ;
    wire new_AGEMA_signal_18762 ;
    wire new_AGEMA_signal_18763 ;
    wire new_AGEMA_signal_18764 ;
    wire new_AGEMA_signal_18765 ;
    wire new_AGEMA_signal_18766 ;
    wire new_AGEMA_signal_18767 ;
    wire new_AGEMA_signal_18768 ;
    wire new_AGEMA_signal_18769 ;
    wire new_AGEMA_signal_18773 ;
    wire new_AGEMA_signal_18774 ;
    wire new_AGEMA_signal_18775 ;
    wire new_AGEMA_signal_18776 ;
    wire new_AGEMA_signal_18777 ;
    wire new_AGEMA_signal_18778 ;
    wire new_AGEMA_signal_18782 ;
    wire new_AGEMA_signal_18783 ;
    wire new_AGEMA_signal_18784 ;
    wire new_AGEMA_signal_18788 ;
    wire new_AGEMA_signal_18789 ;
    wire new_AGEMA_signal_18790 ;
    wire new_AGEMA_signal_18791 ;
    wire new_AGEMA_signal_18792 ;
    wire new_AGEMA_signal_18793 ;
    wire new_AGEMA_signal_18794 ;
    wire new_AGEMA_signal_18795 ;
    wire new_AGEMA_signal_18796 ;
    wire new_AGEMA_signal_18797 ;
    wire new_AGEMA_signal_18798 ;
    wire new_AGEMA_signal_18799 ;
    wire new_AGEMA_signal_18800 ;
    wire new_AGEMA_signal_18801 ;
    wire new_AGEMA_signal_18802 ;
    wire new_AGEMA_signal_18806 ;
    wire new_AGEMA_signal_18807 ;
    wire new_AGEMA_signal_18808 ;
    wire new_AGEMA_signal_18809 ;
    wire new_AGEMA_signal_18810 ;
    wire new_AGEMA_signal_18811 ;
    wire new_AGEMA_signal_18815 ;
    wire new_AGEMA_signal_18816 ;
    wire new_AGEMA_signal_18817 ;
    wire new_AGEMA_signal_18821 ;
    wire new_AGEMA_signal_18822 ;
    wire new_AGEMA_signal_18823 ;
    wire new_AGEMA_signal_18824 ;
    wire new_AGEMA_signal_18825 ;
    wire new_AGEMA_signal_18826 ;
    wire new_AGEMA_signal_18827 ;
    wire new_AGEMA_signal_18828 ;
    wire new_AGEMA_signal_18829 ;
    wire new_AGEMA_signal_18830 ;
    wire new_AGEMA_signal_18831 ;
    wire new_AGEMA_signal_18832 ;
    wire new_AGEMA_signal_18833 ;
    wire new_AGEMA_signal_18834 ;
    wire new_AGEMA_signal_18835 ;
    wire new_AGEMA_signal_18839 ;
    wire new_AGEMA_signal_18840 ;
    wire new_AGEMA_signal_18841 ;
    wire new_AGEMA_signal_18842 ;
    wire new_AGEMA_signal_18843 ;
    wire new_AGEMA_signal_18844 ;
    wire new_AGEMA_signal_18848 ;
    wire new_AGEMA_signal_18849 ;
    wire new_AGEMA_signal_18850 ;
    wire new_AGEMA_signal_18854 ;
    wire new_AGEMA_signal_18855 ;
    wire new_AGEMA_signal_18856 ;
    wire new_AGEMA_signal_18857 ;
    wire new_AGEMA_signal_18858 ;
    wire new_AGEMA_signal_18859 ;
    wire new_AGEMA_signal_18860 ;
    wire new_AGEMA_signal_18861 ;
    wire new_AGEMA_signal_18862 ;
    wire new_AGEMA_signal_18863 ;
    wire new_AGEMA_signal_18864 ;
    wire new_AGEMA_signal_18865 ;
    wire new_AGEMA_signal_18866 ;
    wire new_AGEMA_signal_18867 ;
    wire new_AGEMA_signal_18868 ;
    wire new_AGEMA_signal_18872 ;
    wire new_AGEMA_signal_18873 ;
    wire new_AGEMA_signal_18874 ;
    wire new_AGEMA_signal_18875 ;
    wire new_AGEMA_signal_18876 ;
    wire new_AGEMA_signal_18877 ;
    wire new_AGEMA_signal_18881 ;
    wire new_AGEMA_signal_18882 ;
    wire new_AGEMA_signal_18883 ;
    wire new_AGEMA_signal_18887 ;
    wire new_AGEMA_signal_18888 ;
    wire new_AGEMA_signal_18889 ;
    wire new_AGEMA_signal_18890 ;
    wire new_AGEMA_signal_18891 ;
    wire new_AGEMA_signal_18892 ;
    wire new_AGEMA_signal_18893 ;
    wire new_AGEMA_signal_18894 ;
    wire new_AGEMA_signal_18895 ;
    wire new_AGEMA_signal_18896 ;
    wire new_AGEMA_signal_18897 ;
    wire new_AGEMA_signal_18898 ;
    wire new_AGEMA_signal_18899 ;
    wire new_AGEMA_signal_18900 ;
    wire new_AGEMA_signal_18901 ;
    wire new_AGEMA_signal_18905 ;
    wire new_AGEMA_signal_18906 ;
    wire new_AGEMA_signal_18907 ;
    wire new_AGEMA_signal_18908 ;
    wire new_AGEMA_signal_18909 ;
    wire new_AGEMA_signal_18910 ;
    wire new_AGEMA_signal_18914 ;
    wire new_AGEMA_signal_18915 ;
    wire new_AGEMA_signal_18916 ;
    wire new_AGEMA_signal_18920 ;
    wire new_AGEMA_signal_18921 ;
    wire new_AGEMA_signal_18922 ;
    wire new_AGEMA_signal_18923 ;
    wire new_AGEMA_signal_18924 ;
    wire new_AGEMA_signal_18925 ;
    wire new_AGEMA_signal_18926 ;
    wire new_AGEMA_signal_18927 ;
    wire new_AGEMA_signal_18928 ;
    wire new_AGEMA_signal_18929 ;
    wire new_AGEMA_signal_18930 ;
    wire new_AGEMA_signal_18931 ;
    wire new_AGEMA_signal_18932 ;
    wire new_AGEMA_signal_18933 ;
    wire new_AGEMA_signal_18934 ;
    wire new_AGEMA_signal_18935 ;
    wire new_AGEMA_signal_18936 ;
    wire new_AGEMA_signal_18937 ;
    wire new_AGEMA_signal_18938 ;
    wire new_AGEMA_signal_18939 ;
    wire new_AGEMA_signal_18940 ;
    wire new_AGEMA_signal_18941 ;
    wire new_AGEMA_signal_18942 ;
    wire new_AGEMA_signal_18943 ;
    wire new_AGEMA_signal_18944 ;
    wire new_AGEMA_signal_18945 ;
    wire new_AGEMA_signal_18946 ;
    wire new_AGEMA_signal_18947 ;
    wire new_AGEMA_signal_18948 ;
    wire new_AGEMA_signal_18949 ;
    wire new_AGEMA_signal_18950 ;
    wire new_AGEMA_signal_18951 ;
    wire new_AGEMA_signal_18952 ;
    wire new_AGEMA_signal_18953 ;
    wire new_AGEMA_signal_18954 ;
    wire new_AGEMA_signal_18955 ;
    wire new_AGEMA_signal_18956 ;
    wire new_AGEMA_signal_18957 ;
    wire new_AGEMA_signal_18958 ;
    wire new_AGEMA_signal_18959 ;
    wire new_AGEMA_signal_18960 ;
    wire new_AGEMA_signal_18961 ;
    wire new_AGEMA_signal_18962 ;
    wire new_AGEMA_signal_18963 ;
    wire new_AGEMA_signal_18964 ;
    wire new_AGEMA_signal_18965 ;
    wire new_AGEMA_signal_18966 ;
    wire new_AGEMA_signal_18967 ;
    wire new_AGEMA_signal_18968 ;
    wire new_AGEMA_signal_18969 ;
    wire new_AGEMA_signal_18970 ;
    wire new_AGEMA_signal_18971 ;
    wire new_AGEMA_signal_18972 ;
    wire new_AGEMA_signal_18973 ;
    wire new_AGEMA_signal_18974 ;
    wire new_AGEMA_signal_18975 ;
    wire new_AGEMA_signal_18976 ;
    wire new_AGEMA_signal_18977 ;
    wire new_AGEMA_signal_18978 ;
    wire new_AGEMA_signal_18979 ;
    wire new_AGEMA_signal_18980 ;
    wire new_AGEMA_signal_18981 ;
    wire new_AGEMA_signal_18982 ;
    wire new_AGEMA_signal_18983 ;
    wire new_AGEMA_signal_18984 ;
    wire new_AGEMA_signal_18985 ;
    wire new_AGEMA_signal_18986 ;
    wire new_AGEMA_signal_18987 ;
    wire new_AGEMA_signal_18988 ;
    wire new_AGEMA_signal_18989 ;
    wire new_AGEMA_signal_18990 ;
    wire new_AGEMA_signal_18991 ;
    wire new_AGEMA_signal_18992 ;
    wire new_AGEMA_signal_18993 ;
    wire new_AGEMA_signal_18994 ;
    wire new_AGEMA_signal_18995 ;
    wire new_AGEMA_signal_18996 ;
    wire new_AGEMA_signal_18997 ;
    wire new_AGEMA_signal_18998 ;
    wire new_AGEMA_signal_18999 ;
    wire new_AGEMA_signal_19000 ;
    wire new_AGEMA_signal_19001 ;
    wire new_AGEMA_signal_19002 ;
    wire new_AGEMA_signal_19003 ;
    wire new_AGEMA_signal_19004 ;
    wire new_AGEMA_signal_19005 ;
    wire new_AGEMA_signal_19006 ;
    wire new_AGEMA_signal_19007 ;
    wire new_AGEMA_signal_19008 ;
    wire new_AGEMA_signal_19009 ;
    wire new_AGEMA_signal_19010 ;
    wire new_AGEMA_signal_19011 ;
    wire new_AGEMA_signal_19012 ;
    wire new_AGEMA_signal_19013 ;
    wire new_AGEMA_signal_19014 ;
    wire new_AGEMA_signal_19015 ;
    wire new_AGEMA_signal_19016 ;
    wire new_AGEMA_signal_19017 ;
    wire new_AGEMA_signal_19018 ;
    wire new_AGEMA_signal_19019 ;
    wire new_AGEMA_signal_19020 ;
    wire new_AGEMA_signal_19021 ;
    wire new_AGEMA_signal_19022 ;
    wire new_AGEMA_signal_19023 ;
    wire new_AGEMA_signal_19024 ;
    wire new_AGEMA_signal_19025 ;
    wire new_AGEMA_signal_19026 ;
    wire new_AGEMA_signal_19027 ;
    wire new_AGEMA_signal_19028 ;
    wire new_AGEMA_signal_19029 ;
    wire new_AGEMA_signal_19030 ;
    wire new_AGEMA_signal_19031 ;
    wire new_AGEMA_signal_19032 ;
    wire new_AGEMA_signal_19033 ;
    wire new_AGEMA_signal_19034 ;
    wire new_AGEMA_signal_19035 ;
    wire new_AGEMA_signal_19036 ;
    wire new_AGEMA_signal_19037 ;
    wire new_AGEMA_signal_19038 ;
    wire new_AGEMA_signal_19039 ;
    wire new_AGEMA_signal_19040 ;
    wire new_AGEMA_signal_19041 ;
    wire new_AGEMA_signal_19042 ;
    wire new_AGEMA_signal_19043 ;
    wire new_AGEMA_signal_19044 ;
    wire new_AGEMA_signal_19045 ;
    wire new_AGEMA_signal_19046 ;
    wire new_AGEMA_signal_19047 ;
    wire new_AGEMA_signal_19048 ;
    wire new_AGEMA_signal_19049 ;
    wire new_AGEMA_signal_19050 ;
    wire new_AGEMA_signal_19051 ;
    wire new_AGEMA_signal_19052 ;
    wire new_AGEMA_signal_19053 ;
    wire new_AGEMA_signal_19054 ;
    wire new_AGEMA_signal_19055 ;
    wire new_AGEMA_signal_19056 ;
    wire new_AGEMA_signal_19057 ;
    wire new_AGEMA_signal_19058 ;
    wire new_AGEMA_signal_19059 ;
    wire new_AGEMA_signal_19060 ;
    wire new_AGEMA_signal_19061 ;
    wire new_AGEMA_signal_19062 ;
    wire new_AGEMA_signal_19063 ;
    wire new_AGEMA_signal_19064 ;
    wire new_AGEMA_signal_19065 ;
    wire new_AGEMA_signal_19066 ;
    wire new_AGEMA_signal_19067 ;
    wire new_AGEMA_signal_19068 ;
    wire new_AGEMA_signal_19069 ;
    wire new_AGEMA_signal_19070 ;
    wire new_AGEMA_signal_19071 ;
    wire new_AGEMA_signal_19072 ;
    wire new_AGEMA_signal_19073 ;
    wire new_AGEMA_signal_19074 ;
    wire new_AGEMA_signal_19075 ;

    /* cells in depth 0 */
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1093 ( .A0_t (RoundCounter[0]), .A0_f (new_AGEMA_signal_5054), .B0_t (n592), .B0_f (new_AGEMA_signal_6336), .Z0_t (n577), .Z0_f (new_AGEMA_signal_6924) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1099 ( .A0_t (RoundCounter[3]), .A0_f (new_AGEMA_signal_5055), .B0_t (n585), .B0_f (new_AGEMA_signal_5053), .Z0_t (n592), .Z0_f (new_AGEMA_signal_6336) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1100 ( .A0_t (RoundCounter[1]), .A0_f (new_AGEMA_signal_5051), .B0_t (RoundCounter[2]), .B0_f (new_AGEMA_signal_5052), .Z0_t (n585), .Z0_f (new_AGEMA_signal_5053) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1103 ( .A0_t (RoundCounter[0]), .A0_f (new_AGEMA_signal_5054), .B0_t (n585), .B0_f (new_AGEMA_signal_5053), .Z0_t (Rcon[0]), .Z0_f (new_AGEMA_signal_6337) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1104 ( .A0_t (RoundCounter[0]), .A0_f (new_AGEMA_signal_5054), .B0_t (RoundCounter[3]), .B0_f (new_AGEMA_signal_5055), .Z0_t (n855), .Z0_f (new_AGEMA_signal_5056) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1105 ( .A0_t (n855), .A0_f (new_AGEMA_signal_5056), .B0_t (n585), .B0_f (new_AGEMA_signal_5053), .Z0_t (Rcon[1]), .Z0_f (new_AGEMA_signal_6338) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1107 ( .A0_t (RoundCounter[2]), .A0_f (new_AGEMA_signal_5052), .B0_t (RoundCounter[1]), .B0_f (new_AGEMA_signal_5051), .Z0_t (n851), .Z0_f (new_AGEMA_signal_5057) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1108 ( .A0_t (n855), .A0_f (new_AGEMA_signal_5056), .B0_t (n851), .B0_f (new_AGEMA_signal_5057), .Z0_t (n586), .Z0_f (new_AGEMA_signal_6339) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1109 ( .A0_t (n577), .A0_f (new_AGEMA_signal_6924), .B0_t (n586), .B0_f (new_AGEMA_signal_6339), .Z0_t (Rcon[2]), .Z0_f (new_AGEMA_signal_7469) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1110 ( .A0_t (RoundCounter[3]), .A0_f (new_AGEMA_signal_5055), .B0_t (RoundCounter[0]), .B0_f (new_AGEMA_signal_5054), .Z0_t (n853), .Z0_f (new_AGEMA_signal_5058) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1111 ( .A0_t (n851), .A0_f (new_AGEMA_signal_5057), .B0_t (n853), .B0_f (new_AGEMA_signal_5058), .Z0_t (n589), .Z0_f (new_AGEMA_signal_6340) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1112 ( .A0_t (RoundCounter[3]), .A0_f (new_AGEMA_signal_5055), .B0_t (Rcon[0]), .B0_f (new_AGEMA_signal_6337), .Z0_t (n588), .Z0_f (new_AGEMA_signal_6925) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1113 ( .A0_t (n589), .A0_f (new_AGEMA_signal_6340), .B0_t (n588), .B0_f (new_AGEMA_signal_6925), .Z0_t (Rcon[3]), .Z0_f (new_AGEMA_signal_7470) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1114 ( .A0_t (RoundCounter[1]), .A0_f (new_AGEMA_signal_5051), .B0_t (RoundCounter[2]), .B0_f (new_AGEMA_signal_5052), .Z0_t (n593), .Z0_f (new_AGEMA_signal_5059) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1115 ( .A0_t (n855), .A0_f (new_AGEMA_signal_5056), .B0_t (n593), .B0_f (new_AGEMA_signal_5059), .Z0_t (n591), .Z0_f (new_AGEMA_signal_6341) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1116 ( .A0_t (n592), .A0_f (new_AGEMA_signal_6336), .B0_t (n591), .B0_f (new_AGEMA_signal_6341), .Z0_t (Rcon[4]), .Z0_f (new_AGEMA_signal_6926) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1117 ( .A0_t (n853), .A0_f (new_AGEMA_signal_5058), .B0_t (n593), .B0_f (new_AGEMA_signal_5059), .Z0_t (n594), .Z0_f (new_AGEMA_signal_6342) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1118 ( .A0_t (n577), .A0_f (new_AGEMA_signal_6924), .B0_t (n594), .B0_f (new_AGEMA_signal_6342), .Z0_t (Rcon[5]), .Z0_f (new_AGEMA_signal_7471) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1119 ( .A0_t (MixColumnsOutput[0]), .A0_f (new_AGEMA_signal_16193), .A1_t (new_AGEMA_signal_16194), .A1_f (new_AGEMA_signal_16195), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n596), .Z0_f (new_AGEMA_signal_16571), .Z1_t (new_AGEMA_signal_16572), .Z1_f (new_AGEMA_signal_16573) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1120 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[0]), .B0_f (new_AGEMA_signal_13130), .B1_t (new_AGEMA_signal_13131), .B1_f (new_AGEMA_signal_13132), .Z0_t (n595), .Z0_f (new_AGEMA_signal_13592), .Z1_t (new_AGEMA_signal_13593), .Z1_f (new_AGEMA_signal_13594) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1121 ( .A0_t (n596), .A0_f (new_AGEMA_signal_16571), .A1_t (new_AGEMA_signal_16572), .A1_f (new_AGEMA_signal_16573), .B0_t (n595), .B0_f (new_AGEMA_signal_13592), .B1_t (new_AGEMA_signal_13593), .B1_f (new_AGEMA_signal_13594), .Z0_t (RoundOutput[0]), .Z0_f (new_AGEMA_signal_17246), .Z1_t (new_AGEMA_signal_17247), .Z1_f (new_AGEMA_signal_17248) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1122 ( .A0_t (MixColumnsOutput[100]), .A0_f (new_AGEMA_signal_16814), .A1_t (new_AGEMA_signal_16815), .A1_f (new_AGEMA_signal_16816), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n598), .Z0_f (new_AGEMA_signal_17249), .Z1_t (new_AGEMA_signal_17250), .Z1_f (new_AGEMA_signal_17251) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1123 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .B0_f (new_AGEMA_signal_13649), .B1_t (new_AGEMA_signal_13650), .B1_f (new_AGEMA_signal_13651), .Z0_t (n597), .Z0_f (new_AGEMA_signal_14090), .Z1_t (new_AGEMA_signal_14091), .Z1_f (new_AGEMA_signal_14092) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1124 ( .A0_t (n598), .A0_f (new_AGEMA_signal_17249), .A1_t (new_AGEMA_signal_17250), .A1_f (new_AGEMA_signal_17251), .B0_t (n597), .B0_f (new_AGEMA_signal_14090), .B1_t (new_AGEMA_signal_14091), .B1_f (new_AGEMA_signal_14092), .Z0_t (RoundOutput[100]), .Z0_f (new_AGEMA_signal_17759), .Z1_t (new_AGEMA_signal_17760), .Z1_f (new_AGEMA_signal_17761) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1125 ( .A0_t (MixColumnsOutput[101]), .A0_f (new_AGEMA_signal_15824), .A1_t (new_AGEMA_signal_15825), .A1_f (new_AGEMA_signal_15826), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n600), .Z0_f (new_AGEMA_signal_16574), .Z1_t (new_AGEMA_signal_16575), .Z1_f (new_AGEMA_signal_16576) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1126 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .B0_f (new_AGEMA_signal_13646), .B1_t (new_AGEMA_signal_13647), .B1_f (new_AGEMA_signal_13648), .Z0_t (n599), .Z0_f (new_AGEMA_signal_14093), .Z1_t (new_AGEMA_signal_14094), .Z1_f (new_AGEMA_signal_14095) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1127 ( .A0_t (n600), .A0_f (new_AGEMA_signal_16574), .A1_t (new_AGEMA_signal_16575), .A1_f (new_AGEMA_signal_16576), .B0_t (n599), .B0_f (new_AGEMA_signal_14093), .B1_t (new_AGEMA_signal_14094), .B1_f (new_AGEMA_signal_14095), .Z0_t (RoundOutput[101]), .Z0_f (new_AGEMA_signal_17252), .Z1_t (new_AGEMA_signal_17253), .Z1_f (new_AGEMA_signal_17254) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1128 ( .A0_t (MixColumnsOutput[102]), .A0_f (new_AGEMA_signal_15821), .A1_t (new_AGEMA_signal_15822), .A1_f (new_AGEMA_signal_15823), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n602), .Z0_f (new_AGEMA_signal_16577), .Z1_t (new_AGEMA_signal_16578), .Z1_f (new_AGEMA_signal_16579) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1129 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .B0_f (new_AGEMA_signal_13643), .B1_t (new_AGEMA_signal_13644), .B1_f (new_AGEMA_signal_13645), .Z0_t (n601), .Z0_f (new_AGEMA_signal_14096), .Z1_t (new_AGEMA_signal_14097), .Z1_f (new_AGEMA_signal_14098) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1130 ( .A0_t (n602), .A0_f (new_AGEMA_signal_16577), .A1_t (new_AGEMA_signal_16578), .A1_f (new_AGEMA_signal_16579), .B0_t (n601), .B0_f (new_AGEMA_signal_14096), .B1_t (new_AGEMA_signal_14097), .B1_f (new_AGEMA_signal_14098), .Z0_t (RoundOutput[102]), .Z0_f (new_AGEMA_signal_17255), .Z1_t (new_AGEMA_signal_17256), .Z1_f (new_AGEMA_signal_17257) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1131 ( .A0_t (MixColumnsOutput[103]), .A0_f (new_AGEMA_signal_15818), .A1_t (new_AGEMA_signal_15819), .A1_f (new_AGEMA_signal_15820), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n604), .Z0_f (new_AGEMA_signal_16580), .Z1_t (new_AGEMA_signal_16581), .Z1_f (new_AGEMA_signal_16582) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1132 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B0_f (new_AGEMA_signal_13640), .B1_t (new_AGEMA_signal_13641), .B1_f (new_AGEMA_signal_13642), .Z0_t (n603), .Z0_f (new_AGEMA_signal_14099), .Z1_t (new_AGEMA_signal_14100), .Z1_f (new_AGEMA_signal_14101) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1133 ( .A0_t (n604), .A0_f (new_AGEMA_signal_16580), .A1_t (new_AGEMA_signal_16581), .A1_f (new_AGEMA_signal_16582), .B0_t (n603), .B0_f (new_AGEMA_signal_14099), .B1_t (new_AGEMA_signal_14100), .B1_f (new_AGEMA_signal_14101), .Z0_t (RoundOutput[103]), .Z0_f (new_AGEMA_signal_17258), .Z1_t (new_AGEMA_signal_17259), .Z1_f (new_AGEMA_signal_17260) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1134 ( .A0_t (MixColumnsOutput[104]), .A0_f (new_AGEMA_signal_15815), .A1_t (new_AGEMA_signal_15816), .A1_f (new_AGEMA_signal_15817), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n606), .Z0_f (new_AGEMA_signal_16583), .Z1_t (new_AGEMA_signal_16584), .Z1_f (new_AGEMA_signal_16585) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1135 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[104]), .B0_f (new_AGEMA_signal_13163), .B1_t (new_AGEMA_signal_13164), .B1_f (new_AGEMA_signal_13165), .Z0_t (n605), .Z0_f (new_AGEMA_signal_13595), .Z1_t (new_AGEMA_signal_13596), .Z1_f (new_AGEMA_signal_13597) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1136 ( .A0_t (n606), .A0_f (new_AGEMA_signal_16583), .A1_t (new_AGEMA_signal_16584), .A1_f (new_AGEMA_signal_16585), .B0_t (n605), .B0_f (new_AGEMA_signal_13595), .B1_t (new_AGEMA_signal_13596), .B1_f (new_AGEMA_signal_13597), .Z0_t (RoundOutput[104]), .Z0_f (new_AGEMA_signal_17261), .Z1_t (new_AGEMA_signal_17262), .Z1_f (new_AGEMA_signal_17263) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1137 ( .A0_t (MixColumnsOutput[105]), .A0_f (new_AGEMA_signal_16811), .A1_t (new_AGEMA_signal_16812), .A1_f (new_AGEMA_signal_16813), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n608), .Z0_f (new_AGEMA_signal_17264), .Z1_t (new_AGEMA_signal_17265), .Z1_f (new_AGEMA_signal_17266) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1138 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13763), .B1_t (new_AGEMA_signal_13764), .B1_f (new_AGEMA_signal_13765), .Z0_t (n607), .Z0_f (new_AGEMA_signal_14102), .Z1_t (new_AGEMA_signal_14103), .Z1_f (new_AGEMA_signal_14104) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1139 ( .A0_t (n608), .A0_f (new_AGEMA_signal_17264), .A1_t (new_AGEMA_signal_17265), .A1_f (new_AGEMA_signal_17266), .B0_t (n607), .B0_f (new_AGEMA_signal_14102), .B1_t (new_AGEMA_signal_14103), .B1_f (new_AGEMA_signal_14104), .Z0_t (RoundOutput[105]), .Z0_f (new_AGEMA_signal_17762), .Z1_t (new_AGEMA_signal_17763), .Z1_f (new_AGEMA_signal_17764) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1140 ( .A0_t (MixColumnsOutput[106]), .A0_f (new_AGEMA_signal_15902), .A1_t (new_AGEMA_signal_15903), .A1_f (new_AGEMA_signal_15904), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n610), .Z0_f (new_AGEMA_signal_16586), .Z1_t (new_AGEMA_signal_16587), .Z1_f (new_AGEMA_signal_16588) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1141 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[106]), .B0_f (new_AGEMA_signal_13760), .B1_t (new_AGEMA_signal_13761), .B1_f (new_AGEMA_signal_13762), .Z0_t (n609), .Z0_f (new_AGEMA_signal_14105), .Z1_t (new_AGEMA_signal_14106), .Z1_f (new_AGEMA_signal_14107) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1142 ( .A0_t (n610), .A0_f (new_AGEMA_signal_16586), .A1_t (new_AGEMA_signal_16587), .A1_f (new_AGEMA_signal_16588), .B0_t (n609), .B0_f (new_AGEMA_signal_14105), .B1_t (new_AGEMA_signal_14106), .B1_f (new_AGEMA_signal_14107), .Z0_t (RoundOutput[106]), .Z0_f (new_AGEMA_signal_17267), .Z1_t (new_AGEMA_signal_17268), .Z1_f (new_AGEMA_signal_17269) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1143 ( .A0_t (MixColumnsOutput[107]), .A0_f (new_AGEMA_signal_16844), .A1_t (new_AGEMA_signal_16845), .A1_f (new_AGEMA_signal_16846), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n612), .Z0_f (new_AGEMA_signal_17270), .Z1_t (new_AGEMA_signal_17271), .Z1_f (new_AGEMA_signal_17272) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1144 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[107]), .B0_f (new_AGEMA_signal_13757), .B1_t (new_AGEMA_signal_13758), .B1_f (new_AGEMA_signal_13759), .Z0_t (n611), .Z0_f (new_AGEMA_signal_14108), .Z1_t (new_AGEMA_signal_14109), .Z1_f (new_AGEMA_signal_14110) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1145 ( .A0_t (n612), .A0_f (new_AGEMA_signal_17270), .A1_t (new_AGEMA_signal_17271), .A1_f (new_AGEMA_signal_17272), .B0_t (n611), .B0_f (new_AGEMA_signal_14108), .B1_t (new_AGEMA_signal_14109), .B1_f (new_AGEMA_signal_14110), .Z0_t (RoundOutput[107]), .Z0_f (new_AGEMA_signal_17765), .Z1_t (new_AGEMA_signal_17766), .Z1_f (new_AGEMA_signal_17767) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1146 ( .A0_t (MixColumnsOutput[108]), .A0_f (new_AGEMA_signal_16841), .A1_t (new_AGEMA_signal_16842), .A1_f (new_AGEMA_signal_16843), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n614), .Z0_f (new_AGEMA_signal_17273), .Z1_t (new_AGEMA_signal_17274), .Z1_f (new_AGEMA_signal_17275) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1147 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13754), .B1_t (new_AGEMA_signal_13755), .B1_f (new_AGEMA_signal_13756), .Z0_t (n613), .Z0_f (new_AGEMA_signal_14111), .Z1_t (new_AGEMA_signal_14112), .Z1_f (new_AGEMA_signal_14113) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1148 ( .A0_t (n614), .A0_f (new_AGEMA_signal_17273), .A1_t (new_AGEMA_signal_17274), .A1_f (new_AGEMA_signal_17275), .B0_t (n613), .B0_f (new_AGEMA_signal_14111), .B1_t (new_AGEMA_signal_14112), .B1_f (new_AGEMA_signal_14113), .Z0_t (RoundOutput[108]), .Z0_f (new_AGEMA_signal_17768), .Z1_t (new_AGEMA_signal_17769), .Z1_f (new_AGEMA_signal_17770) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1149 ( .A0_t (MixColumnsOutput[109]), .A0_f (new_AGEMA_signal_15893), .A1_t (new_AGEMA_signal_15894), .A1_f (new_AGEMA_signal_15895), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n616), .Z0_f (new_AGEMA_signal_16589), .Z1_t (new_AGEMA_signal_16590), .Z1_f (new_AGEMA_signal_16591) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1150 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13751), .B1_t (new_AGEMA_signal_13752), .B1_f (new_AGEMA_signal_13753), .Z0_t (n615), .Z0_f (new_AGEMA_signal_14114), .Z1_t (new_AGEMA_signal_14115), .Z1_f (new_AGEMA_signal_14116) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1151 ( .A0_t (n616), .A0_f (new_AGEMA_signal_16589), .A1_t (new_AGEMA_signal_16590), .A1_f (new_AGEMA_signal_16591), .B0_t (n615), .B0_f (new_AGEMA_signal_14114), .B1_t (new_AGEMA_signal_14115), .B1_f (new_AGEMA_signal_14116), .Z0_t (RoundOutput[109]), .Z0_f (new_AGEMA_signal_17276), .Z1_t (new_AGEMA_signal_17277), .Z1_f (new_AGEMA_signal_17278) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1152 ( .A0_t (MixColumnsOutput[10]), .A0_f (new_AGEMA_signal_16190), .A1_t (new_AGEMA_signal_16191), .A1_f (new_AGEMA_signal_16192), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n618), .Z0_f (new_AGEMA_signal_16592), .Z1_t (new_AGEMA_signal_16593), .Z1_f (new_AGEMA_signal_16594) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1153 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[10]), .B0_f (new_AGEMA_signal_13844), .B1_t (new_AGEMA_signal_13845), .B1_f (new_AGEMA_signal_13846), .Z0_t (n617), .Z0_f (new_AGEMA_signal_14117), .Z1_t (new_AGEMA_signal_14118), .Z1_f (new_AGEMA_signal_14119) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1154 ( .A0_t (n618), .A0_f (new_AGEMA_signal_16592), .A1_t (new_AGEMA_signal_16593), .A1_f (new_AGEMA_signal_16594), .B0_t (n617), .B0_f (new_AGEMA_signal_14117), .B1_t (new_AGEMA_signal_14118), .B1_f (new_AGEMA_signal_14119), .Z0_t (RoundOutput[10]), .Z0_f (new_AGEMA_signal_17279), .Z1_t (new_AGEMA_signal_17280), .Z1_f (new_AGEMA_signal_17281) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1155 ( .A0_t (MixColumnsOutput[110]), .A0_f (new_AGEMA_signal_15890), .A1_t (new_AGEMA_signal_15891), .A1_f (new_AGEMA_signal_15892), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n620), .Z0_f (new_AGEMA_signal_16595), .Z1_t (new_AGEMA_signal_16596), .Z1_f (new_AGEMA_signal_16597) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1156 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13748), .B1_t (new_AGEMA_signal_13749), .B1_f (new_AGEMA_signal_13750), .Z0_t (n619), .Z0_f (new_AGEMA_signal_14120), .Z1_t (new_AGEMA_signal_14121), .Z1_f (new_AGEMA_signal_14122) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1157 ( .A0_t (n620), .A0_f (new_AGEMA_signal_16595), .A1_t (new_AGEMA_signal_16596), .A1_f (new_AGEMA_signal_16597), .B0_t (n619), .B0_f (new_AGEMA_signal_14120), .B1_t (new_AGEMA_signal_14121), .B1_f (new_AGEMA_signal_14122), .Z0_t (RoundOutput[110]), .Z0_f (new_AGEMA_signal_17282), .Z1_t (new_AGEMA_signal_17283), .Z1_f (new_AGEMA_signal_17284) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1158 ( .A0_t (MixColumnsOutput[111]), .A0_f (new_AGEMA_signal_15887), .A1_t (new_AGEMA_signal_15888), .A1_f (new_AGEMA_signal_15889), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n622), .Z0_f (new_AGEMA_signal_16598), .Z1_t (new_AGEMA_signal_16599), .Z1_f (new_AGEMA_signal_16600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1159 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B0_f (new_AGEMA_signal_13745), .B1_t (new_AGEMA_signal_13746), .B1_f (new_AGEMA_signal_13747), .Z0_t (n621), .Z0_f (new_AGEMA_signal_14123), .Z1_t (new_AGEMA_signal_14124), .Z1_f (new_AGEMA_signal_14125) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1160 ( .A0_t (n622), .A0_f (new_AGEMA_signal_16598), .A1_t (new_AGEMA_signal_16599), .A1_f (new_AGEMA_signal_16600), .B0_t (n621), .B0_f (new_AGEMA_signal_14123), .B1_t (new_AGEMA_signal_14124), .B1_f (new_AGEMA_signal_14125), .Z0_t (RoundOutput[111]), .Z0_f (new_AGEMA_signal_17285), .Z1_t (new_AGEMA_signal_17286), .Z1_f (new_AGEMA_signal_17287) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1161 ( .A0_t (MixColumnsOutput[112]), .A0_f (new_AGEMA_signal_15884), .A1_t (new_AGEMA_signal_15885), .A1_f (new_AGEMA_signal_15886), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n624), .Z0_f (new_AGEMA_signal_16601), .Z1_t (new_AGEMA_signal_16602), .Z1_f (new_AGEMA_signal_16603) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1162 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[112]), .B0_f (new_AGEMA_signal_13328), .B1_t (new_AGEMA_signal_13329), .B1_f (new_AGEMA_signal_13330), .Z0_t (n623), .Z0_f (new_AGEMA_signal_13598), .Z1_t (new_AGEMA_signal_13599), .Z1_f (new_AGEMA_signal_13600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1163 ( .A0_t (n624), .A0_f (new_AGEMA_signal_16601), .A1_t (new_AGEMA_signal_16602), .A1_f (new_AGEMA_signal_16603), .B0_t (n623), .B0_f (new_AGEMA_signal_13598), .B1_t (new_AGEMA_signal_13599), .B1_f (new_AGEMA_signal_13600), .Z0_t (RoundOutput[112]), .Z0_f (new_AGEMA_signal_17288), .Z1_t (new_AGEMA_signal_17289), .Z1_f (new_AGEMA_signal_17290) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1164 ( .A0_t (MixColumnsOutput[113]), .A0_f (new_AGEMA_signal_16838), .A1_t (new_AGEMA_signal_16839), .A1_f (new_AGEMA_signal_16840), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n626), .Z0_f (new_AGEMA_signal_17291), .Z1_t (new_AGEMA_signal_17292), .Z1_f (new_AGEMA_signal_17293) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1165 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13868), .B1_t (new_AGEMA_signal_13869), .B1_f (new_AGEMA_signal_13870), .Z0_t (n625), .Z0_f (new_AGEMA_signal_14126), .Z1_t (new_AGEMA_signal_14127), .Z1_f (new_AGEMA_signal_14128) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1166 ( .A0_t (n626), .A0_f (new_AGEMA_signal_17291), .A1_t (new_AGEMA_signal_17292), .A1_f (new_AGEMA_signal_17293), .B0_t (n625), .B0_f (new_AGEMA_signal_14126), .B1_t (new_AGEMA_signal_14127), .B1_f (new_AGEMA_signal_14128), .Z0_t (RoundOutput[113]), .Z0_f (new_AGEMA_signal_17771), .Z1_t (new_AGEMA_signal_17772), .Z1_f (new_AGEMA_signal_17773) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1167 ( .A0_t (MixColumnsOutput[114]), .A0_f (new_AGEMA_signal_15878), .A1_t (new_AGEMA_signal_15879), .A1_f (new_AGEMA_signal_15880), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n628), .Z0_f (new_AGEMA_signal_16604), .Z1_t (new_AGEMA_signal_16605), .Z1_f (new_AGEMA_signal_16606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1168 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[114]), .B0_f (new_AGEMA_signal_13865), .B1_t (new_AGEMA_signal_13866), .B1_f (new_AGEMA_signal_13867), .Z0_t (n627), .Z0_f (new_AGEMA_signal_14129), .Z1_t (new_AGEMA_signal_14130), .Z1_f (new_AGEMA_signal_14131) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1169 ( .A0_t (n628), .A0_f (new_AGEMA_signal_16604), .A1_t (new_AGEMA_signal_16605), .A1_f (new_AGEMA_signal_16606), .B0_t (n627), .B0_f (new_AGEMA_signal_14129), .B1_t (new_AGEMA_signal_14130), .B1_f (new_AGEMA_signal_14131), .Z0_t (RoundOutput[114]), .Z0_f (new_AGEMA_signal_17294), .Z1_t (new_AGEMA_signal_17295), .Z1_f (new_AGEMA_signal_17296) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1170 ( .A0_t (MixColumnsOutput[115]), .A0_f (new_AGEMA_signal_16835), .A1_t (new_AGEMA_signal_16836), .A1_f (new_AGEMA_signal_16837), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n630), .Z0_f (new_AGEMA_signal_17297), .Z1_t (new_AGEMA_signal_17298), .Z1_f (new_AGEMA_signal_17299) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1171 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[115]), .B0_f (new_AGEMA_signal_13862), .B1_t (new_AGEMA_signal_13863), .B1_f (new_AGEMA_signal_13864), .Z0_t (n629), .Z0_f (new_AGEMA_signal_14132), .Z1_t (new_AGEMA_signal_14133), .Z1_f (new_AGEMA_signal_14134) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1172 ( .A0_t (n630), .A0_f (new_AGEMA_signal_17297), .A1_t (new_AGEMA_signal_17298), .A1_f (new_AGEMA_signal_17299), .B0_t (n629), .B0_f (new_AGEMA_signal_14132), .B1_t (new_AGEMA_signal_14133), .B1_f (new_AGEMA_signal_14134), .Z0_t (RoundOutput[115]), .Z0_f (new_AGEMA_signal_17774), .Z1_t (new_AGEMA_signal_17775), .Z1_f (new_AGEMA_signal_17776) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1173 ( .A0_t (MixColumnsOutput[116]), .A0_f (new_AGEMA_signal_16829), .A1_t (new_AGEMA_signal_16830), .A1_f (new_AGEMA_signal_16831), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n632), .Z0_f (new_AGEMA_signal_17300), .Z1_t (new_AGEMA_signal_17301), .Z1_f (new_AGEMA_signal_17302) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1174 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13859), .B1_t (new_AGEMA_signal_13860), .B1_f (new_AGEMA_signal_13861), .Z0_t (n631), .Z0_f (new_AGEMA_signal_14135), .Z1_t (new_AGEMA_signal_14136), .Z1_f (new_AGEMA_signal_14137) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1175 ( .A0_t (n632), .A0_f (new_AGEMA_signal_17300), .A1_t (new_AGEMA_signal_17301), .A1_f (new_AGEMA_signal_17302), .B0_t (n631), .B0_f (new_AGEMA_signal_14135), .B1_t (new_AGEMA_signal_14136), .B1_f (new_AGEMA_signal_14137), .Z0_t (RoundOutput[116]), .Z0_f (new_AGEMA_signal_17777), .Z1_t (new_AGEMA_signal_17778), .Z1_f (new_AGEMA_signal_17779) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1176 ( .A0_t (MixColumnsOutput[117]), .A0_f (new_AGEMA_signal_15866), .A1_t (new_AGEMA_signal_15867), .A1_f (new_AGEMA_signal_15868), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n634), .Z0_f (new_AGEMA_signal_16607), .Z1_t (new_AGEMA_signal_16608), .Z1_f (new_AGEMA_signal_16609) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1177 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13856), .B1_t (new_AGEMA_signal_13857), .B1_f (new_AGEMA_signal_13858), .Z0_t (n633), .Z0_f (new_AGEMA_signal_14138), .Z1_t (new_AGEMA_signal_14139), .Z1_f (new_AGEMA_signal_14140) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1178 ( .A0_t (n634), .A0_f (new_AGEMA_signal_16607), .A1_t (new_AGEMA_signal_16608), .A1_f (new_AGEMA_signal_16609), .B0_t (n633), .B0_f (new_AGEMA_signal_14138), .B1_t (new_AGEMA_signal_14139), .B1_f (new_AGEMA_signal_14140), .Z0_t (RoundOutput[117]), .Z0_f (new_AGEMA_signal_17303), .Z1_t (new_AGEMA_signal_17304), .Z1_f (new_AGEMA_signal_17305) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1179 ( .A0_t (MixColumnsOutput[118]), .A0_f (new_AGEMA_signal_15863), .A1_t (new_AGEMA_signal_15864), .A1_f (new_AGEMA_signal_15865), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n636), .Z0_f (new_AGEMA_signal_16610), .Z1_t (new_AGEMA_signal_16611), .Z1_f (new_AGEMA_signal_16612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1180 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13853), .B1_t (new_AGEMA_signal_13854), .B1_f (new_AGEMA_signal_13855), .Z0_t (n635), .Z0_f (new_AGEMA_signal_14141), .Z1_t (new_AGEMA_signal_14142), .Z1_f (new_AGEMA_signal_14143) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1181 ( .A0_t (n636), .A0_f (new_AGEMA_signal_16610), .A1_t (new_AGEMA_signal_16611), .A1_f (new_AGEMA_signal_16612), .B0_t (n635), .B0_f (new_AGEMA_signal_14141), .B1_t (new_AGEMA_signal_14142), .B1_f (new_AGEMA_signal_14143), .Z0_t (RoundOutput[118]), .Z0_f (new_AGEMA_signal_17306), .Z1_t (new_AGEMA_signal_17307), .Z1_f (new_AGEMA_signal_17308) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1182 ( .A0_t (MixColumnsOutput[119]), .A0_f (new_AGEMA_signal_15860), .A1_t (new_AGEMA_signal_15861), .A1_f (new_AGEMA_signal_15862), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n638), .Z0_f (new_AGEMA_signal_16613), .Z1_t (new_AGEMA_signal_16614), .Z1_f (new_AGEMA_signal_16615) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1183 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13850), .B1_t (new_AGEMA_signal_13851), .B1_f (new_AGEMA_signal_13852), .Z0_t (n637), .Z0_f (new_AGEMA_signal_14144), .Z1_t (new_AGEMA_signal_14145), .Z1_f (new_AGEMA_signal_14146) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1184 ( .A0_t (n638), .A0_f (new_AGEMA_signal_16613), .A1_t (new_AGEMA_signal_16614), .A1_f (new_AGEMA_signal_16615), .B0_t (n637), .B0_f (new_AGEMA_signal_14144), .B1_t (new_AGEMA_signal_14145), .B1_f (new_AGEMA_signal_14146), .Z0_t (RoundOutput[119]), .Z0_f (new_AGEMA_signal_17309), .Z1_t (new_AGEMA_signal_17310), .Z1_f (new_AGEMA_signal_17311) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1185 ( .A0_t (MixColumnsOutput[11]), .A0_f (new_AGEMA_signal_16952), .A1_t (new_AGEMA_signal_16953), .A1_f (new_AGEMA_signal_16954), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n640), .Z0_f (new_AGEMA_signal_17312), .Z1_t (new_AGEMA_signal_17313), .Z1_f (new_AGEMA_signal_17314) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1186 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[11]), .B0_f (new_AGEMA_signal_13841), .B1_t (new_AGEMA_signal_13842), .B1_f (new_AGEMA_signal_13843), .Z0_t (n639), .Z0_f (new_AGEMA_signal_14147), .Z1_t (new_AGEMA_signal_14148), .Z1_f (new_AGEMA_signal_14149) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1187 ( .A0_t (n640), .A0_f (new_AGEMA_signal_17312), .A1_t (new_AGEMA_signal_17313), .A1_f (new_AGEMA_signal_17314), .B0_t (n639), .B0_f (new_AGEMA_signal_14147), .B1_t (new_AGEMA_signal_14148), .B1_f (new_AGEMA_signal_14149), .Z0_t (RoundOutput[11]), .Z0_f (new_AGEMA_signal_17780), .Z1_t (new_AGEMA_signal_17781), .Z1_f (new_AGEMA_signal_17782) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1188 ( .A0_t (MixColumnsOutput[120]), .A0_f (new_AGEMA_signal_15857), .A1_t (new_AGEMA_signal_15858), .A1_f (new_AGEMA_signal_15859), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n642), .Z0_f (new_AGEMA_signal_16616), .Z1_t (new_AGEMA_signal_16617), .Z1_f (new_AGEMA_signal_16618) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1189 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[120]), .B0_f (new_AGEMA_signal_13493), .B1_t (new_AGEMA_signal_13494), .B1_f (new_AGEMA_signal_13495), .Z0_t (n641), .Z0_f (new_AGEMA_signal_13601), .Z1_t (new_AGEMA_signal_13602), .Z1_f (new_AGEMA_signal_13603) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1190 ( .A0_t (n642), .A0_f (new_AGEMA_signal_16616), .A1_t (new_AGEMA_signal_16617), .A1_f (new_AGEMA_signal_16618), .B0_t (n641), .B0_f (new_AGEMA_signal_13601), .B1_t (new_AGEMA_signal_13602), .B1_f (new_AGEMA_signal_13603), .Z0_t (RoundOutput[120]), .Z0_f (new_AGEMA_signal_17315), .Z1_t (new_AGEMA_signal_17316), .Z1_f (new_AGEMA_signal_17317) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1191 ( .A0_t (MixColumnsOutput[121]), .A0_f (new_AGEMA_signal_16826), .A1_t (new_AGEMA_signal_16827), .A1_f (new_AGEMA_signal_16828), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n644), .Z0_f (new_AGEMA_signal_17318), .Z1_t (new_AGEMA_signal_17319), .Z1_f (new_AGEMA_signal_17320) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1192 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13973), .B1_t (new_AGEMA_signal_13974), .B1_f (new_AGEMA_signal_13975), .Z0_t (n643), .Z0_f (new_AGEMA_signal_14150), .Z1_t (new_AGEMA_signal_14151), .Z1_f (new_AGEMA_signal_14152) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1193 ( .A0_t (n644), .A0_f (new_AGEMA_signal_17318), .A1_t (new_AGEMA_signal_17319), .A1_f (new_AGEMA_signal_17320), .B0_t (n643), .B0_f (new_AGEMA_signal_14150), .B1_t (new_AGEMA_signal_14151), .B1_f (new_AGEMA_signal_14152), .Z0_t (RoundOutput[121]), .Z0_f (new_AGEMA_signal_17783), .Z1_t (new_AGEMA_signal_17784), .Z1_f (new_AGEMA_signal_17785) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1194 ( .A0_t (MixColumnsOutput[122]), .A0_f (new_AGEMA_signal_15851), .A1_t (new_AGEMA_signal_15852), .A1_f (new_AGEMA_signal_15853), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n646), .Z0_f (new_AGEMA_signal_16619), .Z1_t (new_AGEMA_signal_16620), .Z1_f (new_AGEMA_signal_16621) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1195 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[122]), .B0_f (new_AGEMA_signal_13970), .B1_t (new_AGEMA_signal_13971), .B1_f (new_AGEMA_signal_13972), .Z0_t (n645), .Z0_f (new_AGEMA_signal_14153), .Z1_t (new_AGEMA_signal_14154), .Z1_f (new_AGEMA_signal_14155) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1196 ( .A0_t (n646), .A0_f (new_AGEMA_signal_16619), .A1_t (new_AGEMA_signal_16620), .A1_f (new_AGEMA_signal_16621), .B0_t (n645), .B0_f (new_AGEMA_signal_14153), .B1_t (new_AGEMA_signal_14154), .B1_f (new_AGEMA_signal_14155), .Z0_t (RoundOutput[122]), .Z0_f (new_AGEMA_signal_17321), .Z1_t (new_AGEMA_signal_17322), .Z1_f (new_AGEMA_signal_17323) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1197 ( .A0_t (MixColumnsOutput[123]), .A0_f (new_AGEMA_signal_16823), .A1_t (new_AGEMA_signal_16824), .A1_f (new_AGEMA_signal_16825), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n648), .Z0_f (new_AGEMA_signal_17324), .Z1_t (new_AGEMA_signal_17325), .Z1_f (new_AGEMA_signal_17326) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1198 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[123]), .B0_f (new_AGEMA_signal_13967), .B1_t (new_AGEMA_signal_13968), .B1_f (new_AGEMA_signal_13969), .Z0_t (n647), .Z0_f (new_AGEMA_signal_14156), .Z1_t (new_AGEMA_signal_14157), .Z1_f (new_AGEMA_signal_14158) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1199 ( .A0_t (n648), .A0_f (new_AGEMA_signal_17324), .A1_t (new_AGEMA_signal_17325), .A1_f (new_AGEMA_signal_17326), .B0_t (n647), .B0_f (new_AGEMA_signal_14156), .B1_t (new_AGEMA_signal_14157), .B1_f (new_AGEMA_signal_14158), .Z0_t (RoundOutput[123]), .Z0_f (new_AGEMA_signal_17786), .Z1_t (new_AGEMA_signal_17787), .Z1_f (new_AGEMA_signal_17788) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1200 ( .A0_t (MixColumnsOutput[124]), .A0_f (new_AGEMA_signal_16820), .A1_t (new_AGEMA_signal_16821), .A1_f (new_AGEMA_signal_16822), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n650), .Z0_f (new_AGEMA_signal_17327), .Z1_t (new_AGEMA_signal_17328), .Z1_f (new_AGEMA_signal_17329) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1201 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13964), .B1_t (new_AGEMA_signal_13965), .B1_f (new_AGEMA_signal_13966), .Z0_t (n649), .Z0_f (new_AGEMA_signal_14159), .Z1_t (new_AGEMA_signal_14160), .Z1_f (new_AGEMA_signal_14161) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1202 ( .A0_t (n650), .A0_f (new_AGEMA_signal_17327), .A1_t (new_AGEMA_signal_17328), .A1_f (new_AGEMA_signal_17329), .B0_t (n649), .B0_f (new_AGEMA_signal_14159), .B1_t (new_AGEMA_signal_14160), .B1_f (new_AGEMA_signal_14161), .Z0_t (RoundOutput[124]), .Z0_f (new_AGEMA_signal_17789), .Z1_t (new_AGEMA_signal_17790), .Z1_f (new_AGEMA_signal_17791) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1203 ( .A0_t (MixColumnsOutput[125]), .A0_f (new_AGEMA_signal_15842), .A1_t (new_AGEMA_signal_15843), .A1_f (new_AGEMA_signal_15844), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n652), .Z0_f (new_AGEMA_signal_16622), .Z1_t (new_AGEMA_signal_16623), .Z1_f (new_AGEMA_signal_16624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1204 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13961), .B1_t (new_AGEMA_signal_13962), .B1_f (new_AGEMA_signal_13963), .Z0_t (n651), .Z0_f (new_AGEMA_signal_14162), .Z1_t (new_AGEMA_signal_14163), .Z1_f (new_AGEMA_signal_14164) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1205 ( .A0_t (n652), .A0_f (new_AGEMA_signal_16622), .A1_t (new_AGEMA_signal_16623), .A1_f (new_AGEMA_signal_16624), .B0_t (n651), .B0_f (new_AGEMA_signal_14162), .B1_t (new_AGEMA_signal_14163), .B1_f (new_AGEMA_signal_14164), .Z0_t (RoundOutput[125]), .Z0_f (new_AGEMA_signal_17330), .Z1_t (new_AGEMA_signal_17331), .Z1_f (new_AGEMA_signal_17332) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1206 ( .A0_t (MixColumnsOutput[126]), .A0_f (new_AGEMA_signal_15836), .A1_t (new_AGEMA_signal_15837), .A1_f (new_AGEMA_signal_15838), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n654), .Z0_f (new_AGEMA_signal_16625), .Z1_t (new_AGEMA_signal_16626), .Z1_f (new_AGEMA_signal_16627) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1207 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13958), .B1_t (new_AGEMA_signal_13959), .B1_f (new_AGEMA_signal_13960), .Z0_t (n653), .Z0_f (new_AGEMA_signal_14165), .Z1_t (new_AGEMA_signal_14166), .Z1_f (new_AGEMA_signal_14167) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1208 ( .A0_t (n654), .A0_f (new_AGEMA_signal_16625), .A1_t (new_AGEMA_signal_16626), .A1_f (new_AGEMA_signal_16627), .B0_t (n653), .B0_f (new_AGEMA_signal_14165), .B1_t (new_AGEMA_signal_14166), .B1_f (new_AGEMA_signal_14167), .Z0_t (RoundOutput[126]), .Z0_f (new_AGEMA_signal_17333), .Z1_t (new_AGEMA_signal_17334), .Z1_f (new_AGEMA_signal_17335) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1209 ( .A0_t (MixColumnsOutput[127]), .A0_f (new_AGEMA_signal_15833), .A1_t (new_AGEMA_signal_15834), .A1_f (new_AGEMA_signal_15835), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n656), .Z0_f (new_AGEMA_signal_16628), .Z1_t (new_AGEMA_signal_16629), .Z1_f (new_AGEMA_signal_16630) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1210 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13955), .B1_t (new_AGEMA_signal_13956), .B1_f (new_AGEMA_signal_13957), .Z0_t (n655), .Z0_f (new_AGEMA_signal_14168), .Z1_t (new_AGEMA_signal_14169), .Z1_f (new_AGEMA_signal_14170) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1211 ( .A0_t (n656), .A0_f (new_AGEMA_signal_16628), .A1_t (new_AGEMA_signal_16629), .A1_f (new_AGEMA_signal_16630), .B0_t (n655), .B0_f (new_AGEMA_signal_14168), .B1_t (new_AGEMA_signal_14169), .B1_f (new_AGEMA_signal_14170), .Z0_t (RoundOutput[127]), .Z0_f (new_AGEMA_signal_17336), .Z1_t (new_AGEMA_signal_17337), .Z1_f (new_AGEMA_signal_17338) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1212 ( .A0_t (MixColumnsOutput[12]), .A0_f (new_AGEMA_signal_16949), .A1_t (new_AGEMA_signal_16950), .A1_f (new_AGEMA_signal_16951), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n658), .Z0_f (new_AGEMA_signal_17339), .Z1_t (new_AGEMA_signal_17340), .Z1_f (new_AGEMA_signal_17341) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1213 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13838), .B1_t (new_AGEMA_signal_13839), .B1_f (new_AGEMA_signal_13840), .Z0_t (n657), .Z0_f (new_AGEMA_signal_14171), .Z1_t (new_AGEMA_signal_14172), .Z1_f (new_AGEMA_signal_14173) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1214 ( .A0_t (n658), .A0_f (new_AGEMA_signal_17339), .A1_t (new_AGEMA_signal_17340), .A1_f (new_AGEMA_signal_17341), .B0_t (n657), .B0_f (new_AGEMA_signal_14171), .B1_t (new_AGEMA_signal_14172), .B1_f (new_AGEMA_signal_14173), .Z0_t (RoundOutput[12]), .Z0_f (new_AGEMA_signal_17792), .Z1_t (new_AGEMA_signal_17793), .Z1_f (new_AGEMA_signal_17794) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1215 ( .A0_t (MixColumnsOutput[13]), .A0_f (new_AGEMA_signal_16181), .A1_t (new_AGEMA_signal_16182), .A1_f (new_AGEMA_signal_16183), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n660), .Z0_f (new_AGEMA_signal_16631), .Z1_t (new_AGEMA_signal_16632), .Z1_f (new_AGEMA_signal_16633) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1216 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13835), .B1_t (new_AGEMA_signal_13836), .B1_f (new_AGEMA_signal_13837), .Z0_t (n659), .Z0_f (new_AGEMA_signal_14174), .Z1_t (new_AGEMA_signal_14175), .Z1_f (new_AGEMA_signal_14176) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1217 ( .A0_t (n660), .A0_f (new_AGEMA_signal_16631), .A1_t (new_AGEMA_signal_16632), .A1_f (new_AGEMA_signal_16633), .B0_t (n659), .B0_f (new_AGEMA_signal_14174), .B1_t (new_AGEMA_signal_14175), .B1_f (new_AGEMA_signal_14176), .Z0_t (RoundOutput[13]), .Z0_f (new_AGEMA_signal_17342), .Z1_t (new_AGEMA_signal_17343), .Z1_f (new_AGEMA_signal_17344) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1218 ( .A0_t (MixColumnsOutput[14]), .A0_f (new_AGEMA_signal_16178), .A1_t (new_AGEMA_signal_16179), .A1_f (new_AGEMA_signal_16180), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n662), .Z0_f (new_AGEMA_signal_16634), .Z1_t (new_AGEMA_signal_16635), .Z1_f (new_AGEMA_signal_16636) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1219 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13832), .B1_t (new_AGEMA_signal_13833), .B1_f (new_AGEMA_signal_13834), .Z0_t (n661), .Z0_f (new_AGEMA_signal_14177), .Z1_t (new_AGEMA_signal_14178), .Z1_f (new_AGEMA_signal_14179) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1220 ( .A0_t (n662), .A0_f (new_AGEMA_signal_16634), .A1_t (new_AGEMA_signal_16635), .A1_f (new_AGEMA_signal_16636), .B0_t (n661), .B0_f (new_AGEMA_signal_14177), .B1_t (new_AGEMA_signal_14178), .B1_f (new_AGEMA_signal_14179), .Z0_t (RoundOutput[14]), .Z0_f (new_AGEMA_signal_17345), .Z1_t (new_AGEMA_signal_17346), .Z1_f (new_AGEMA_signal_17347) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1221 ( .A0_t (MixColumnsOutput[15]), .A0_f (new_AGEMA_signal_16175), .A1_t (new_AGEMA_signal_16176), .A1_f (new_AGEMA_signal_16177), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n664), .Z0_f (new_AGEMA_signal_16637), .Z1_t (new_AGEMA_signal_16638), .Z1_f (new_AGEMA_signal_16639) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1222 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B0_f (new_AGEMA_signal_13829), .B1_t (new_AGEMA_signal_13830), .B1_f (new_AGEMA_signal_13831), .Z0_t (n663), .Z0_f (new_AGEMA_signal_14180), .Z1_t (new_AGEMA_signal_14181), .Z1_f (new_AGEMA_signal_14182) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1223 ( .A0_t (n664), .A0_f (new_AGEMA_signal_16637), .A1_t (new_AGEMA_signal_16638), .A1_f (new_AGEMA_signal_16639), .B0_t (n663), .B0_f (new_AGEMA_signal_14180), .B1_t (new_AGEMA_signal_14181), .B1_f (new_AGEMA_signal_14182), .Z0_t (RoundOutput[15]), .Z0_f (new_AGEMA_signal_17348), .Z1_t (new_AGEMA_signal_17349), .Z1_f (new_AGEMA_signal_17350) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1224 ( .A0_t (MixColumnsOutput[16]), .A0_f (new_AGEMA_signal_16172), .A1_t (new_AGEMA_signal_16173), .A1_f (new_AGEMA_signal_16174), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n666), .Z0_f (new_AGEMA_signal_16640), .Z1_t (new_AGEMA_signal_16641), .Z1_f (new_AGEMA_signal_16642) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1225 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[16]), .B0_f (new_AGEMA_signal_13460), .B1_t (new_AGEMA_signal_13461), .B1_f (new_AGEMA_signal_13462), .Z0_t (n665), .Z0_f (new_AGEMA_signal_13604), .Z1_t (new_AGEMA_signal_13605), .Z1_f (new_AGEMA_signal_13606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1226 ( .A0_t (n666), .A0_f (new_AGEMA_signal_16640), .A1_t (new_AGEMA_signal_16641), .A1_f (new_AGEMA_signal_16642), .B0_t (n665), .B0_f (new_AGEMA_signal_13604), .B1_t (new_AGEMA_signal_13605), .B1_f (new_AGEMA_signal_13606), .Z0_t (RoundOutput[16]), .Z0_f (new_AGEMA_signal_17351), .Z1_t (new_AGEMA_signal_17352), .Z1_f (new_AGEMA_signal_17353) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1227 ( .A0_t (MixColumnsOutput[17]), .A0_f (new_AGEMA_signal_16946), .A1_t (new_AGEMA_signal_16947), .A1_f (new_AGEMA_signal_16948), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n668), .Z0_f (new_AGEMA_signal_17354), .Z1_t (new_AGEMA_signal_17355), .Z1_f (new_AGEMA_signal_17356) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1228 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13952), .B1_t (new_AGEMA_signal_13953), .B1_f (new_AGEMA_signal_13954), .Z0_t (n667), .Z0_f (new_AGEMA_signal_14183), .Z1_t (new_AGEMA_signal_14184), .Z1_f (new_AGEMA_signal_14185) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1229 ( .A0_t (n668), .A0_f (new_AGEMA_signal_17354), .A1_t (new_AGEMA_signal_17355), .A1_f (new_AGEMA_signal_17356), .B0_t (n667), .B0_f (new_AGEMA_signal_14183), .B1_t (new_AGEMA_signal_14184), .B1_f (new_AGEMA_signal_14185), .Z0_t (RoundOutput[17]), .Z0_f (new_AGEMA_signal_17795), .Z1_t (new_AGEMA_signal_17796), .Z1_f (new_AGEMA_signal_17797) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1230 ( .A0_t (MixColumnsOutput[18]), .A0_f (new_AGEMA_signal_16166), .A1_t (new_AGEMA_signal_16167), .A1_f (new_AGEMA_signal_16168), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n670), .Z0_f (new_AGEMA_signal_16643), .Z1_t (new_AGEMA_signal_16644), .Z1_f (new_AGEMA_signal_16645) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1231 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[18]), .B0_f (new_AGEMA_signal_13949), .B1_t (new_AGEMA_signal_13950), .B1_f (new_AGEMA_signal_13951), .Z0_t (n669), .Z0_f (new_AGEMA_signal_14186), .Z1_t (new_AGEMA_signal_14187), .Z1_f (new_AGEMA_signal_14188) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1232 ( .A0_t (n670), .A0_f (new_AGEMA_signal_16643), .A1_t (new_AGEMA_signal_16644), .A1_f (new_AGEMA_signal_16645), .B0_t (n669), .B0_f (new_AGEMA_signal_14186), .B1_t (new_AGEMA_signal_14187), .B1_f (new_AGEMA_signal_14188), .Z0_t (RoundOutput[18]), .Z0_f (new_AGEMA_signal_17357), .Z1_t (new_AGEMA_signal_17358), .Z1_f (new_AGEMA_signal_17359) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1233 ( .A0_t (MixColumnsOutput[19]), .A0_f (new_AGEMA_signal_16943), .A1_t (new_AGEMA_signal_16944), .A1_f (new_AGEMA_signal_16945), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n672), .Z0_f (new_AGEMA_signal_17360), .Z1_t (new_AGEMA_signal_17361), .Z1_f (new_AGEMA_signal_17362) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1234 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[19]), .B0_f (new_AGEMA_signal_13946), .B1_t (new_AGEMA_signal_13947), .B1_f (new_AGEMA_signal_13948), .Z0_t (n671), .Z0_f (new_AGEMA_signal_14189), .Z1_t (new_AGEMA_signal_14190), .Z1_f (new_AGEMA_signal_14191) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1235 ( .A0_t (n672), .A0_f (new_AGEMA_signal_17360), .A1_t (new_AGEMA_signal_17361), .A1_f (new_AGEMA_signal_17362), .B0_t (n671), .B0_f (new_AGEMA_signal_14189), .B1_t (new_AGEMA_signal_14190), .B1_f (new_AGEMA_signal_14191), .Z0_t (RoundOutput[19]), .Z0_f (new_AGEMA_signal_17798), .Z1_t (new_AGEMA_signal_17799), .Z1_f (new_AGEMA_signal_17800) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1236 ( .A0_t (MixColumnsOutput[1]), .A0_f (new_AGEMA_signal_16940), .A1_t (new_AGEMA_signal_16941), .A1_f (new_AGEMA_signal_16942), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n674), .Z0_f (new_AGEMA_signal_17363), .Z1_t (new_AGEMA_signal_17364), .Z1_f (new_AGEMA_signal_17365) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1237 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .B0_f (new_AGEMA_signal_13742), .B1_t (new_AGEMA_signal_13743), .B1_f (new_AGEMA_signal_13744), .Z0_t (n673), .Z0_f (new_AGEMA_signal_14192), .Z1_t (new_AGEMA_signal_14193), .Z1_f (new_AGEMA_signal_14194) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1238 ( .A0_t (n674), .A0_f (new_AGEMA_signal_17363), .A1_t (new_AGEMA_signal_17364), .A1_f (new_AGEMA_signal_17365), .B0_t (n673), .B0_f (new_AGEMA_signal_14192), .B1_t (new_AGEMA_signal_14193), .B1_f (new_AGEMA_signal_14194), .Z0_t (RoundOutput[1]), .Z0_f (new_AGEMA_signal_17801), .Z1_t (new_AGEMA_signal_17802), .Z1_f (new_AGEMA_signal_17803) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1239 ( .A0_t (MixColumnsOutput[20]), .A0_f (new_AGEMA_signal_16937), .A1_t (new_AGEMA_signal_16938), .A1_f (new_AGEMA_signal_16939), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n676), .Z0_f (new_AGEMA_signal_17366), .Z1_t (new_AGEMA_signal_17367), .Z1_f (new_AGEMA_signal_17368) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1240 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13943), .B1_t (new_AGEMA_signal_13944), .B1_f (new_AGEMA_signal_13945), .Z0_t (n675), .Z0_f (new_AGEMA_signal_14195), .Z1_t (new_AGEMA_signal_14196), .Z1_f (new_AGEMA_signal_14197) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1241 ( .A0_t (n676), .A0_f (new_AGEMA_signal_17366), .A1_t (new_AGEMA_signal_17367), .A1_f (new_AGEMA_signal_17368), .B0_t (n675), .B0_f (new_AGEMA_signal_14195), .B1_t (new_AGEMA_signal_14196), .B1_f (new_AGEMA_signal_14197), .Z0_t (RoundOutput[20]), .Z0_f (new_AGEMA_signal_17804), .Z1_t (new_AGEMA_signal_17805), .Z1_f (new_AGEMA_signal_17806) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1242 ( .A0_t (MixColumnsOutput[21]), .A0_f (new_AGEMA_signal_16154), .A1_t (new_AGEMA_signal_16155), .A1_f (new_AGEMA_signal_16156), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n678), .Z0_f (new_AGEMA_signal_16646), .Z1_t (new_AGEMA_signal_16647), .Z1_f (new_AGEMA_signal_16648) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1243 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13940), .B1_t (new_AGEMA_signal_13941), .B1_f (new_AGEMA_signal_13942), .Z0_t (n677), .Z0_f (new_AGEMA_signal_14198), .Z1_t (new_AGEMA_signal_14199), .Z1_f (new_AGEMA_signal_14200) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1244 ( .A0_t (n678), .A0_f (new_AGEMA_signal_16646), .A1_t (new_AGEMA_signal_16647), .A1_f (new_AGEMA_signal_16648), .B0_t (n677), .B0_f (new_AGEMA_signal_14198), .B1_t (new_AGEMA_signal_14199), .B1_f (new_AGEMA_signal_14200), .Z0_t (RoundOutput[21]), .Z0_f (new_AGEMA_signal_17369), .Z1_t (new_AGEMA_signal_17370), .Z1_f (new_AGEMA_signal_17371) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1245 ( .A0_t (MixColumnsOutput[22]), .A0_f (new_AGEMA_signal_16151), .A1_t (new_AGEMA_signal_16152), .A1_f (new_AGEMA_signal_16153), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n680), .Z0_f (new_AGEMA_signal_16649), .Z1_t (new_AGEMA_signal_16650), .Z1_f (new_AGEMA_signal_16651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1246 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13937), .B1_t (new_AGEMA_signal_13938), .B1_f (new_AGEMA_signal_13939), .Z0_t (n679), .Z0_f (new_AGEMA_signal_14201), .Z1_t (new_AGEMA_signal_14202), .Z1_f (new_AGEMA_signal_14203) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1247 ( .A0_t (n680), .A0_f (new_AGEMA_signal_16649), .A1_t (new_AGEMA_signal_16650), .A1_f (new_AGEMA_signal_16651), .B0_t (n679), .B0_f (new_AGEMA_signal_14201), .B1_t (new_AGEMA_signal_14202), .B1_f (new_AGEMA_signal_14203), .Z0_t (RoundOutput[22]), .Z0_f (new_AGEMA_signal_17372), .Z1_t (new_AGEMA_signal_17373), .Z1_f (new_AGEMA_signal_17374) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1248 ( .A0_t (MixColumnsOutput[23]), .A0_f (new_AGEMA_signal_16148), .A1_t (new_AGEMA_signal_16149), .A1_f (new_AGEMA_signal_16150), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n682), .Z0_f (new_AGEMA_signal_16652), .Z1_t (new_AGEMA_signal_16653), .Z1_f (new_AGEMA_signal_16654) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1249 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13934), .B1_t (new_AGEMA_signal_13935), .B1_f (new_AGEMA_signal_13936), .Z0_t (n681), .Z0_f (new_AGEMA_signal_14204), .Z1_t (new_AGEMA_signal_14205), .Z1_f (new_AGEMA_signal_14206) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1250 ( .A0_t (n682), .A0_f (new_AGEMA_signal_16652), .A1_t (new_AGEMA_signal_16653), .A1_f (new_AGEMA_signal_16654), .B0_t (n681), .B0_f (new_AGEMA_signal_14204), .B1_t (new_AGEMA_signal_14205), .B1_f (new_AGEMA_signal_14206), .Z0_t (RoundOutput[23]), .Z0_f (new_AGEMA_signal_17375), .Z1_t (new_AGEMA_signal_17376), .Z1_f (new_AGEMA_signal_17377) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1251 ( .A0_t (MixColumnsOutput[24]), .A0_f (new_AGEMA_signal_16145), .A1_t (new_AGEMA_signal_16146), .A1_f (new_AGEMA_signal_16147), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n684), .Z0_f (new_AGEMA_signal_16655), .Z1_t (new_AGEMA_signal_16656), .Z1_f (new_AGEMA_signal_16657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1252 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[24]), .B0_f (new_AGEMA_signal_13097), .B1_t (new_AGEMA_signal_13098), .B1_f (new_AGEMA_signal_13099), .Z0_t (n683), .Z0_f (new_AGEMA_signal_13607), .Z1_t (new_AGEMA_signal_13608), .Z1_f (new_AGEMA_signal_13609) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1253 ( .A0_t (n684), .A0_f (new_AGEMA_signal_16655), .A1_t (new_AGEMA_signal_16656), .A1_f (new_AGEMA_signal_16657), .B0_t (n683), .B0_f (new_AGEMA_signal_13607), .B1_t (new_AGEMA_signal_13608), .B1_f (new_AGEMA_signal_13609), .Z0_t (RoundOutput[24]), .Z0_f (new_AGEMA_signal_17378), .Z1_t (new_AGEMA_signal_17379), .Z1_f (new_AGEMA_signal_17380) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1254 ( .A0_t (MixColumnsOutput[25]), .A0_f (new_AGEMA_signal_16934), .A1_t (new_AGEMA_signal_16935), .A1_f (new_AGEMA_signal_16936), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n686), .Z0_f (new_AGEMA_signal_17381), .Z1_t (new_AGEMA_signal_17382), .Z1_f (new_AGEMA_signal_17383) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1255 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13721), .B1_t (new_AGEMA_signal_13722), .B1_f (new_AGEMA_signal_13723), .Z0_t (n685), .Z0_f (new_AGEMA_signal_14207), .Z1_t (new_AGEMA_signal_14208), .Z1_f (new_AGEMA_signal_14209) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1256 ( .A0_t (n686), .A0_f (new_AGEMA_signal_17381), .A1_t (new_AGEMA_signal_17382), .A1_f (new_AGEMA_signal_17383), .B0_t (n685), .B0_f (new_AGEMA_signal_14207), .B1_t (new_AGEMA_signal_14208), .B1_f (new_AGEMA_signal_14209), .Z0_t (RoundOutput[25]), .Z0_f (new_AGEMA_signal_17807), .Z1_t (new_AGEMA_signal_17808), .Z1_f (new_AGEMA_signal_17809) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1257 ( .A0_t (MixColumnsOutput[26]), .A0_f (new_AGEMA_signal_16139), .A1_t (new_AGEMA_signal_16140), .A1_f (new_AGEMA_signal_16141), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n688), .Z0_f (new_AGEMA_signal_16658), .Z1_t (new_AGEMA_signal_16659), .Z1_f (new_AGEMA_signal_16660) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1258 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[26]), .B0_f (new_AGEMA_signal_13718), .B1_t (new_AGEMA_signal_13719), .B1_f (new_AGEMA_signal_13720), .Z0_t (n687), .Z0_f (new_AGEMA_signal_14210), .Z1_t (new_AGEMA_signal_14211), .Z1_f (new_AGEMA_signal_14212) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1259 ( .A0_t (n688), .A0_f (new_AGEMA_signal_16658), .A1_t (new_AGEMA_signal_16659), .A1_f (new_AGEMA_signal_16660), .B0_t (n687), .B0_f (new_AGEMA_signal_14210), .B1_t (new_AGEMA_signal_14211), .B1_f (new_AGEMA_signal_14212), .Z0_t (RoundOutput[26]), .Z0_f (new_AGEMA_signal_17384), .Z1_t (new_AGEMA_signal_17385), .Z1_f (new_AGEMA_signal_17386) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1260 ( .A0_t (MixColumnsOutput[27]), .A0_f (new_AGEMA_signal_16931), .A1_t (new_AGEMA_signal_16932), .A1_f (new_AGEMA_signal_16933), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n690), .Z0_f (new_AGEMA_signal_17387), .Z1_t (new_AGEMA_signal_17388), .Z1_f (new_AGEMA_signal_17389) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1261 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[27]), .B0_f (new_AGEMA_signal_13715), .B1_t (new_AGEMA_signal_13716), .B1_f (new_AGEMA_signal_13717), .Z0_t (n689), .Z0_f (new_AGEMA_signal_14213), .Z1_t (new_AGEMA_signal_14214), .Z1_f (new_AGEMA_signal_14215) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1262 ( .A0_t (n690), .A0_f (new_AGEMA_signal_17387), .A1_t (new_AGEMA_signal_17388), .A1_f (new_AGEMA_signal_17389), .B0_t (n689), .B0_f (new_AGEMA_signal_14213), .B1_t (new_AGEMA_signal_14214), .B1_f (new_AGEMA_signal_14215), .Z0_t (RoundOutput[27]), .Z0_f (new_AGEMA_signal_17810), .Z1_t (new_AGEMA_signal_17811), .Z1_f (new_AGEMA_signal_17812) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1263 ( .A0_t (MixColumnsOutput[28]), .A0_f (new_AGEMA_signal_16928), .A1_t (new_AGEMA_signal_16929), .A1_f (new_AGEMA_signal_16930), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n692), .Z0_f (new_AGEMA_signal_17390), .Z1_t (new_AGEMA_signal_17391), .Z1_f (new_AGEMA_signal_17392) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1264 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13712), .B1_t (new_AGEMA_signal_13713), .B1_f (new_AGEMA_signal_13714), .Z0_t (n691), .Z0_f (new_AGEMA_signal_14216), .Z1_t (new_AGEMA_signal_14217), .Z1_f (new_AGEMA_signal_14218) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1265 ( .A0_t (n692), .A0_f (new_AGEMA_signal_17390), .A1_t (new_AGEMA_signal_17391), .A1_f (new_AGEMA_signal_17392), .B0_t (n691), .B0_f (new_AGEMA_signal_14216), .B1_t (new_AGEMA_signal_14217), .B1_f (new_AGEMA_signal_14218), .Z0_t (RoundOutput[28]), .Z0_f (new_AGEMA_signal_17813), .Z1_t (new_AGEMA_signal_17814), .Z1_f (new_AGEMA_signal_17815) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1266 ( .A0_t (MixColumnsOutput[29]), .A0_f (new_AGEMA_signal_16130), .A1_t (new_AGEMA_signal_16131), .A1_f (new_AGEMA_signal_16132), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n694), .Z0_f (new_AGEMA_signal_16661), .Z1_t (new_AGEMA_signal_16662), .Z1_f (new_AGEMA_signal_16663) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1267 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13709), .B1_t (new_AGEMA_signal_13710), .B1_f (new_AGEMA_signal_13711), .Z0_t (n693), .Z0_f (new_AGEMA_signal_14219), .Z1_t (new_AGEMA_signal_14220), .Z1_f (new_AGEMA_signal_14221) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1268 ( .A0_t (n694), .A0_f (new_AGEMA_signal_16661), .A1_t (new_AGEMA_signal_16662), .A1_f (new_AGEMA_signal_16663), .B0_t (n693), .B0_f (new_AGEMA_signal_14219), .B1_t (new_AGEMA_signal_14220), .B1_f (new_AGEMA_signal_14221), .Z0_t (RoundOutput[29]), .Z0_f (new_AGEMA_signal_17393), .Z1_t (new_AGEMA_signal_17394), .Z1_f (new_AGEMA_signal_17395) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1269 ( .A0_t (MixColumnsOutput[2]), .A0_f (new_AGEMA_signal_16127), .A1_t (new_AGEMA_signal_16128), .A1_f (new_AGEMA_signal_16129), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n696), .Z0_f (new_AGEMA_signal_16664), .Z1_t (new_AGEMA_signal_16665), .Z1_f (new_AGEMA_signal_16666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1270 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[2]), .B0_f (new_AGEMA_signal_13739), .B1_t (new_AGEMA_signal_13740), .B1_f (new_AGEMA_signal_13741), .Z0_t (n695), .Z0_f (new_AGEMA_signal_14222), .Z1_t (new_AGEMA_signal_14223), .Z1_f (new_AGEMA_signal_14224) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1271 ( .A0_t (n696), .A0_f (new_AGEMA_signal_16664), .A1_t (new_AGEMA_signal_16665), .A1_f (new_AGEMA_signal_16666), .B0_t (n695), .B0_f (new_AGEMA_signal_14222), .B1_t (new_AGEMA_signal_14223), .B1_f (new_AGEMA_signal_14224), .Z0_t (RoundOutput[2]), .Z0_f (new_AGEMA_signal_17396), .Z1_t (new_AGEMA_signal_17397), .Z1_f (new_AGEMA_signal_17398) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1272 ( .A0_t (MixColumnsOutput[30]), .A0_f (new_AGEMA_signal_16124), .A1_t (new_AGEMA_signal_16125), .A1_f (new_AGEMA_signal_16126), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n698), .Z0_f (new_AGEMA_signal_16667), .Z1_t (new_AGEMA_signal_16668), .Z1_f (new_AGEMA_signal_16669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1273 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13706), .B1_t (new_AGEMA_signal_13707), .B1_f (new_AGEMA_signal_13708), .Z0_t (n697), .Z0_f (new_AGEMA_signal_14225), .Z1_t (new_AGEMA_signal_14226), .Z1_f (new_AGEMA_signal_14227) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1274 ( .A0_t (n698), .A0_f (new_AGEMA_signal_16667), .A1_t (new_AGEMA_signal_16668), .A1_f (new_AGEMA_signal_16669), .B0_t (n697), .B0_f (new_AGEMA_signal_14225), .B1_t (new_AGEMA_signal_14226), .B1_f (new_AGEMA_signal_14227), .Z0_t (RoundOutput[30]), .Z0_f (new_AGEMA_signal_17399), .Z1_t (new_AGEMA_signal_17400), .Z1_f (new_AGEMA_signal_17401) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1275 ( .A0_t (MixColumnsOutput[31]), .A0_f (new_AGEMA_signal_16121), .A1_t (new_AGEMA_signal_16122), .A1_f (new_AGEMA_signal_16123), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n700), .Z0_f (new_AGEMA_signal_16670), .Z1_t (new_AGEMA_signal_16671), .Z1_f (new_AGEMA_signal_16672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1276 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13703), .B1_t (new_AGEMA_signal_13704), .B1_f (new_AGEMA_signal_13705), .Z0_t (n699), .Z0_f (new_AGEMA_signal_14228), .Z1_t (new_AGEMA_signal_14229), .Z1_f (new_AGEMA_signal_14230) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1277 ( .A0_t (n700), .A0_f (new_AGEMA_signal_16670), .A1_t (new_AGEMA_signal_16671), .A1_f (new_AGEMA_signal_16672), .B0_t (n699), .B0_f (new_AGEMA_signal_14228), .B1_t (new_AGEMA_signal_14229), .B1_f (new_AGEMA_signal_14230), .Z0_t (RoundOutput[31]), .Z0_f (new_AGEMA_signal_17402), .Z1_t (new_AGEMA_signal_17403), .Z1_f (new_AGEMA_signal_17404) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1278 ( .A0_t (MixColumnsOutput[32]), .A0_f (new_AGEMA_signal_16097), .A1_t (new_AGEMA_signal_16098), .A1_f (new_AGEMA_signal_16099), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n702), .Z0_f (new_AGEMA_signal_16673), .Z1_t (new_AGEMA_signal_16674), .Z1_f (new_AGEMA_signal_16675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1279 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[32]), .B0_f (new_AGEMA_signal_13262), .B1_t (new_AGEMA_signal_13263), .B1_f (new_AGEMA_signal_13264), .Z0_t (n701), .Z0_f (new_AGEMA_signal_13610), .Z1_t (new_AGEMA_signal_13611), .Z1_f (new_AGEMA_signal_13612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1280 ( .A0_t (n702), .A0_f (new_AGEMA_signal_16673), .A1_t (new_AGEMA_signal_16674), .A1_f (new_AGEMA_signal_16675), .B0_t (n701), .B0_f (new_AGEMA_signal_13610), .B1_t (new_AGEMA_signal_13611), .B1_f (new_AGEMA_signal_13612), .Z0_t (RoundOutput[32]), .Z0_f (new_AGEMA_signal_17405), .Z1_t (new_AGEMA_signal_17406), .Z1_f (new_AGEMA_signal_17407) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1281 ( .A0_t (MixColumnsOutput[33]), .A0_f (new_AGEMA_signal_16904), .A1_t (new_AGEMA_signal_16905), .A1_f (new_AGEMA_signal_16906), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n704), .Z0_f (new_AGEMA_signal_17408), .Z1_t (new_AGEMA_signal_17409), .Z1_f (new_AGEMA_signal_17410) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1282 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .B0_f (new_AGEMA_signal_13826), .B1_t (new_AGEMA_signal_13827), .B1_f (new_AGEMA_signal_13828), .Z0_t (n703), .Z0_f (new_AGEMA_signal_14231), .Z1_t (new_AGEMA_signal_14232), .Z1_f (new_AGEMA_signal_14233) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1283 ( .A0_t (n704), .A0_f (new_AGEMA_signal_17408), .A1_t (new_AGEMA_signal_17409), .A1_f (new_AGEMA_signal_17410), .B0_t (n703), .B0_f (new_AGEMA_signal_14231), .B1_t (new_AGEMA_signal_14232), .B1_f (new_AGEMA_signal_14233), .Z0_t (RoundOutput[33]), .Z0_f (new_AGEMA_signal_17816), .Z1_t (new_AGEMA_signal_17817), .Z1_f (new_AGEMA_signal_17818) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1284 ( .A0_t (MixColumnsOutput[34]), .A0_f (new_AGEMA_signal_16031), .A1_t (new_AGEMA_signal_16032), .A1_f (new_AGEMA_signal_16033), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n706), .Z0_f (new_AGEMA_signal_16676), .Z1_t (new_AGEMA_signal_16677), .Z1_f (new_AGEMA_signal_16678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1285 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[34]), .B0_f (new_AGEMA_signal_13823), .B1_t (new_AGEMA_signal_13824), .B1_f (new_AGEMA_signal_13825), .Z0_t (n705), .Z0_f (new_AGEMA_signal_14234), .Z1_t (new_AGEMA_signal_14235), .Z1_f (new_AGEMA_signal_14236) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1286 ( .A0_t (n706), .A0_f (new_AGEMA_signal_16676), .A1_t (new_AGEMA_signal_16677), .A1_f (new_AGEMA_signal_16678), .B0_t (n705), .B0_f (new_AGEMA_signal_14234), .B1_t (new_AGEMA_signal_14235), .B1_f (new_AGEMA_signal_14236), .Z0_t (RoundOutput[34]), .Z0_f (new_AGEMA_signal_17411), .Z1_t (new_AGEMA_signal_17412), .Z1_f (new_AGEMA_signal_17413) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1287 ( .A0_t (MixColumnsOutput[35]), .A0_f (new_AGEMA_signal_16889), .A1_t (new_AGEMA_signal_16890), .A1_f (new_AGEMA_signal_16891), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n708), .Z0_f (new_AGEMA_signal_17414), .Z1_t (new_AGEMA_signal_17415), .Z1_f (new_AGEMA_signal_17416) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1288 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[35]), .B0_f (new_AGEMA_signal_13820), .B1_t (new_AGEMA_signal_13821), .B1_f (new_AGEMA_signal_13822), .Z0_t (n707), .Z0_f (new_AGEMA_signal_14237), .Z1_t (new_AGEMA_signal_14238), .Z1_f (new_AGEMA_signal_14239) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1289 ( .A0_t (n708), .A0_f (new_AGEMA_signal_17414), .A1_t (new_AGEMA_signal_17415), .A1_f (new_AGEMA_signal_17416), .B0_t (n707), .B0_f (new_AGEMA_signal_14237), .B1_t (new_AGEMA_signal_14238), .B1_f (new_AGEMA_signal_14239), .Z0_t (RoundOutput[35]), .Z0_f (new_AGEMA_signal_17819), .Z1_t (new_AGEMA_signal_17820), .Z1_f (new_AGEMA_signal_17821) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1290 ( .A0_t (MixColumnsOutput[36]), .A0_f (new_AGEMA_signal_16886), .A1_t (new_AGEMA_signal_16887), .A1_f (new_AGEMA_signal_16888), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n710), .Z0_f (new_AGEMA_signal_17417), .Z1_t (new_AGEMA_signal_17418), .Z1_f (new_AGEMA_signal_17419) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1291 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .B0_f (new_AGEMA_signal_13817), .B1_t (new_AGEMA_signal_13818), .B1_f (new_AGEMA_signal_13819), .Z0_t (n709), .Z0_f (new_AGEMA_signal_14240), .Z1_t (new_AGEMA_signal_14241), .Z1_f (new_AGEMA_signal_14242) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1292 ( .A0_t (n710), .A0_f (new_AGEMA_signal_17417), .A1_t (new_AGEMA_signal_17418), .A1_f (new_AGEMA_signal_17419), .B0_t (n709), .B0_f (new_AGEMA_signal_14240), .B1_t (new_AGEMA_signal_14241), .B1_f (new_AGEMA_signal_14242), .Z0_t (RoundOutput[36]), .Z0_f (new_AGEMA_signal_17822), .Z1_t (new_AGEMA_signal_17823), .Z1_f (new_AGEMA_signal_17824) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1293 ( .A0_t (MixColumnsOutput[37]), .A0_f (new_AGEMA_signal_16016), .A1_t (new_AGEMA_signal_16017), .A1_f (new_AGEMA_signal_16018), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n712), .Z0_f (new_AGEMA_signal_16679), .Z1_t (new_AGEMA_signal_16680), .Z1_f (new_AGEMA_signal_16681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1294 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .B0_f (new_AGEMA_signal_13814), .B1_t (new_AGEMA_signal_13815), .B1_f (new_AGEMA_signal_13816), .Z0_t (n711), .Z0_f (new_AGEMA_signal_14243), .Z1_t (new_AGEMA_signal_14244), .Z1_f (new_AGEMA_signal_14245) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1295 ( .A0_t (n712), .A0_f (new_AGEMA_signal_16679), .A1_t (new_AGEMA_signal_16680), .A1_f (new_AGEMA_signal_16681), .B0_t (n711), .B0_f (new_AGEMA_signal_14243), .B1_t (new_AGEMA_signal_14244), .B1_f (new_AGEMA_signal_14245), .Z0_t (RoundOutput[37]), .Z0_f (new_AGEMA_signal_17420), .Z1_t (new_AGEMA_signal_17421), .Z1_f (new_AGEMA_signal_17422) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1296 ( .A0_t (MixColumnsOutput[38]), .A0_f (new_AGEMA_signal_16013), .A1_t (new_AGEMA_signal_16014), .A1_f (new_AGEMA_signal_16015), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n714), .Z0_f (new_AGEMA_signal_16682), .Z1_t (new_AGEMA_signal_16683), .Z1_f (new_AGEMA_signal_16684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1297 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .B0_f (new_AGEMA_signal_13811), .B1_t (new_AGEMA_signal_13812), .B1_f (new_AGEMA_signal_13813), .Z0_t (n713), .Z0_f (new_AGEMA_signal_14246), .Z1_t (new_AGEMA_signal_14247), .Z1_f (new_AGEMA_signal_14248) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1298 ( .A0_t (n714), .A0_f (new_AGEMA_signal_16682), .A1_t (new_AGEMA_signal_16683), .A1_f (new_AGEMA_signal_16684), .B0_t (n713), .B0_f (new_AGEMA_signal_14246), .B1_t (new_AGEMA_signal_14247), .B1_f (new_AGEMA_signal_14248), .Z0_t (RoundOutput[38]), .Z0_f (new_AGEMA_signal_17423), .Z1_t (new_AGEMA_signal_17424), .Z1_f (new_AGEMA_signal_17425) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1299 ( .A0_t (MixColumnsOutput[39]), .A0_f (new_AGEMA_signal_16010), .A1_t (new_AGEMA_signal_16011), .A1_f (new_AGEMA_signal_16012), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n716), .Z0_f (new_AGEMA_signal_16685), .Z1_t (new_AGEMA_signal_16686), .Z1_f (new_AGEMA_signal_16687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1300 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B0_f (new_AGEMA_signal_13808), .B1_t (new_AGEMA_signal_13809), .B1_f (new_AGEMA_signal_13810), .Z0_t (n715), .Z0_f (new_AGEMA_signal_14249), .Z1_t (new_AGEMA_signal_14250), .Z1_f (new_AGEMA_signal_14251) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1301 ( .A0_t (n716), .A0_f (new_AGEMA_signal_16685), .A1_t (new_AGEMA_signal_16686), .A1_f (new_AGEMA_signal_16687), .B0_t (n715), .B0_f (new_AGEMA_signal_14249), .B1_t (new_AGEMA_signal_14250), .B1_f (new_AGEMA_signal_14251), .Z0_t (RoundOutput[39]), .Z0_f (new_AGEMA_signal_17426), .Z1_t (new_AGEMA_signal_17427), .Z1_f (new_AGEMA_signal_17428) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1302 ( .A0_t (MixColumnsOutput[3]), .A0_f (new_AGEMA_signal_16925), .A1_t (new_AGEMA_signal_16926), .A1_f (new_AGEMA_signal_16927), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n718), .Z0_f (new_AGEMA_signal_17429), .Z1_t (new_AGEMA_signal_17430), .Z1_f (new_AGEMA_signal_17431) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1303 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[3]), .B0_f (new_AGEMA_signal_13736), .B1_t (new_AGEMA_signal_13737), .B1_f (new_AGEMA_signal_13738), .Z0_t (n717), .Z0_f (new_AGEMA_signal_14252), .Z1_t (new_AGEMA_signal_14253), .Z1_f (new_AGEMA_signal_14254) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1304 ( .A0_t (n718), .A0_f (new_AGEMA_signal_17429), .A1_t (new_AGEMA_signal_17430), .A1_f (new_AGEMA_signal_17431), .B0_t (n717), .B0_f (new_AGEMA_signal_14252), .B1_t (new_AGEMA_signal_14253), .B1_f (new_AGEMA_signal_14254), .Z0_t (RoundOutput[3]), .Z0_f (new_AGEMA_signal_17825), .Z1_t (new_AGEMA_signal_17826), .Z1_f (new_AGEMA_signal_17827) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1305 ( .A0_t (MixColumnsOutput[40]), .A0_f (new_AGEMA_signal_16007), .A1_t (new_AGEMA_signal_16008), .A1_f (new_AGEMA_signal_16009), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n720), .Z0_f (new_AGEMA_signal_16688), .Z1_t (new_AGEMA_signal_16689), .Z1_f (new_AGEMA_signal_16690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1306 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[40]), .B0_f (new_AGEMA_signal_13427), .B1_t (new_AGEMA_signal_13428), .B1_f (new_AGEMA_signal_13429), .Z0_t (n719), .Z0_f (new_AGEMA_signal_13613), .Z1_t (new_AGEMA_signal_13614), .Z1_f (new_AGEMA_signal_13615) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1307 ( .A0_t (n720), .A0_f (new_AGEMA_signal_16688), .A1_t (new_AGEMA_signal_16689), .A1_f (new_AGEMA_signal_16690), .B0_t (n719), .B0_f (new_AGEMA_signal_13613), .B1_t (new_AGEMA_signal_13614), .B1_f (new_AGEMA_signal_13615), .Z0_t (RoundOutput[40]), .Z0_f (new_AGEMA_signal_17432), .Z1_t (new_AGEMA_signal_17433), .Z1_f (new_AGEMA_signal_17434) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1308 ( .A0_t (MixColumnsOutput[41]), .A0_f (new_AGEMA_signal_16883), .A1_t (new_AGEMA_signal_16884), .A1_f (new_AGEMA_signal_16885), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n722), .Z0_f (new_AGEMA_signal_17435), .Z1_t (new_AGEMA_signal_17436), .Z1_f (new_AGEMA_signal_17437) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1309 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13931), .B1_t (new_AGEMA_signal_13932), .B1_f (new_AGEMA_signal_13933), .Z0_t (n721), .Z0_f (new_AGEMA_signal_14255), .Z1_t (new_AGEMA_signal_14256), .Z1_f (new_AGEMA_signal_14257) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1310 ( .A0_t (n722), .A0_f (new_AGEMA_signal_17435), .A1_t (new_AGEMA_signal_17436), .A1_f (new_AGEMA_signal_17437), .B0_t (n721), .B0_f (new_AGEMA_signal_14255), .B1_t (new_AGEMA_signal_14256), .B1_f (new_AGEMA_signal_14257), .Z0_t (RoundOutput[41]), .Z0_f (new_AGEMA_signal_17828), .Z1_t (new_AGEMA_signal_17829), .Z1_f (new_AGEMA_signal_17830) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1311 ( .A0_t (MixColumnsOutput[42]), .A0_f (new_AGEMA_signal_16094), .A1_t (new_AGEMA_signal_16095), .A1_f (new_AGEMA_signal_16096), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n724), .Z0_f (new_AGEMA_signal_16691), .Z1_t (new_AGEMA_signal_16692), .Z1_f (new_AGEMA_signal_16693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1312 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[42]), .B0_f (new_AGEMA_signal_13928), .B1_t (new_AGEMA_signal_13929), .B1_f (new_AGEMA_signal_13930), .Z0_t (n723), .Z0_f (new_AGEMA_signal_14258), .Z1_t (new_AGEMA_signal_14259), .Z1_f (new_AGEMA_signal_14260) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1313 ( .A0_t (n724), .A0_f (new_AGEMA_signal_16691), .A1_t (new_AGEMA_signal_16692), .A1_f (new_AGEMA_signal_16693), .B0_t (n723), .B0_f (new_AGEMA_signal_14258), .B1_t (new_AGEMA_signal_14259), .B1_f (new_AGEMA_signal_14260), .Z0_t (RoundOutput[42]), .Z0_f (new_AGEMA_signal_17438), .Z1_t (new_AGEMA_signal_17439), .Z1_f (new_AGEMA_signal_17440) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1314 ( .A0_t (MixColumnsOutput[43]), .A0_f (new_AGEMA_signal_16916), .A1_t (new_AGEMA_signal_16917), .A1_f (new_AGEMA_signal_16918), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n726), .Z0_f (new_AGEMA_signal_17441), .Z1_t (new_AGEMA_signal_17442), .Z1_f (new_AGEMA_signal_17443) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1315 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[43]), .B0_f (new_AGEMA_signal_13925), .B1_t (new_AGEMA_signal_13926), .B1_f (new_AGEMA_signal_13927), .Z0_t (n725), .Z0_f (new_AGEMA_signal_14261), .Z1_t (new_AGEMA_signal_14262), .Z1_f (new_AGEMA_signal_14263) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1316 ( .A0_t (n726), .A0_f (new_AGEMA_signal_17441), .A1_t (new_AGEMA_signal_17442), .A1_f (new_AGEMA_signal_17443), .B0_t (n725), .B0_f (new_AGEMA_signal_14261), .B1_t (new_AGEMA_signal_14262), .B1_f (new_AGEMA_signal_14263), .Z0_t (RoundOutput[43]), .Z0_f (new_AGEMA_signal_17831), .Z1_t (new_AGEMA_signal_17832), .Z1_f (new_AGEMA_signal_17833) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1317 ( .A0_t (MixColumnsOutput[44]), .A0_f (new_AGEMA_signal_16913), .A1_t (new_AGEMA_signal_16914), .A1_f (new_AGEMA_signal_16915), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n728), .Z0_f (new_AGEMA_signal_17444), .Z1_t (new_AGEMA_signal_17445), .Z1_f (new_AGEMA_signal_17446) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1318 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13922), .B1_t (new_AGEMA_signal_13923), .B1_f (new_AGEMA_signal_13924), .Z0_t (n727), .Z0_f (new_AGEMA_signal_14264), .Z1_t (new_AGEMA_signal_14265), .Z1_f (new_AGEMA_signal_14266) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1319 ( .A0_t (n728), .A0_f (new_AGEMA_signal_17444), .A1_t (new_AGEMA_signal_17445), .A1_f (new_AGEMA_signal_17446), .B0_t (n727), .B0_f (new_AGEMA_signal_14264), .B1_t (new_AGEMA_signal_14265), .B1_f (new_AGEMA_signal_14266), .Z0_t (RoundOutput[44]), .Z0_f (new_AGEMA_signal_17834), .Z1_t (new_AGEMA_signal_17835), .Z1_f (new_AGEMA_signal_17836) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1320 ( .A0_t (MixColumnsOutput[45]), .A0_f (new_AGEMA_signal_16085), .A1_t (new_AGEMA_signal_16086), .A1_f (new_AGEMA_signal_16087), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n730), .Z0_f (new_AGEMA_signal_16694), .Z1_t (new_AGEMA_signal_16695), .Z1_f (new_AGEMA_signal_16696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1321 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13919), .B1_t (new_AGEMA_signal_13920), .B1_f (new_AGEMA_signal_13921), .Z0_t (n729), .Z0_f (new_AGEMA_signal_14267), .Z1_t (new_AGEMA_signal_14268), .Z1_f (new_AGEMA_signal_14269) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1322 ( .A0_t (n730), .A0_f (new_AGEMA_signal_16694), .A1_t (new_AGEMA_signal_16695), .A1_f (new_AGEMA_signal_16696), .B0_t (n729), .B0_f (new_AGEMA_signal_14267), .B1_t (new_AGEMA_signal_14268), .B1_f (new_AGEMA_signal_14269), .Z0_t (RoundOutput[45]), .Z0_f (new_AGEMA_signal_17447), .Z1_t (new_AGEMA_signal_17448), .Z1_f (new_AGEMA_signal_17449) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1323 ( .A0_t (MixColumnsOutput[46]), .A0_f (new_AGEMA_signal_16082), .A1_t (new_AGEMA_signal_16083), .A1_f (new_AGEMA_signal_16084), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n732), .Z0_f (new_AGEMA_signal_16697), .Z1_t (new_AGEMA_signal_16698), .Z1_f (new_AGEMA_signal_16699) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1324 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13916), .B1_t (new_AGEMA_signal_13917), .B1_f (new_AGEMA_signal_13918), .Z0_t (n731), .Z0_f (new_AGEMA_signal_14270), .Z1_t (new_AGEMA_signal_14271), .Z1_f (new_AGEMA_signal_14272) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1325 ( .A0_t (n732), .A0_f (new_AGEMA_signal_16697), .A1_t (new_AGEMA_signal_16698), .A1_f (new_AGEMA_signal_16699), .B0_t (n731), .B0_f (new_AGEMA_signal_14270), .B1_t (new_AGEMA_signal_14271), .B1_f (new_AGEMA_signal_14272), .Z0_t (RoundOutput[46]), .Z0_f (new_AGEMA_signal_17450), .Z1_t (new_AGEMA_signal_17451), .Z1_f (new_AGEMA_signal_17452) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1326 ( .A0_t (MixColumnsOutput[47]), .A0_f (new_AGEMA_signal_16079), .A1_t (new_AGEMA_signal_16080), .A1_f (new_AGEMA_signal_16081), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n734), .Z0_f (new_AGEMA_signal_16700), .Z1_t (new_AGEMA_signal_16701), .Z1_f (new_AGEMA_signal_16702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1327 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B0_f (new_AGEMA_signal_13913), .B1_t (new_AGEMA_signal_13914), .B1_f (new_AGEMA_signal_13915), .Z0_t (n733), .Z0_f (new_AGEMA_signal_14273), .Z1_t (new_AGEMA_signal_14274), .Z1_f (new_AGEMA_signal_14275) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1328 ( .A0_t (n734), .A0_f (new_AGEMA_signal_16700), .A1_t (new_AGEMA_signal_16701), .A1_f (new_AGEMA_signal_16702), .B0_t (n733), .B0_f (new_AGEMA_signal_14273), .B1_t (new_AGEMA_signal_14274), .B1_f (new_AGEMA_signal_14275), .Z0_t (RoundOutput[47]), .Z0_f (new_AGEMA_signal_17453), .Z1_t (new_AGEMA_signal_17454), .Z1_f (new_AGEMA_signal_17455) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1329 ( .A0_t (MixColumnsOutput[48]), .A0_f (new_AGEMA_signal_16076), .A1_t (new_AGEMA_signal_16077), .A1_f (new_AGEMA_signal_16078), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n736), .Z0_f (new_AGEMA_signal_16703), .Z1_t (new_AGEMA_signal_16704), .Z1_f (new_AGEMA_signal_16705) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1330 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[48]), .B0_f (new_AGEMA_signal_13064), .B1_t (new_AGEMA_signal_13065), .B1_f (new_AGEMA_signal_13066), .Z0_t (n735), .Z0_f (new_AGEMA_signal_13616), .Z1_t (new_AGEMA_signal_13617), .Z1_f (new_AGEMA_signal_13618) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1331 ( .A0_t (n736), .A0_f (new_AGEMA_signal_16703), .A1_t (new_AGEMA_signal_16704), .A1_f (new_AGEMA_signal_16705), .B0_t (n735), .B0_f (new_AGEMA_signal_13616), .B1_t (new_AGEMA_signal_13617), .B1_f (new_AGEMA_signal_13618), .Z0_t (RoundOutput[48]), .Z0_f (new_AGEMA_signal_17456), .Z1_t (new_AGEMA_signal_17457), .Z1_f (new_AGEMA_signal_17458) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1332 ( .A0_t (MixColumnsOutput[49]), .A0_f (new_AGEMA_signal_16910), .A1_t (new_AGEMA_signal_16911), .A1_f (new_AGEMA_signal_16912), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n738), .Z0_f (new_AGEMA_signal_17459), .Z1_t (new_AGEMA_signal_17460), .Z1_f (new_AGEMA_signal_17461) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1333 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13700), .B1_t (new_AGEMA_signal_13701), .B1_f (new_AGEMA_signal_13702), .Z0_t (n737), .Z0_f (new_AGEMA_signal_14276), .Z1_t (new_AGEMA_signal_14277), .Z1_f (new_AGEMA_signal_14278) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1334 ( .A0_t (n738), .A0_f (new_AGEMA_signal_17459), .A1_t (new_AGEMA_signal_17460), .A1_f (new_AGEMA_signal_17461), .B0_t (n737), .B0_f (new_AGEMA_signal_14276), .B1_t (new_AGEMA_signal_14277), .B1_f (new_AGEMA_signal_14278), .Z0_t (RoundOutput[49]), .Z0_f (new_AGEMA_signal_17837), .Z1_t (new_AGEMA_signal_17838), .Z1_f (new_AGEMA_signal_17839) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1335 ( .A0_t (MixColumnsOutput[4]), .A0_f (new_AGEMA_signal_16922), .A1_t (new_AGEMA_signal_16923), .A1_f (new_AGEMA_signal_16924), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n740), .Z0_f (new_AGEMA_signal_17462), .Z1_t (new_AGEMA_signal_17463), .Z1_f (new_AGEMA_signal_17464) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1336 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .B0_f (new_AGEMA_signal_13733), .B1_t (new_AGEMA_signal_13734), .B1_f (new_AGEMA_signal_13735), .Z0_t (n739), .Z0_f (new_AGEMA_signal_14279), .Z1_t (new_AGEMA_signal_14280), .Z1_f (new_AGEMA_signal_14281) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1337 ( .A0_t (n740), .A0_f (new_AGEMA_signal_17462), .A1_t (new_AGEMA_signal_17463), .A1_f (new_AGEMA_signal_17464), .B0_t (n739), .B0_f (new_AGEMA_signal_14279), .B1_t (new_AGEMA_signal_14280), .B1_f (new_AGEMA_signal_14281), .Z0_t (RoundOutput[4]), .Z0_f (new_AGEMA_signal_17840), .Z1_t (new_AGEMA_signal_17841), .Z1_f (new_AGEMA_signal_17842) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1338 ( .A0_t (MixColumnsOutput[50]), .A0_f (new_AGEMA_signal_16070), .A1_t (new_AGEMA_signal_16071), .A1_f (new_AGEMA_signal_16072), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n742), .Z0_f (new_AGEMA_signal_16706), .Z1_t (new_AGEMA_signal_16707), .Z1_f (new_AGEMA_signal_16708) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1339 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[50]), .B0_f (new_AGEMA_signal_13697), .B1_t (new_AGEMA_signal_13698), .B1_f (new_AGEMA_signal_13699), .Z0_t (n741), .Z0_f (new_AGEMA_signal_14282), .Z1_t (new_AGEMA_signal_14283), .Z1_f (new_AGEMA_signal_14284) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1340 ( .A0_t (n742), .A0_f (new_AGEMA_signal_16706), .A1_t (new_AGEMA_signal_16707), .A1_f (new_AGEMA_signal_16708), .B0_t (n741), .B0_f (new_AGEMA_signal_14282), .B1_t (new_AGEMA_signal_14283), .B1_f (new_AGEMA_signal_14284), .Z0_t (RoundOutput[50]), .Z0_f (new_AGEMA_signal_17465), .Z1_t (new_AGEMA_signal_17466), .Z1_f (new_AGEMA_signal_17467) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1341 ( .A0_t (MixColumnsOutput[51]), .A0_f (new_AGEMA_signal_16907), .A1_t (new_AGEMA_signal_16908), .A1_f (new_AGEMA_signal_16909), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n744), .Z0_f (new_AGEMA_signal_17468), .Z1_t (new_AGEMA_signal_17469), .Z1_f (new_AGEMA_signal_17470) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1342 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[51]), .B0_f (new_AGEMA_signal_13694), .B1_t (new_AGEMA_signal_13695), .B1_f (new_AGEMA_signal_13696), .Z0_t (n743), .Z0_f (new_AGEMA_signal_14285), .Z1_t (new_AGEMA_signal_14286), .Z1_f (new_AGEMA_signal_14287) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1343 ( .A0_t (n744), .A0_f (new_AGEMA_signal_17468), .A1_t (new_AGEMA_signal_17469), .A1_f (new_AGEMA_signal_17470), .B0_t (n743), .B0_f (new_AGEMA_signal_14285), .B1_t (new_AGEMA_signal_14286), .B1_f (new_AGEMA_signal_14287), .Z0_t (RoundOutput[51]), .Z0_f (new_AGEMA_signal_17843), .Z1_t (new_AGEMA_signal_17844), .Z1_f (new_AGEMA_signal_17845) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1344 ( .A0_t (MixColumnsOutput[52]), .A0_f (new_AGEMA_signal_16901), .A1_t (new_AGEMA_signal_16902), .A1_f (new_AGEMA_signal_16903), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n746), .Z0_f (new_AGEMA_signal_17471), .Z1_t (new_AGEMA_signal_17472), .Z1_f (new_AGEMA_signal_17473) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1345 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13691), .B1_t (new_AGEMA_signal_13692), .B1_f (new_AGEMA_signal_13693), .Z0_t (n745), .Z0_f (new_AGEMA_signal_14288), .Z1_t (new_AGEMA_signal_14289), .Z1_f (new_AGEMA_signal_14290) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1346 ( .A0_t (n746), .A0_f (new_AGEMA_signal_17471), .A1_t (new_AGEMA_signal_17472), .A1_f (new_AGEMA_signal_17473), .B0_t (n745), .B0_f (new_AGEMA_signal_14288), .B1_t (new_AGEMA_signal_14289), .B1_f (new_AGEMA_signal_14290), .Z0_t (RoundOutput[52]), .Z0_f (new_AGEMA_signal_17846), .Z1_t (new_AGEMA_signal_17847), .Z1_f (new_AGEMA_signal_17848) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1347 ( .A0_t (MixColumnsOutput[53]), .A0_f (new_AGEMA_signal_16058), .A1_t (new_AGEMA_signal_16059), .A1_f (new_AGEMA_signal_16060), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n748), .Z0_f (new_AGEMA_signal_16709), .Z1_t (new_AGEMA_signal_16710), .Z1_f (new_AGEMA_signal_16711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1348 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13688), .B1_t (new_AGEMA_signal_13689), .B1_f (new_AGEMA_signal_13690), .Z0_t (n747), .Z0_f (new_AGEMA_signal_14291), .Z1_t (new_AGEMA_signal_14292), .Z1_f (new_AGEMA_signal_14293) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1349 ( .A0_t (n748), .A0_f (new_AGEMA_signal_16709), .A1_t (new_AGEMA_signal_16710), .A1_f (new_AGEMA_signal_16711), .B0_t (n747), .B0_f (new_AGEMA_signal_14291), .B1_t (new_AGEMA_signal_14292), .B1_f (new_AGEMA_signal_14293), .Z0_t (RoundOutput[53]), .Z0_f (new_AGEMA_signal_17474), .Z1_t (new_AGEMA_signal_17475), .Z1_f (new_AGEMA_signal_17476) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1350 ( .A0_t (MixColumnsOutput[54]), .A0_f (new_AGEMA_signal_16055), .A1_t (new_AGEMA_signal_16056), .A1_f (new_AGEMA_signal_16057), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n750), .Z0_f (new_AGEMA_signal_16712), .Z1_t (new_AGEMA_signal_16713), .Z1_f (new_AGEMA_signal_16714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1351 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13685), .B1_t (new_AGEMA_signal_13686), .B1_f (new_AGEMA_signal_13687), .Z0_t (n749), .Z0_f (new_AGEMA_signal_14294), .Z1_t (new_AGEMA_signal_14295), .Z1_f (new_AGEMA_signal_14296) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1352 ( .A0_t (n750), .A0_f (new_AGEMA_signal_16712), .A1_t (new_AGEMA_signal_16713), .A1_f (new_AGEMA_signal_16714), .B0_t (n749), .B0_f (new_AGEMA_signal_14294), .B1_t (new_AGEMA_signal_14295), .B1_f (new_AGEMA_signal_14296), .Z0_t (RoundOutput[54]), .Z0_f (new_AGEMA_signal_17477), .Z1_t (new_AGEMA_signal_17478), .Z1_f (new_AGEMA_signal_17479) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1353 ( .A0_t (MixColumnsOutput[55]), .A0_f (new_AGEMA_signal_16052), .A1_t (new_AGEMA_signal_16053), .A1_f (new_AGEMA_signal_16054), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n752), .Z0_f (new_AGEMA_signal_16715), .Z1_t (new_AGEMA_signal_16716), .Z1_f (new_AGEMA_signal_16717) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1354 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13682), .B1_t (new_AGEMA_signal_13683), .B1_f (new_AGEMA_signal_13684), .Z0_t (n751), .Z0_f (new_AGEMA_signal_14297), .Z1_t (new_AGEMA_signal_14298), .Z1_f (new_AGEMA_signal_14299) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1355 ( .A0_t (n752), .A0_f (new_AGEMA_signal_16715), .A1_t (new_AGEMA_signal_16716), .A1_f (new_AGEMA_signal_16717), .B0_t (n751), .B0_f (new_AGEMA_signal_14297), .B1_t (new_AGEMA_signal_14298), .B1_f (new_AGEMA_signal_14299), .Z0_t (RoundOutput[55]), .Z0_f (new_AGEMA_signal_17480), .Z1_t (new_AGEMA_signal_17481), .Z1_f (new_AGEMA_signal_17482) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1356 ( .A0_t (MixColumnsOutput[56]), .A0_f (new_AGEMA_signal_16049), .A1_t (new_AGEMA_signal_16050), .A1_f (new_AGEMA_signal_16051), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n754), .Z0_f (new_AGEMA_signal_16718), .Z1_t (new_AGEMA_signal_16719), .Z1_f (new_AGEMA_signal_16720) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1357 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[56]), .B0_f (new_AGEMA_signal_13229), .B1_t (new_AGEMA_signal_13230), .B1_f (new_AGEMA_signal_13231), .Z0_t (n753), .Z0_f (new_AGEMA_signal_13619), .Z1_t (new_AGEMA_signal_13620), .Z1_f (new_AGEMA_signal_13621) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1358 ( .A0_t (n754), .A0_f (new_AGEMA_signal_16718), .A1_t (new_AGEMA_signal_16719), .A1_f (new_AGEMA_signal_16720), .B0_t (n753), .B0_f (new_AGEMA_signal_13619), .B1_t (new_AGEMA_signal_13620), .B1_f (new_AGEMA_signal_13621), .Z0_t (RoundOutput[56]), .Z0_f (new_AGEMA_signal_17483), .Z1_t (new_AGEMA_signal_17484), .Z1_f (new_AGEMA_signal_17485) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1359 ( .A0_t (MixColumnsOutput[57]), .A0_f (new_AGEMA_signal_16898), .A1_t (new_AGEMA_signal_16899), .A1_f (new_AGEMA_signal_16900), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n756), .Z0_f (new_AGEMA_signal_17486), .Z1_t (new_AGEMA_signal_17487), .Z1_f (new_AGEMA_signal_17488) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1360 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13805), .B1_t (new_AGEMA_signal_13806), .B1_f (new_AGEMA_signal_13807), .Z0_t (n755), .Z0_f (new_AGEMA_signal_14300), .Z1_t (new_AGEMA_signal_14301), .Z1_f (new_AGEMA_signal_14302) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1361 ( .A0_t (n756), .A0_f (new_AGEMA_signal_17486), .A1_t (new_AGEMA_signal_17487), .A1_f (new_AGEMA_signal_17488), .B0_t (n755), .B0_f (new_AGEMA_signal_14300), .B1_t (new_AGEMA_signal_14301), .B1_f (new_AGEMA_signal_14302), .Z0_t (RoundOutput[57]), .Z0_f (new_AGEMA_signal_17849), .Z1_t (new_AGEMA_signal_17850), .Z1_f (new_AGEMA_signal_17851) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1362 ( .A0_t (MixColumnsOutput[58]), .A0_f (new_AGEMA_signal_16043), .A1_t (new_AGEMA_signal_16044), .A1_f (new_AGEMA_signal_16045), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n758), .Z0_f (new_AGEMA_signal_16721), .Z1_t (new_AGEMA_signal_16722), .Z1_f (new_AGEMA_signal_16723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1363 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[58]), .B0_f (new_AGEMA_signal_13802), .B1_t (new_AGEMA_signal_13803), .B1_f (new_AGEMA_signal_13804), .Z0_t (n757), .Z0_f (new_AGEMA_signal_14303), .Z1_t (new_AGEMA_signal_14304), .Z1_f (new_AGEMA_signal_14305) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1364 ( .A0_t (n758), .A0_f (new_AGEMA_signal_16721), .A1_t (new_AGEMA_signal_16722), .A1_f (new_AGEMA_signal_16723), .B0_t (n757), .B0_f (new_AGEMA_signal_14303), .B1_t (new_AGEMA_signal_14304), .B1_f (new_AGEMA_signal_14305), .Z0_t (RoundOutput[58]), .Z0_f (new_AGEMA_signal_17489), .Z1_t (new_AGEMA_signal_17490), .Z1_f (new_AGEMA_signal_17491) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1365 ( .A0_t (MixColumnsOutput[59]), .A0_f (new_AGEMA_signal_16895), .A1_t (new_AGEMA_signal_16896), .A1_f (new_AGEMA_signal_16897), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n760), .Z0_f (new_AGEMA_signal_17492), .Z1_t (new_AGEMA_signal_17493), .Z1_f (new_AGEMA_signal_17494) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1366 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[59]), .B0_f (new_AGEMA_signal_13799), .B1_t (new_AGEMA_signal_13800), .B1_f (new_AGEMA_signal_13801), .Z0_t (n759), .Z0_f (new_AGEMA_signal_14306), .Z1_t (new_AGEMA_signal_14307), .Z1_f (new_AGEMA_signal_14308) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1367 ( .A0_t (n760), .A0_f (new_AGEMA_signal_17492), .A1_t (new_AGEMA_signal_17493), .A1_f (new_AGEMA_signal_17494), .B0_t (n759), .B0_f (new_AGEMA_signal_14306), .B1_t (new_AGEMA_signal_14307), .B1_f (new_AGEMA_signal_14308), .Z0_t (RoundOutput[59]), .Z0_f (new_AGEMA_signal_17852), .Z1_t (new_AGEMA_signal_17853), .Z1_f (new_AGEMA_signal_17854) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1368 ( .A0_t (MixColumnsOutput[5]), .A0_f (new_AGEMA_signal_16112), .A1_t (new_AGEMA_signal_16113), .A1_f (new_AGEMA_signal_16114), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n762), .Z0_f (new_AGEMA_signal_16724), .Z1_t (new_AGEMA_signal_16725), .Z1_f (new_AGEMA_signal_16726) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1369 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .B0_f (new_AGEMA_signal_13730), .B1_t (new_AGEMA_signal_13731), .B1_f (new_AGEMA_signal_13732), .Z0_t (n761), .Z0_f (new_AGEMA_signal_14309), .Z1_t (new_AGEMA_signal_14310), .Z1_f (new_AGEMA_signal_14311) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1370 ( .A0_t (n762), .A0_f (new_AGEMA_signal_16724), .A1_t (new_AGEMA_signal_16725), .A1_f (new_AGEMA_signal_16726), .B0_t (n761), .B0_f (new_AGEMA_signal_14309), .B1_t (new_AGEMA_signal_14310), .B1_f (new_AGEMA_signal_14311), .Z0_t (RoundOutput[5]), .Z0_f (new_AGEMA_signal_17495), .Z1_t (new_AGEMA_signal_17496), .Z1_f (new_AGEMA_signal_17497) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1371 ( .A0_t (MixColumnsOutput[60]), .A0_f (new_AGEMA_signal_16892), .A1_t (new_AGEMA_signal_16893), .A1_f (new_AGEMA_signal_16894), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n764), .Z0_f (new_AGEMA_signal_17498), .Z1_t (new_AGEMA_signal_17499), .Z1_f (new_AGEMA_signal_17500) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1372 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13796), .B1_t (new_AGEMA_signal_13797), .B1_f (new_AGEMA_signal_13798), .Z0_t (n763), .Z0_f (new_AGEMA_signal_14312), .Z1_t (new_AGEMA_signal_14313), .Z1_f (new_AGEMA_signal_14314) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1373 ( .A0_t (n764), .A0_f (new_AGEMA_signal_17498), .A1_t (new_AGEMA_signal_17499), .A1_f (new_AGEMA_signal_17500), .B0_t (n763), .B0_f (new_AGEMA_signal_14312), .B1_t (new_AGEMA_signal_14313), .B1_f (new_AGEMA_signal_14314), .Z0_t (RoundOutput[60]), .Z0_f (new_AGEMA_signal_17855), .Z1_t (new_AGEMA_signal_17856), .Z1_f (new_AGEMA_signal_17857) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1374 ( .A0_t (MixColumnsOutput[61]), .A0_f (new_AGEMA_signal_16034), .A1_t (new_AGEMA_signal_16035), .A1_f (new_AGEMA_signal_16036), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n766), .Z0_f (new_AGEMA_signal_16727), .Z1_t (new_AGEMA_signal_16728), .Z1_f (new_AGEMA_signal_16729) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1375 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13793), .B1_t (new_AGEMA_signal_13794), .B1_f (new_AGEMA_signal_13795), .Z0_t (n765), .Z0_f (new_AGEMA_signal_14315), .Z1_t (new_AGEMA_signal_14316), .Z1_f (new_AGEMA_signal_14317) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1376 ( .A0_t (n766), .A0_f (new_AGEMA_signal_16727), .A1_t (new_AGEMA_signal_16728), .A1_f (new_AGEMA_signal_16729), .B0_t (n765), .B0_f (new_AGEMA_signal_14315), .B1_t (new_AGEMA_signal_14316), .B1_f (new_AGEMA_signal_14317), .Z0_t (RoundOutput[61]), .Z0_f (new_AGEMA_signal_17501), .Z1_t (new_AGEMA_signal_17502), .Z1_f (new_AGEMA_signal_17503) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1377 ( .A0_t (MixColumnsOutput[62]), .A0_f (new_AGEMA_signal_16028), .A1_t (new_AGEMA_signal_16029), .A1_f (new_AGEMA_signal_16030), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n768), .Z0_f (new_AGEMA_signal_16730), .Z1_t (new_AGEMA_signal_16731), .Z1_f (new_AGEMA_signal_16732) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1378 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13790), .B1_t (new_AGEMA_signal_13791), .B1_f (new_AGEMA_signal_13792), .Z0_t (n767), .Z0_f (new_AGEMA_signal_14318), .Z1_t (new_AGEMA_signal_14319), .Z1_f (new_AGEMA_signal_14320) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1379 ( .A0_t (n768), .A0_f (new_AGEMA_signal_16730), .A1_t (new_AGEMA_signal_16731), .A1_f (new_AGEMA_signal_16732), .B0_t (n767), .B0_f (new_AGEMA_signal_14318), .B1_t (new_AGEMA_signal_14319), .B1_f (new_AGEMA_signal_14320), .Z0_t (RoundOutput[62]), .Z0_f (new_AGEMA_signal_17504), .Z1_t (new_AGEMA_signal_17505), .Z1_f (new_AGEMA_signal_17506) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1380 ( .A0_t (MixColumnsOutput[63]), .A0_f (new_AGEMA_signal_16025), .A1_t (new_AGEMA_signal_16026), .A1_f (new_AGEMA_signal_16027), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n770), .Z0_f (new_AGEMA_signal_16733), .Z1_t (new_AGEMA_signal_16734), .Z1_f (new_AGEMA_signal_16735) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1381 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13787), .B1_t (new_AGEMA_signal_13788), .B1_f (new_AGEMA_signal_13789), .Z0_t (n769), .Z0_f (new_AGEMA_signal_14321), .Z1_t (new_AGEMA_signal_14322), .Z1_f (new_AGEMA_signal_14323) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1382 ( .A0_t (n770), .A0_f (new_AGEMA_signal_16733), .A1_t (new_AGEMA_signal_16734), .A1_f (new_AGEMA_signal_16735), .B0_t (n769), .B0_f (new_AGEMA_signal_14321), .B1_t (new_AGEMA_signal_14322), .B1_f (new_AGEMA_signal_14323), .Z0_t (RoundOutput[63]), .Z0_f (new_AGEMA_signal_17507), .Z1_t (new_AGEMA_signal_17508), .Z1_f (new_AGEMA_signal_17509) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1383 ( .A0_t (MixColumnsOutput[64]), .A0_f (new_AGEMA_signal_16001), .A1_t (new_AGEMA_signal_16002), .A1_f (new_AGEMA_signal_16003), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n772), .Z0_f (new_AGEMA_signal_16736), .Z1_t (new_AGEMA_signal_16737), .Z1_f (new_AGEMA_signal_16738) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1384 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[64]), .B0_f (new_AGEMA_signal_13394), .B1_t (new_AGEMA_signal_13395), .B1_f (new_AGEMA_signal_13396), .Z0_t (n771), .Z0_f (new_AGEMA_signal_13622), .Z1_t (new_AGEMA_signal_13623), .Z1_f (new_AGEMA_signal_13624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1385 ( .A0_t (n772), .A0_f (new_AGEMA_signal_16736), .A1_t (new_AGEMA_signal_16737), .A1_f (new_AGEMA_signal_16738), .B0_t (n771), .B0_f (new_AGEMA_signal_13622), .B1_t (new_AGEMA_signal_13623), .B1_f (new_AGEMA_signal_13624), .Z0_t (RoundOutput[64]), .Z0_f (new_AGEMA_signal_17510), .Z1_t (new_AGEMA_signal_17511), .Z1_f (new_AGEMA_signal_17512) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1386 ( .A0_t (MixColumnsOutput[65]), .A0_f (new_AGEMA_signal_16868), .A1_t (new_AGEMA_signal_16869), .A1_f (new_AGEMA_signal_16870), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n774), .Z0_f (new_AGEMA_signal_17513), .Z1_t (new_AGEMA_signal_17514), .Z1_f (new_AGEMA_signal_17515) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1387 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .B0_f (new_AGEMA_signal_13910), .B1_t (new_AGEMA_signal_13911), .B1_f (new_AGEMA_signal_13912), .Z0_t (n773), .Z0_f (new_AGEMA_signal_14324), .Z1_t (new_AGEMA_signal_14325), .Z1_f (new_AGEMA_signal_14326) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1388 ( .A0_t (n774), .A0_f (new_AGEMA_signal_17513), .A1_t (new_AGEMA_signal_17514), .A1_f (new_AGEMA_signal_17515), .B0_t (n773), .B0_f (new_AGEMA_signal_14324), .B1_t (new_AGEMA_signal_14325), .B1_f (new_AGEMA_signal_14326), .Z0_t (RoundOutput[65]), .Z0_f (new_AGEMA_signal_17858), .Z1_t (new_AGEMA_signal_17859), .Z1_f (new_AGEMA_signal_17860) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1389 ( .A0_t (MixColumnsOutput[66]), .A0_f (new_AGEMA_signal_15935), .A1_t (new_AGEMA_signal_15936), .A1_f (new_AGEMA_signal_15937), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n776), .Z0_f (new_AGEMA_signal_16739), .Z1_t (new_AGEMA_signal_16740), .Z1_f (new_AGEMA_signal_16741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1390 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[66]), .B0_f (new_AGEMA_signal_13907), .B1_t (new_AGEMA_signal_13908), .B1_f (new_AGEMA_signal_13909), .Z0_t (n775), .Z0_f (new_AGEMA_signal_14327), .Z1_t (new_AGEMA_signal_14328), .Z1_f (new_AGEMA_signal_14329) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1391 ( .A0_t (n776), .A0_f (new_AGEMA_signal_16739), .A1_t (new_AGEMA_signal_16740), .A1_f (new_AGEMA_signal_16741), .B0_t (n775), .B0_f (new_AGEMA_signal_14327), .B1_t (new_AGEMA_signal_14328), .B1_f (new_AGEMA_signal_14329), .Z0_t (RoundOutput[66]), .Z0_f (new_AGEMA_signal_17516), .Z1_t (new_AGEMA_signal_17517), .Z1_f (new_AGEMA_signal_17518) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1392 ( .A0_t (MixColumnsOutput[67]), .A0_f (new_AGEMA_signal_16853), .A1_t (new_AGEMA_signal_16854), .A1_f (new_AGEMA_signal_16855), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n778), .Z0_f (new_AGEMA_signal_17519), .Z1_t (new_AGEMA_signal_17520), .Z1_f (new_AGEMA_signal_17521) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1393 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[67]), .B0_f (new_AGEMA_signal_13904), .B1_t (new_AGEMA_signal_13905), .B1_f (new_AGEMA_signal_13906), .Z0_t (n777), .Z0_f (new_AGEMA_signal_14330), .Z1_t (new_AGEMA_signal_14331), .Z1_f (new_AGEMA_signal_14332) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1394 ( .A0_t (n778), .A0_f (new_AGEMA_signal_17519), .A1_t (new_AGEMA_signal_17520), .A1_f (new_AGEMA_signal_17521), .B0_t (n777), .B0_f (new_AGEMA_signal_14330), .B1_t (new_AGEMA_signal_14331), .B1_f (new_AGEMA_signal_14332), .Z0_t (RoundOutput[67]), .Z0_f (new_AGEMA_signal_17861), .Z1_t (new_AGEMA_signal_17862), .Z1_f (new_AGEMA_signal_17863) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1395 ( .A0_t (MixColumnsOutput[68]), .A0_f (new_AGEMA_signal_16850), .A1_t (new_AGEMA_signal_16851), .A1_f (new_AGEMA_signal_16852), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n780), .Z0_f (new_AGEMA_signal_17522), .Z1_t (new_AGEMA_signal_17523), .Z1_f (new_AGEMA_signal_17524) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1396 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .B0_f (new_AGEMA_signal_13901), .B1_t (new_AGEMA_signal_13902), .B1_f (new_AGEMA_signal_13903), .Z0_t (n779), .Z0_f (new_AGEMA_signal_14333), .Z1_t (new_AGEMA_signal_14334), .Z1_f (new_AGEMA_signal_14335) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1397 ( .A0_t (n780), .A0_f (new_AGEMA_signal_17522), .A1_t (new_AGEMA_signal_17523), .A1_f (new_AGEMA_signal_17524), .B0_t (n779), .B0_f (new_AGEMA_signal_14333), .B1_t (new_AGEMA_signal_14334), .B1_f (new_AGEMA_signal_14335), .Z0_t (RoundOutput[68]), .Z0_f (new_AGEMA_signal_17864), .Z1_t (new_AGEMA_signal_17865), .Z1_f (new_AGEMA_signal_17866) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1398 ( .A0_t (MixColumnsOutput[69]), .A0_f (new_AGEMA_signal_15920), .A1_t (new_AGEMA_signal_15921), .A1_f (new_AGEMA_signal_15922), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n782), .Z0_f (new_AGEMA_signal_16742), .Z1_t (new_AGEMA_signal_16743), .Z1_f (new_AGEMA_signal_16744) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1399 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .B0_f (new_AGEMA_signal_13898), .B1_t (new_AGEMA_signal_13899), .B1_f (new_AGEMA_signal_13900), .Z0_t (n781), .Z0_f (new_AGEMA_signal_14336), .Z1_t (new_AGEMA_signal_14337), .Z1_f (new_AGEMA_signal_14338) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1400 ( .A0_t (n782), .A0_f (new_AGEMA_signal_16742), .A1_t (new_AGEMA_signal_16743), .A1_f (new_AGEMA_signal_16744), .B0_t (n781), .B0_f (new_AGEMA_signal_14336), .B1_t (new_AGEMA_signal_14337), .B1_f (new_AGEMA_signal_14338), .Z0_t (RoundOutput[69]), .Z0_f (new_AGEMA_signal_17525), .Z1_t (new_AGEMA_signal_17526), .Z1_f (new_AGEMA_signal_17527) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1401 ( .A0_t (MixColumnsOutput[6]), .A0_f (new_AGEMA_signal_16109), .A1_t (new_AGEMA_signal_16110), .A1_f (new_AGEMA_signal_16111), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n784), .Z0_f (new_AGEMA_signal_16745), .Z1_t (new_AGEMA_signal_16746), .Z1_f (new_AGEMA_signal_16747) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1402 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .B0_f (new_AGEMA_signal_13727), .B1_t (new_AGEMA_signal_13728), .B1_f (new_AGEMA_signal_13729), .Z0_t (n783), .Z0_f (new_AGEMA_signal_14339), .Z1_t (new_AGEMA_signal_14340), .Z1_f (new_AGEMA_signal_14341) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1403 ( .A0_t (n784), .A0_f (new_AGEMA_signal_16745), .A1_t (new_AGEMA_signal_16746), .A1_f (new_AGEMA_signal_16747), .B0_t (n783), .B0_f (new_AGEMA_signal_14339), .B1_t (new_AGEMA_signal_14340), .B1_f (new_AGEMA_signal_14341), .Z0_t (RoundOutput[6]), .Z0_f (new_AGEMA_signal_17528), .Z1_t (new_AGEMA_signal_17529), .Z1_f (new_AGEMA_signal_17530) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1404 ( .A0_t (MixColumnsOutput[70]), .A0_f (new_AGEMA_signal_15917), .A1_t (new_AGEMA_signal_15918), .A1_f (new_AGEMA_signal_15919), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n786), .Z0_f (new_AGEMA_signal_16748), .Z1_t (new_AGEMA_signal_16749), .Z1_f (new_AGEMA_signal_16750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1405 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .B0_f (new_AGEMA_signal_13895), .B1_t (new_AGEMA_signal_13896), .B1_f (new_AGEMA_signal_13897), .Z0_t (n785), .Z0_f (new_AGEMA_signal_14342), .Z1_t (new_AGEMA_signal_14343), .Z1_f (new_AGEMA_signal_14344) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1406 ( .A0_t (n786), .A0_f (new_AGEMA_signal_16748), .A1_t (new_AGEMA_signal_16749), .A1_f (new_AGEMA_signal_16750), .B0_t (n785), .B0_f (new_AGEMA_signal_14342), .B1_t (new_AGEMA_signal_14343), .B1_f (new_AGEMA_signal_14344), .Z0_t (RoundOutput[70]), .Z0_f (new_AGEMA_signal_17531), .Z1_t (new_AGEMA_signal_17532), .Z1_f (new_AGEMA_signal_17533) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1407 ( .A0_t (MixColumnsOutput[71]), .A0_f (new_AGEMA_signal_15914), .A1_t (new_AGEMA_signal_15915), .A1_f (new_AGEMA_signal_15916), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n788), .Z0_f (new_AGEMA_signal_16751), .Z1_t (new_AGEMA_signal_16752), .Z1_f (new_AGEMA_signal_16753) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1408 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B0_f (new_AGEMA_signal_13892), .B1_t (new_AGEMA_signal_13893), .B1_f (new_AGEMA_signal_13894), .Z0_t (n787), .Z0_f (new_AGEMA_signal_14345), .Z1_t (new_AGEMA_signal_14346), .Z1_f (new_AGEMA_signal_14347) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1409 ( .A0_t (n788), .A0_f (new_AGEMA_signal_16751), .A1_t (new_AGEMA_signal_16752), .A1_f (new_AGEMA_signal_16753), .B0_t (n787), .B0_f (new_AGEMA_signal_14345), .B1_t (new_AGEMA_signal_14346), .B1_f (new_AGEMA_signal_14347), .Z0_t (RoundOutput[71]), .Z0_f (new_AGEMA_signal_17534), .Z1_t (new_AGEMA_signal_17535), .Z1_f (new_AGEMA_signal_17536) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1410 ( .A0_t (MixColumnsOutput[72]), .A0_f (new_AGEMA_signal_15911), .A1_t (new_AGEMA_signal_15912), .A1_f (new_AGEMA_signal_15913), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n790), .Z0_f (new_AGEMA_signal_16754), .Z1_t (new_AGEMA_signal_16755), .Z1_f (new_AGEMA_signal_16756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1411 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[72]), .B0_f (new_AGEMA_signal_13031), .B1_t (new_AGEMA_signal_13032), .B1_f (new_AGEMA_signal_13033), .Z0_t (n789), .Z0_f (new_AGEMA_signal_13625), .Z1_t (new_AGEMA_signal_13626), .Z1_f (new_AGEMA_signal_13627) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1412 ( .A0_t (n790), .A0_f (new_AGEMA_signal_16754), .A1_t (new_AGEMA_signal_16755), .A1_f (new_AGEMA_signal_16756), .B0_t (n789), .B0_f (new_AGEMA_signal_13625), .B1_t (new_AGEMA_signal_13626), .B1_f (new_AGEMA_signal_13627), .Z0_t (RoundOutput[72]), .Z0_f (new_AGEMA_signal_17537), .Z1_t (new_AGEMA_signal_17538), .Z1_f (new_AGEMA_signal_17539) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1413 ( .A0_t (MixColumnsOutput[73]), .A0_f (new_AGEMA_signal_16847), .A1_t (new_AGEMA_signal_16848), .A1_f (new_AGEMA_signal_16849), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n792), .Z0_f (new_AGEMA_signal_17540), .Z1_t (new_AGEMA_signal_17541), .Z1_f (new_AGEMA_signal_17542) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1414 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13679), .B1_t (new_AGEMA_signal_13680), .B1_f (new_AGEMA_signal_13681), .Z0_t (n791), .Z0_f (new_AGEMA_signal_14348), .Z1_t (new_AGEMA_signal_14349), .Z1_f (new_AGEMA_signal_14350) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1415 ( .A0_t (n792), .A0_f (new_AGEMA_signal_17540), .A1_t (new_AGEMA_signal_17541), .A1_f (new_AGEMA_signal_17542), .B0_t (n791), .B0_f (new_AGEMA_signal_14348), .B1_t (new_AGEMA_signal_14349), .B1_f (new_AGEMA_signal_14350), .Z0_t (RoundOutput[73]), .Z0_f (new_AGEMA_signal_17867), .Z1_t (new_AGEMA_signal_17868), .Z1_f (new_AGEMA_signal_17869) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1416 ( .A0_t (MixColumnsOutput[74]), .A0_f (new_AGEMA_signal_15998), .A1_t (new_AGEMA_signal_15999), .A1_f (new_AGEMA_signal_16000), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n794), .Z0_f (new_AGEMA_signal_16757), .Z1_t (new_AGEMA_signal_16758), .Z1_f (new_AGEMA_signal_16759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1417 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[74]), .B0_f (new_AGEMA_signal_13676), .B1_t (new_AGEMA_signal_13677), .B1_f (new_AGEMA_signal_13678), .Z0_t (n793), .Z0_f (new_AGEMA_signal_14351), .Z1_t (new_AGEMA_signal_14352), .Z1_f (new_AGEMA_signal_14353) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1418 ( .A0_t (n794), .A0_f (new_AGEMA_signal_16757), .A1_t (new_AGEMA_signal_16758), .A1_f (new_AGEMA_signal_16759), .B0_t (n793), .B0_f (new_AGEMA_signal_14351), .B1_t (new_AGEMA_signal_14352), .B1_f (new_AGEMA_signal_14353), .Z0_t (RoundOutput[74]), .Z0_f (new_AGEMA_signal_17543), .Z1_t (new_AGEMA_signal_17544), .Z1_f (new_AGEMA_signal_17545) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1419 ( .A0_t (MixColumnsOutput[75]), .A0_f (new_AGEMA_signal_16880), .A1_t (new_AGEMA_signal_16881), .A1_f (new_AGEMA_signal_16882), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n796), .Z0_f (new_AGEMA_signal_17546), .Z1_t (new_AGEMA_signal_17547), .Z1_f (new_AGEMA_signal_17548) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1420 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[75]), .B0_f (new_AGEMA_signal_13673), .B1_t (new_AGEMA_signal_13674), .B1_f (new_AGEMA_signal_13675), .Z0_t (n795), .Z0_f (new_AGEMA_signal_14354), .Z1_t (new_AGEMA_signal_14355), .Z1_f (new_AGEMA_signal_14356) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1421 ( .A0_t (n796), .A0_f (new_AGEMA_signal_17546), .A1_t (new_AGEMA_signal_17547), .A1_f (new_AGEMA_signal_17548), .B0_t (n795), .B0_f (new_AGEMA_signal_14354), .B1_t (new_AGEMA_signal_14355), .B1_f (new_AGEMA_signal_14356), .Z0_t (RoundOutput[75]), .Z0_f (new_AGEMA_signal_17870), .Z1_t (new_AGEMA_signal_17871), .Z1_f (new_AGEMA_signal_17872) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1422 ( .A0_t (MixColumnsOutput[76]), .A0_f (new_AGEMA_signal_16877), .A1_t (new_AGEMA_signal_16878), .A1_f (new_AGEMA_signal_16879), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n798), .Z0_f (new_AGEMA_signal_17549), .Z1_t (new_AGEMA_signal_17550), .Z1_f (new_AGEMA_signal_17551) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1423 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13670), .B1_t (new_AGEMA_signal_13671), .B1_f (new_AGEMA_signal_13672), .Z0_t (n797), .Z0_f (new_AGEMA_signal_14357), .Z1_t (new_AGEMA_signal_14358), .Z1_f (new_AGEMA_signal_14359) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1424 ( .A0_t (n798), .A0_f (new_AGEMA_signal_17549), .A1_t (new_AGEMA_signal_17550), .A1_f (new_AGEMA_signal_17551), .B0_t (n797), .B0_f (new_AGEMA_signal_14357), .B1_t (new_AGEMA_signal_14358), .B1_f (new_AGEMA_signal_14359), .Z0_t (RoundOutput[76]), .Z0_f (new_AGEMA_signal_17873), .Z1_t (new_AGEMA_signal_17874), .Z1_f (new_AGEMA_signal_17875) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1425 ( .A0_t (MixColumnsOutput[77]), .A0_f (new_AGEMA_signal_15989), .A1_t (new_AGEMA_signal_15990), .A1_f (new_AGEMA_signal_15991), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n800), .Z0_f (new_AGEMA_signal_16760), .Z1_t (new_AGEMA_signal_16761), .Z1_f (new_AGEMA_signal_16762) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1426 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13667), .B1_t (new_AGEMA_signal_13668), .B1_f (new_AGEMA_signal_13669), .Z0_t (n799), .Z0_f (new_AGEMA_signal_14360), .Z1_t (new_AGEMA_signal_14361), .Z1_f (new_AGEMA_signal_14362) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1427 ( .A0_t (n800), .A0_f (new_AGEMA_signal_16760), .A1_t (new_AGEMA_signal_16761), .A1_f (new_AGEMA_signal_16762), .B0_t (n799), .B0_f (new_AGEMA_signal_14360), .B1_t (new_AGEMA_signal_14361), .B1_f (new_AGEMA_signal_14362), .Z0_t (RoundOutput[77]), .Z0_f (new_AGEMA_signal_17552), .Z1_t (new_AGEMA_signal_17553), .Z1_f (new_AGEMA_signal_17554) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1428 ( .A0_t (MixColumnsOutput[78]), .A0_f (new_AGEMA_signal_15986), .A1_t (new_AGEMA_signal_15987), .A1_f (new_AGEMA_signal_15988), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n802), .Z0_f (new_AGEMA_signal_16763), .Z1_t (new_AGEMA_signal_16764), .Z1_f (new_AGEMA_signal_16765) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1429 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13664), .B1_t (new_AGEMA_signal_13665), .B1_f (new_AGEMA_signal_13666), .Z0_t (n801), .Z0_f (new_AGEMA_signal_14363), .Z1_t (new_AGEMA_signal_14364), .Z1_f (new_AGEMA_signal_14365) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1430 ( .A0_t (n802), .A0_f (new_AGEMA_signal_16763), .A1_t (new_AGEMA_signal_16764), .A1_f (new_AGEMA_signal_16765), .B0_t (n801), .B0_f (new_AGEMA_signal_14363), .B1_t (new_AGEMA_signal_14364), .B1_f (new_AGEMA_signal_14365), .Z0_t (RoundOutput[78]), .Z0_f (new_AGEMA_signal_17555), .Z1_t (new_AGEMA_signal_17556), .Z1_f (new_AGEMA_signal_17557) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1431 ( .A0_t (MixColumnsOutput[79]), .A0_f (new_AGEMA_signal_15983), .A1_t (new_AGEMA_signal_15984), .A1_f (new_AGEMA_signal_15985), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n804), .Z0_f (new_AGEMA_signal_16766), .Z1_t (new_AGEMA_signal_16767), .Z1_f (new_AGEMA_signal_16768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1432 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B0_f (new_AGEMA_signal_13661), .B1_t (new_AGEMA_signal_13662), .B1_f (new_AGEMA_signal_13663), .Z0_t (n803), .Z0_f (new_AGEMA_signal_14366), .Z1_t (new_AGEMA_signal_14367), .Z1_f (new_AGEMA_signal_14368) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1433 ( .A0_t (n804), .A0_f (new_AGEMA_signal_16766), .A1_t (new_AGEMA_signal_16767), .A1_f (new_AGEMA_signal_16768), .B0_t (n803), .B0_f (new_AGEMA_signal_14366), .B1_t (new_AGEMA_signal_14367), .B1_f (new_AGEMA_signal_14368), .Z0_t (RoundOutput[79]), .Z0_f (new_AGEMA_signal_17558), .Z1_t (new_AGEMA_signal_17559), .Z1_f (new_AGEMA_signal_17560) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1434 ( .A0_t (MixColumnsOutput[7]), .A0_f (new_AGEMA_signal_16106), .A1_t (new_AGEMA_signal_16107), .A1_f (new_AGEMA_signal_16108), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n806), .Z0_f (new_AGEMA_signal_16769), .Z1_t (new_AGEMA_signal_16770), .Z1_f (new_AGEMA_signal_16771) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1435 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B0_f (new_AGEMA_signal_13724), .B1_t (new_AGEMA_signal_13725), .B1_f (new_AGEMA_signal_13726), .Z0_t (n805), .Z0_f (new_AGEMA_signal_14369), .Z1_t (new_AGEMA_signal_14370), .Z1_f (new_AGEMA_signal_14371) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1436 ( .A0_t (n806), .A0_f (new_AGEMA_signal_16769), .A1_t (new_AGEMA_signal_16770), .A1_f (new_AGEMA_signal_16771), .B0_t (n805), .B0_f (new_AGEMA_signal_14369), .B1_t (new_AGEMA_signal_14370), .B1_f (new_AGEMA_signal_14371), .Z0_t (RoundOutput[7]), .Z0_f (new_AGEMA_signal_17561), .Z1_t (new_AGEMA_signal_17562), .Z1_f (new_AGEMA_signal_17563) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1437 ( .A0_t (MixColumnsOutput[80]), .A0_f (new_AGEMA_signal_15980), .A1_t (new_AGEMA_signal_15981), .A1_f (new_AGEMA_signal_15982), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n808), .Z0_f (new_AGEMA_signal_16772), .Z1_t (new_AGEMA_signal_16773), .Z1_f (new_AGEMA_signal_16774) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1438 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[80]), .B0_f (new_AGEMA_signal_13196), .B1_t (new_AGEMA_signal_13197), .B1_f (new_AGEMA_signal_13198), .Z0_t (n807), .Z0_f (new_AGEMA_signal_13628), .Z1_t (new_AGEMA_signal_13629), .Z1_f (new_AGEMA_signal_13630) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1439 ( .A0_t (n808), .A0_f (new_AGEMA_signal_16772), .A1_t (new_AGEMA_signal_16773), .A1_f (new_AGEMA_signal_16774), .B0_t (n807), .B0_f (new_AGEMA_signal_13628), .B1_t (new_AGEMA_signal_13629), .B1_f (new_AGEMA_signal_13630), .Z0_t (RoundOutput[80]), .Z0_f (new_AGEMA_signal_17564), .Z1_t (new_AGEMA_signal_17565), .Z1_f (new_AGEMA_signal_17566) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1440 ( .A0_t (MixColumnsOutput[81]), .A0_f (new_AGEMA_signal_16874), .A1_t (new_AGEMA_signal_16875), .A1_f (new_AGEMA_signal_16876), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n810), .Z0_f (new_AGEMA_signal_17567), .Z1_t (new_AGEMA_signal_17568), .Z1_f (new_AGEMA_signal_17569) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1441 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13784), .B1_t (new_AGEMA_signal_13785), .B1_f (new_AGEMA_signal_13786), .Z0_t (n809), .Z0_f (new_AGEMA_signal_14372), .Z1_t (new_AGEMA_signal_14373), .Z1_f (new_AGEMA_signal_14374) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1442 ( .A0_t (n810), .A0_f (new_AGEMA_signal_17567), .A1_t (new_AGEMA_signal_17568), .A1_f (new_AGEMA_signal_17569), .B0_t (n809), .B0_f (new_AGEMA_signal_14372), .B1_t (new_AGEMA_signal_14373), .B1_f (new_AGEMA_signal_14374), .Z0_t (RoundOutput[81]), .Z0_f (new_AGEMA_signal_17876), .Z1_t (new_AGEMA_signal_17877), .Z1_f (new_AGEMA_signal_17878) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1443 ( .A0_t (MixColumnsOutput[82]), .A0_f (new_AGEMA_signal_15974), .A1_t (new_AGEMA_signal_15975), .A1_f (new_AGEMA_signal_15976), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n812), .Z0_f (new_AGEMA_signal_16775), .Z1_t (new_AGEMA_signal_16776), .Z1_f (new_AGEMA_signal_16777) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1444 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[82]), .B0_f (new_AGEMA_signal_13781), .B1_t (new_AGEMA_signal_13782), .B1_f (new_AGEMA_signal_13783), .Z0_t (n811), .Z0_f (new_AGEMA_signal_14375), .Z1_t (new_AGEMA_signal_14376), .Z1_f (new_AGEMA_signal_14377) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1445 ( .A0_t (n812), .A0_f (new_AGEMA_signal_16775), .A1_t (new_AGEMA_signal_16776), .A1_f (new_AGEMA_signal_16777), .B0_t (n811), .B0_f (new_AGEMA_signal_14375), .B1_t (new_AGEMA_signal_14376), .B1_f (new_AGEMA_signal_14377), .Z0_t (RoundOutput[82]), .Z0_f (new_AGEMA_signal_17570), .Z1_t (new_AGEMA_signal_17571), .Z1_f (new_AGEMA_signal_17572) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1446 ( .A0_t (MixColumnsOutput[83]), .A0_f (new_AGEMA_signal_16871), .A1_t (new_AGEMA_signal_16872), .A1_f (new_AGEMA_signal_16873), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n814), .Z0_f (new_AGEMA_signal_17573), .Z1_t (new_AGEMA_signal_17574), .Z1_f (new_AGEMA_signal_17575) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1447 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[83]), .B0_f (new_AGEMA_signal_13778), .B1_t (new_AGEMA_signal_13779), .B1_f (new_AGEMA_signal_13780), .Z0_t (n813), .Z0_f (new_AGEMA_signal_14378), .Z1_t (new_AGEMA_signal_14379), .Z1_f (new_AGEMA_signal_14380) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1448 ( .A0_t (n814), .A0_f (new_AGEMA_signal_17573), .A1_t (new_AGEMA_signal_17574), .A1_f (new_AGEMA_signal_17575), .B0_t (n813), .B0_f (new_AGEMA_signal_14378), .B1_t (new_AGEMA_signal_14379), .B1_f (new_AGEMA_signal_14380), .Z0_t (RoundOutput[83]), .Z0_f (new_AGEMA_signal_17879), .Z1_t (new_AGEMA_signal_17880), .Z1_f (new_AGEMA_signal_17881) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1449 ( .A0_t (MixColumnsOutput[84]), .A0_f (new_AGEMA_signal_16865), .A1_t (new_AGEMA_signal_16866), .A1_f (new_AGEMA_signal_16867), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n816), .Z0_f (new_AGEMA_signal_17576), .Z1_t (new_AGEMA_signal_17577), .Z1_f (new_AGEMA_signal_17578) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1450 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13775), .B1_t (new_AGEMA_signal_13776), .B1_f (new_AGEMA_signal_13777), .Z0_t (n815), .Z0_f (new_AGEMA_signal_14381), .Z1_t (new_AGEMA_signal_14382), .Z1_f (new_AGEMA_signal_14383) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1451 ( .A0_t (n816), .A0_f (new_AGEMA_signal_17576), .A1_t (new_AGEMA_signal_17577), .A1_f (new_AGEMA_signal_17578), .B0_t (n815), .B0_f (new_AGEMA_signal_14381), .B1_t (new_AGEMA_signal_14382), .B1_f (new_AGEMA_signal_14383), .Z0_t (RoundOutput[84]), .Z0_f (new_AGEMA_signal_17882), .Z1_t (new_AGEMA_signal_17883), .Z1_f (new_AGEMA_signal_17884) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1452 ( .A0_t (MixColumnsOutput[85]), .A0_f (new_AGEMA_signal_15962), .A1_t (new_AGEMA_signal_15963), .A1_f (new_AGEMA_signal_15964), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n818), .Z0_f (new_AGEMA_signal_16778), .Z1_t (new_AGEMA_signal_16779), .Z1_f (new_AGEMA_signal_16780) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1453 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13772), .B1_t (new_AGEMA_signal_13773), .B1_f (new_AGEMA_signal_13774), .Z0_t (n817), .Z0_f (new_AGEMA_signal_14384), .Z1_t (new_AGEMA_signal_14385), .Z1_f (new_AGEMA_signal_14386) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1454 ( .A0_t (n818), .A0_f (new_AGEMA_signal_16778), .A1_t (new_AGEMA_signal_16779), .A1_f (new_AGEMA_signal_16780), .B0_t (n817), .B0_f (new_AGEMA_signal_14384), .B1_t (new_AGEMA_signal_14385), .B1_f (new_AGEMA_signal_14386), .Z0_t (RoundOutput[85]), .Z0_f (new_AGEMA_signal_17579), .Z1_t (new_AGEMA_signal_17580), .Z1_f (new_AGEMA_signal_17581) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1455 ( .A0_t (MixColumnsOutput[86]), .A0_f (new_AGEMA_signal_15959), .A1_t (new_AGEMA_signal_15960), .A1_f (new_AGEMA_signal_15961), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n820), .Z0_f (new_AGEMA_signal_16781), .Z1_t (new_AGEMA_signal_16782), .Z1_f (new_AGEMA_signal_16783) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1456 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13769), .B1_t (new_AGEMA_signal_13770), .B1_f (new_AGEMA_signal_13771), .Z0_t (n819), .Z0_f (new_AGEMA_signal_14387), .Z1_t (new_AGEMA_signal_14388), .Z1_f (new_AGEMA_signal_14389) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1457 ( .A0_t (n820), .A0_f (new_AGEMA_signal_16781), .A1_t (new_AGEMA_signal_16782), .A1_f (new_AGEMA_signal_16783), .B0_t (n819), .B0_f (new_AGEMA_signal_14387), .B1_t (new_AGEMA_signal_14388), .B1_f (new_AGEMA_signal_14389), .Z0_t (RoundOutput[86]), .Z0_f (new_AGEMA_signal_17582), .Z1_t (new_AGEMA_signal_17583), .Z1_f (new_AGEMA_signal_17584) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1458 ( .A0_t (MixColumnsOutput[87]), .A0_f (new_AGEMA_signal_15956), .A1_t (new_AGEMA_signal_15957), .A1_f (new_AGEMA_signal_15958), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n822), .Z0_f (new_AGEMA_signal_16784), .Z1_t (new_AGEMA_signal_16785), .Z1_f (new_AGEMA_signal_16786) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1459 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13766), .B1_t (new_AGEMA_signal_13767), .B1_f (new_AGEMA_signal_13768), .Z0_t (n821), .Z0_f (new_AGEMA_signal_14390), .Z1_t (new_AGEMA_signal_14391), .Z1_f (new_AGEMA_signal_14392) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1460 ( .A0_t (n822), .A0_f (new_AGEMA_signal_16784), .A1_t (new_AGEMA_signal_16785), .A1_f (new_AGEMA_signal_16786), .B0_t (n821), .B0_f (new_AGEMA_signal_14390), .B1_t (new_AGEMA_signal_14391), .B1_f (new_AGEMA_signal_14392), .Z0_t (RoundOutput[87]), .Z0_f (new_AGEMA_signal_17585), .Z1_t (new_AGEMA_signal_17586), .Z1_f (new_AGEMA_signal_17587) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1461 ( .A0_t (MixColumnsOutput[88]), .A0_f (new_AGEMA_signal_15953), .A1_t (new_AGEMA_signal_15954), .A1_f (new_AGEMA_signal_15955), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n824), .Z0_f (new_AGEMA_signal_16787), .Z1_t (new_AGEMA_signal_16788), .Z1_f (new_AGEMA_signal_16789) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1462 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[88]), .B0_f (new_AGEMA_signal_13361), .B1_t (new_AGEMA_signal_13362), .B1_f (new_AGEMA_signal_13363), .Z0_t (n823), .Z0_f (new_AGEMA_signal_13631), .Z1_t (new_AGEMA_signal_13632), .Z1_f (new_AGEMA_signal_13633) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1463 ( .A0_t (n824), .A0_f (new_AGEMA_signal_16787), .A1_t (new_AGEMA_signal_16788), .A1_f (new_AGEMA_signal_16789), .B0_t (n823), .B0_f (new_AGEMA_signal_13631), .B1_t (new_AGEMA_signal_13632), .B1_f (new_AGEMA_signal_13633), .Z0_t (RoundOutput[88]), .Z0_f (new_AGEMA_signal_17588), .Z1_t (new_AGEMA_signal_17589), .Z1_f (new_AGEMA_signal_17590) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1464 ( .A0_t (MixColumnsOutput[89]), .A0_f (new_AGEMA_signal_16862), .A1_t (new_AGEMA_signal_16863), .A1_f (new_AGEMA_signal_16864), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n826), .Z0_f (new_AGEMA_signal_17591), .Z1_t (new_AGEMA_signal_17592), .Z1_f (new_AGEMA_signal_17593) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1465 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13889), .B1_t (new_AGEMA_signal_13890), .B1_f (new_AGEMA_signal_13891), .Z0_t (n825), .Z0_f (new_AGEMA_signal_14393), .Z1_t (new_AGEMA_signal_14394), .Z1_f (new_AGEMA_signal_14395) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1466 ( .A0_t (n826), .A0_f (new_AGEMA_signal_17591), .A1_t (new_AGEMA_signal_17592), .A1_f (new_AGEMA_signal_17593), .B0_t (n825), .B0_f (new_AGEMA_signal_14393), .B1_t (new_AGEMA_signal_14394), .B1_f (new_AGEMA_signal_14395), .Z0_t (RoundOutput[89]), .Z0_f (new_AGEMA_signal_17885), .Z1_t (new_AGEMA_signal_17886), .Z1_f (new_AGEMA_signal_17887) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1467 ( .A0_t (MixColumnsOutput[8]), .A0_f (new_AGEMA_signal_16103), .A1_t (new_AGEMA_signal_16104), .A1_f (new_AGEMA_signal_16105), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n828), .Z0_f (new_AGEMA_signal_16790), .Z1_t (new_AGEMA_signal_16791), .Z1_f (new_AGEMA_signal_16792) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1468 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[8]), .B0_f (new_AGEMA_signal_13295), .B1_t (new_AGEMA_signal_13296), .B1_f (new_AGEMA_signal_13297), .Z0_t (n827), .Z0_f (new_AGEMA_signal_13634), .Z1_t (new_AGEMA_signal_13635), .Z1_f (new_AGEMA_signal_13636) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1469 ( .A0_t (n828), .A0_f (new_AGEMA_signal_16790), .A1_t (new_AGEMA_signal_16791), .A1_f (new_AGEMA_signal_16792), .B0_t (n827), .B0_f (new_AGEMA_signal_13634), .B1_t (new_AGEMA_signal_13635), .B1_f (new_AGEMA_signal_13636), .Z0_t (RoundOutput[8]), .Z0_f (new_AGEMA_signal_17594), .Z1_t (new_AGEMA_signal_17595), .Z1_f (new_AGEMA_signal_17596) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1470 ( .A0_t (MixColumnsOutput[90]), .A0_f (new_AGEMA_signal_15947), .A1_t (new_AGEMA_signal_15948), .A1_f (new_AGEMA_signal_15949), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n830), .Z0_f (new_AGEMA_signal_16793), .Z1_t (new_AGEMA_signal_16794), .Z1_f (new_AGEMA_signal_16795) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1471 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[90]), .B0_f (new_AGEMA_signal_13886), .B1_t (new_AGEMA_signal_13887), .B1_f (new_AGEMA_signal_13888), .Z0_t (n829), .Z0_f (new_AGEMA_signal_14396), .Z1_t (new_AGEMA_signal_14397), .Z1_f (new_AGEMA_signal_14398) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1472 ( .A0_t (n830), .A0_f (new_AGEMA_signal_16793), .A1_t (new_AGEMA_signal_16794), .A1_f (new_AGEMA_signal_16795), .B0_t (n829), .B0_f (new_AGEMA_signal_14396), .B1_t (new_AGEMA_signal_14397), .B1_f (new_AGEMA_signal_14398), .Z0_t (RoundOutput[90]), .Z0_f (new_AGEMA_signal_17597), .Z1_t (new_AGEMA_signal_17598), .Z1_f (new_AGEMA_signal_17599) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1473 ( .A0_t (MixColumnsOutput[91]), .A0_f (new_AGEMA_signal_16859), .A1_t (new_AGEMA_signal_16860), .A1_f (new_AGEMA_signal_16861), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n832), .Z0_f (new_AGEMA_signal_17600), .Z1_t (new_AGEMA_signal_17601), .Z1_f (new_AGEMA_signal_17602) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1474 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[91]), .B0_f (new_AGEMA_signal_13883), .B1_t (new_AGEMA_signal_13884), .B1_f (new_AGEMA_signal_13885), .Z0_t (n831), .Z0_f (new_AGEMA_signal_14399), .Z1_t (new_AGEMA_signal_14400), .Z1_f (new_AGEMA_signal_14401) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1475 ( .A0_t (n832), .A0_f (new_AGEMA_signal_17600), .A1_t (new_AGEMA_signal_17601), .A1_f (new_AGEMA_signal_17602), .B0_t (n831), .B0_f (new_AGEMA_signal_14399), .B1_t (new_AGEMA_signal_14400), .B1_f (new_AGEMA_signal_14401), .Z0_t (RoundOutput[91]), .Z0_f (new_AGEMA_signal_17888), .Z1_t (new_AGEMA_signal_17889), .Z1_f (new_AGEMA_signal_17890) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1476 ( .A0_t (MixColumnsOutput[92]), .A0_f (new_AGEMA_signal_16856), .A1_t (new_AGEMA_signal_16857), .A1_f (new_AGEMA_signal_16858), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n834), .Z0_f (new_AGEMA_signal_17603), .Z1_t (new_AGEMA_signal_17604), .Z1_f (new_AGEMA_signal_17605) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1477 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13880), .B1_t (new_AGEMA_signal_13881), .B1_f (new_AGEMA_signal_13882), .Z0_t (n833), .Z0_f (new_AGEMA_signal_14402), .Z1_t (new_AGEMA_signal_14403), .Z1_f (new_AGEMA_signal_14404) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1478 ( .A0_t (n834), .A0_f (new_AGEMA_signal_17603), .A1_t (new_AGEMA_signal_17604), .A1_f (new_AGEMA_signal_17605), .B0_t (n833), .B0_f (new_AGEMA_signal_14402), .B1_t (new_AGEMA_signal_14403), .B1_f (new_AGEMA_signal_14404), .Z0_t (RoundOutput[92]), .Z0_f (new_AGEMA_signal_17891), .Z1_t (new_AGEMA_signal_17892), .Z1_f (new_AGEMA_signal_17893) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1479 ( .A0_t (MixColumnsOutput[93]), .A0_f (new_AGEMA_signal_15938), .A1_t (new_AGEMA_signal_15939), .A1_f (new_AGEMA_signal_15940), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n836), .Z0_f (new_AGEMA_signal_16796), .Z1_t (new_AGEMA_signal_16797), .Z1_f (new_AGEMA_signal_16798) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1480 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13877), .B1_t (new_AGEMA_signal_13878), .B1_f (new_AGEMA_signal_13879), .Z0_t (n835), .Z0_f (new_AGEMA_signal_14405), .Z1_t (new_AGEMA_signal_14406), .Z1_f (new_AGEMA_signal_14407) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1481 ( .A0_t (n836), .A0_f (new_AGEMA_signal_16796), .A1_t (new_AGEMA_signal_16797), .A1_f (new_AGEMA_signal_16798), .B0_t (n835), .B0_f (new_AGEMA_signal_14405), .B1_t (new_AGEMA_signal_14406), .B1_f (new_AGEMA_signal_14407), .Z0_t (RoundOutput[93]), .Z0_f (new_AGEMA_signal_17606), .Z1_t (new_AGEMA_signal_17607), .Z1_f (new_AGEMA_signal_17608) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1482 ( .A0_t (MixColumnsOutput[94]), .A0_f (new_AGEMA_signal_15932), .A1_t (new_AGEMA_signal_15933), .A1_f (new_AGEMA_signal_15934), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n838), .Z0_f (new_AGEMA_signal_16799), .Z1_t (new_AGEMA_signal_16800), .Z1_f (new_AGEMA_signal_16801) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1483 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13874), .B1_t (new_AGEMA_signal_13875), .B1_f (new_AGEMA_signal_13876), .Z0_t (n837), .Z0_f (new_AGEMA_signal_14408), .Z1_t (new_AGEMA_signal_14409), .Z1_f (new_AGEMA_signal_14410) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1484 ( .A0_t (n838), .A0_f (new_AGEMA_signal_16799), .A1_t (new_AGEMA_signal_16800), .A1_f (new_AGEMA_signal_16801), .B0_t (n837), .B0_f (new_AGEMA_signal_14408), .B1_t (new_AGEMA_signal_14409), .B1_f (new_AGEMA_signal_14410), .Z0_t (RoundOutput[94]), .Z0_f (new_AGEMA_signal_17609), .Z1_t (new_AGEMA_signal_17610), .Z1_f (new_AGEMA_signal_17611) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1485 ( .A0_t (MixColumnsOutput[95]), .A0_f (new_AGEMA_signal_15929), .A1_t (new_AGEMA_signal_15930), .A1_f (new_AGEMA_signal_15931), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n840), .Z0_f (new_AGEMA_signal_16802), .Z1_t (new_AGEMA_signal_16803), .Z1_f (new_AGEMA_signal_16804) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1486 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13871), .B1_t (new_AGEMA_signal_13872), .B1_f (new_AGEMA_signal_13873), .Z0_t (n839), .Z0_f (new_AGEMA_signal_14411), .Z1_t (new_AGEMA_signal_14412), .Z1_f (new_AGEMA_signal_14413) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1487 ( .A0_t (n840), .A0_f (new_AGEMA_signal_16802), .A1_t (new_AGEMA_signal_16803), .A1_f (new_AGEMA_signal_16804), .B0_t (n839), .B0_f (new_AGEMA_signal_14411), .B1_t (new_AGEMA_signal_14412), .B1_f (new_AGEMA_signal_14413), .Z0_t (RoundOutput[95]), .Z0_f (new_AGEMA_signal_17612), .Z1_t (new_AGEMA_signal_17613), .Z1_f (new_AGEMA_signal_17614) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1488 ( .A0_t (MixColumnsOutput[96]), .A0_f (new_AGEMA_signal_15905), .A1_t (new_AGEMA_signal_15906), .A1_f (new_AGEMA_signal_15907), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n842), .Z0_f (new_AGEMA_signal_16805), .Z1_t (new_AGEMA_signal_16806), .Z1_f (new_AGEMA_signal_16807) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1489 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[96]), .B0_f (new_AGEMA_signal_12998), .B1_t (new_AGEMA_signal_12999), .B1_f (new_AGEMA_signal_13000), .Z0_t (n841), .Z0_f (new_AGEMA_signal_13637), .Z1_t (new_AGEMA_signal_13638), .Z1_f (new_AGEMA_signal_13639) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1490 ( .A0_t (n842), .A0_f (new_AGEMA_signal_16805), .A1_t (new_AGEMA_signal_16806), .A1_f (new_AGEMA_signal_16807), .B0_t (n841), .B0_f (new_AGEMA_signal_13637), .B1_t (new_AGEMA_signal_13638), .B1_f (new_AGEMA_signal_13639), .Z0_t (RoundOutput[96]), .Z0_f (new_AGEMA_signal_17615), .Z1_t (new_AGEMA_signal_17616), .Z1_f (new_AGEMA_signal_17617) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1491 ( .A0_t (MixColumnsOutput[97]), .A0_f (new_AGEMA_signal_16832), .A1_t (new_AGEMA_signal_16833), .A1_f (new_AGEMA_signal_16834), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n844), .Z0_f (new_AGEMA_signal_17618), .Z1_t (new_AGEMA_signal_17619), .Z1_f (new_AGEMA_signal_17620) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1492 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .B0_f (new_AGEMA_signal_13658), .B1_t (new_AGEMA_signal_13659), .B1_f (new_AGEMA_signal_13660), .Z0_t (n843), .Z0_f (new_AGEMA_signal_14414), .Z1_t (new_AGEMA_signal_14415), .Z1_f (new_AGEMA_signal_14416) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1493 ( .A0_t (n844), .A0_f (new_AGEMA_signal_17618), .A1_t (new_AGEMA_signal_17619), .A1_f (new_AGEMA_signal_17620), .B0_t (n843), .B0_f (new_AGEMA_signal_14414), .B1_t (new_AGEMA_signal_14415), .B1_f (new_AGEMA_signal_14416), .Z0_t (RoundOutput[97]), .Z0_f (new_AGEMA_signal_17894), .Z1_t (new_AGEMA_signal_17895), .Z1_f (new_AGEMA_signal_17896) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1494 ( .A0_t (MixColumnsOutput[98]), .A0_f (new_AGEMA_signal_15839), .A1_t (new_AGEMA_signal_15840), .A1_f (new_AGEMA_signal_15841), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n846), .Z0_f (new_AGEMA_signal_16808), .Z1_t (new_AGEMA_signal_16809), .Z1_f (new_AGEMA_signal_16810) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1495 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[98]), .B0_f (new_AGEMA_signal_13655), .B1_t (new_AGEMA_signal_13656), .B1_f (new_AGEMA_signal_13657), .Z0_t (n845), .Z0_f (new_AGEMA_signal_14417), .Z1_t (new_AGEMA_signal_14418), .Z1_f (new_AGEMA_signal_14419) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1496 ( .A0_t (n846), .A0_f (new_AGEMA_signal_16808), .A1_t (new_AGEMA_signal_16809), .A1_f (new_AGEMA_signal_16810), .B0_t (n845), .B0_f (new_AGEMA_signal_14417), .B1_t (new_AGEMA_signal_14418), .B1_f (new_AGEMA_signal_14419), .Z0_t (RoundOutput[98]), .Z0_f (new_AGEMA_signal_17621), .Z1_t (new_AGEMA_signal_17622), .Z1_f (new_AGEMA_signal_17623) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1497 ( .A0_t (MixColumnsOutput[99]), .A0_f (new_AGEMA_signal_16817), .A1_t (new_AGEMA_signal_16818), .A1_f (new_AGEMA_signal_16819), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n848), .Z0_f (new_AGEMA_signal_17624), .Z1_t (new_AGEMA_signal_17625), .Z1_f (new_AGEMA_signal_17626) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1498 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsInput[99]), .B0_f (new_AGEMA_signal_13652), .B1_t (new_AGEMA_signal_13653), .B1_f (new_AGEMA_signal_13654), .Z0_t (n847), .Z0_f (new_AGEMA_signal_14420), .Z1_t (new_AGEMA_signal_14421), .Z1_f (new_AGEMA_signal_14422) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1499 ( .A0_t (n848), .A0_f (new_AGEMA_signal_17624), .A1_t (new_AGEMA_signal_17625), .A1_f (new_AGEMA_signal_17626), .B0_t (n847), .B0_f (new_AGEMA_signal_14420), .B1_t (new_AGEMA_signal_14421), .B1_f (new_AGEMA_signal_14422), .Z0_t (RoundOutput[99]), .Z0_f (new_AGEMA_signal_17897), .Z1_t (new_AGEMA_signal_17898), .Z1_f (new_AGEMA_signal_17899) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1500 ( .A0_t (MixColumnsOutput[9]), .A0_f (new_AGEMA_signal_16919), .A1_t (new_AGEMA_signal_16920), .A1_f (new_AGEMA_signal_16921), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n577), .B1_f (new_AGEMA_signal_6924), .Z0_t (n850), .Z0_f (new_AGEMA_signal_17627), .Z1_t (new_AGEMA_signal_17628), .Z1_f (new_AGEMA_signal_17629) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1501 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n577), .A1_f (new_AGEMA_signal_6924), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13847), .B1_t (new_AGEMA_signal_13848), .B1_f (new_AGEMA_signal_13849), .Z0_t (n849), .Z0_f (new_AGEMA_signal_14423), .Z1_t (new_AGEMA_signal_14424), .Z1_f (new_AGEMA_signal_14425) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1502 ( .A0_t (n850), .A0_f (new_AGEMA_signal_17627), .A1_t (new_AGEMA_signal_17628), .A1_f (new_AGEMA_signal_17629), .B0_t (n849), .B0_f (new_AGEMA_signal_14423), .B1_t (new_AGEMA_signal_14424), .B1_f (new_AGEMA_signal_14425), .Z0_t (RoundOutput[9]), .Z0_f (new_AGEMA_signal_17900), .Z1_t (new_AGEMA_signal_17901), .Z1_f (new_AGEMA_signal_17902) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1503 ( .A0_t (RoundInput[0]), .A0_f (new_AGEMA_signal_5060), .A1_t (new_AGEMA_signal_5061), .A1_f (new_AGEMA_signal_5062), .B0_t (RoundKey[0]), .B0_f (new_AGEMA_signal_5063), .B1_t (new_AGEMA_signal_5064), .B1_f (new_AGEMA_signal_5065), .Z0_t (ciphertext_s0_t[0]), .Z0_f (ciphertext_s0_f[0]), .Z1_t (ciphertext_s1_t[0]), .Z1_f (ciphertext_s1_f[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1504 ( .A0_t (RoundInput[100]), .A0_f (new_AGEMA_signal_5069), .A1_t (new_AGEMA_signal_5070), .A1_f (new_AGEMA_signal_5071), .B0_t (RoundKey[100]), .B0_f (new_AGEMA_signal_5072), .B1_t (new_AGEMA_signal_5073), .B1_f (new_AGEMA_signal_5074), .Z0_t (ciphertext_s0_t[100]), .Z0_f (ciphertext_s0_f[100]), .Z1_t (ciphertext_s1_t[100]), .Z1_f (ciphertext_s1_f[100]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1505 ( .A0_t (RoundInput[101]), .A0_f (new_AGEMA_signal_5078), .A1_t (new_AGEMA_signal_5079), .A1_f (new_AGEMA_signal_5080), .B0_t (RoundKey[101]), .B0_f (new_AGEMA_signal_5081), .B1_t (new_AGEMA_signal_5082), .B1_f (new_AGEMA_signal_5083), .Z0_t (ciphertext_s0_t[101]), .Z0_f (ciphertext_s0_f[101]), .Z1_t (ciphertext_s1_t[101]), .Z1_f (ciphertext_s1_f[101]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1506 ( .A0_t (RoundInput[102]), .A0_f (new_AGEMA_signal_5087), .A1_t (new_AGEMA_signal_5088), .A1_f (new_AGEMA_signal_5089), .B0_t (RoundKey[102]), .B0_f (new_AGEMA_signal_5090), .B1_t (new_AGEMA_signal_5091), .B1_f (new_AGEMA_signal_5092), .Z0_t (ciphertext_s0_t[102]), .Z0_f (ciphertext_s0_f[102]), .Z1_t (ciphertext_s1_t[102]), .Z1_f (ciphertext_s1_f[102]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1507 ( .A0_t (RoundInput[103]), .A0_f (new_AGEMA_signal_5096), .A1_t (new_AGEMA_signal_5097), .A1_f (new_AGEMA_signal_5098), .B0_t (RoundKey[103]), .B0_f (new_AGEMA_signal_5099), .B1_t (new_AGEMA_signal_5100), .B1_f (new_AGEMA_signal_5101), .Z0_t (ciphertext_s0_t[103]), .Z0_f (ciphertext_s0_f[103]), .Z1_t (ciphertext_s1_t[103]), .Z1_f (ciphertext_s1_f[103]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1508 ( .A0_t (RoundInput[104]), .A0_f (new_AGEMA_signal_5105), .A1_t (new_AGEMA_signal_5106), .A1_f (new_AGEMA_signal_5107), .B0_t (RoundKey[104]), .B0_f (new_AGEMA_signal_5108), .B1_t (new_AGEMA_signal_5109), .B1_f (new_AGEMA_signal_5110), .Z0_t (ciphertext_s0_t[104]), .Z0_f (ciphertext_s0_f[104]), .Z1_t (ciphertext_s1_t[104]), .Z1_f (ciphertext_s1_f[104]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1509 ( .A0_t (RoundInput[105]), .A0_f (new_AGEMA_signal_5114), .A1_t (new_AGEMA_signal_5115), .A1_f (new_AGEMA_signal_5116), .B0_t (RoundKey[105]), .B0_f (new_AGEMA_signal_5117), .B1_t (new_AGEMA_signal_5118), .B1_f (new_AGEMA_signal_5119), .Z0_t (ciphertext_s0_t[105]), .Z0_f (ciphertext_s0_f[105]), .Z1_t (ciphertext_s1_t[105]), .Z1_f (ciphertext_s1_f[105]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1510 ( .A0_t (RoundInput[106]), .A0_f (new_AGEMA_signal_5123), .A1_t (new_AGEMA_signal_5124), .A1_f (new_AGEMA_signal_5125), .B0_t (RoundKey[106]), .B0_f (new_AGEMA_signal_5126), .B1_t (new_AGEMA_signal_5127), .B1_f (new_AGEMA_signal_5128), .Z0_t (ciphertext_s0_t[106]), .Z0_f (ciphertext_s0_f[106]), .Z1_t (ciphertext_s1_t[106]), .Z1_f (ciphertext_s1_f[106]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1511 ( .A0_t (RoundInput[107]), .A0_f (new_AGEMA_signal_5132), .A1_t (new_AGEMA_signal_5133), .A1_f (new_AGEMA_signal_5134), .B0_t (RoundKey[107]), .B0_f (new_AGEMA_signal_5135), .B1_t (new_AGEMA_signal_5136), .B1_f (new_AGEMA_signal_5137), .Z0_t (ciphertext_s0_t[107]), .Z0_f (ciphertext_s0_f[107]), .Z1_t (ciphertext_s1_t[107]), .Z1_f (ciphertext_s1_f[107]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1512 ( .A0_t (RoundInput[108]), .A0_f (new_AGEMA_signal_5141), .A1_t (new_AGEMA_signal_5142), .A1_f (new_AGEMA_signal_5143), .B0_t (RoundKey[108]), .B0_f (new_AGEMA_signal_5144), .B1_t (new_AGEMA_signal_5145), .B1_f (new_AGEMA_signal_5146), .Z0_t (ciphertext_s0_t[108]), .Z0_f (ciphertext_s0_f[108]), .Z1_t (ciphertext_s1_t[108]), .Z1_f (ciphertext_s1_f[108]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1513 ( .A0_t (RoundInput[109]), .A0_f (new_AGEMA_signal_5150), .A1_t (new_AGEMA_signal_5151), .A1_f (new_AGEMA_signal_5152), .B0_t (RoundKey[109]), .B0_f (new_AGEMA_signal_5153), .B1_t (new_AGEMA_signal_5154), .B1_f (new_AGEMA_signal_5155), .Z0_t (ciphertext_s0_t[109]), .Z0_f (ciphertext_s0_f[109]), .Z1_t (ciphertext_s1_t[109]), .Z1_f (ciphertext_s1_f[109]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1514 ( .A0_t (RoundInput[10]), .A0_f (new_AGEMA_signal_5159), .A1_t (new_AGEMA_signal_5160), .A1_f (new_AGEMA_signal_5161), .B0_t (RoundKey[10]), .B0_f (new_AGEMA_signal_5162), .B1_t (new_AGEMA_signal_5163), .B1_f (new_AGEMA_signal_5164), .Z0_t (ciphertext_s0_t[10]), .Z0_f (ciphertext_s0_f[10]), .Z1_t (ciphertext_s1_t[10]), .Z1_f (ciphertext_s1_f[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1515 ( .A0_t (RoundInput[110]), .A0_f (new_AGEMA_signal_5168), .A1_t (new_AGEMA_signal_5169), .A1_f (new_AGEMA_signal_5170), .B0_t (RoundKey[110]), .B0_f (new_AGEMA_signal_5171), .B1_t (new_AGEMA_signal_5172), .B1_f (new_AGEMA_signal_5173), .Z0_t (ciphertext_s0_t[110]), .Z0_f (ciphertext_s0_f[110]), .Z1_t (ciphertext_s1_t[110]), .Z1_f (ciphertext_s1_f[110]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1516 ( .A0_t (RoundInput[111]), .A0_f (new_AGEMA_signal_5177), .A1_t (new_AGEMA_signal_5178), .A1_f (new_AGEMA_signal_5179), .B0_t (RoundKey[111]), .B0_f (new_AGEMA_signal_5180), .B1_t (new_AGEMA_signal_5181), .B1_f (new_AGEMA_signal_5182), .Z0_t (ciphertext_s0_t[111]), .Z0_f (ciphertext_s0_f[111]), .Z1_t (ciphertext_s1_t[111]), .Z1_f (ciphertext_s1_f[111]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1517 ( .A0_t (RoundInput[112]), .A0_f (new_AGEMA_signal_5186), .A1_t (new_AGEMA_signal_5187), .A1_f (new_AGEMA_signal_5188), .B0_t (RoundKey[112]), .B0_f (new_AGEMA_signal_5189), .B1_t (new_AGEMA_signal_5190), .B1_f (new_AGEMA_signal_5191), .Z0_t (ciphertext_s0_t[112]), .Z0_f (ciphertext_s0_f[112]), .Z1_t (ciphertext_s1_t[112]), .Z1_f (ciphertext_s1_f[112]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1518 ( .A0_t (RoundInput[113]), .A0_f (new_AGEMA_signal_5195), .A1_t (new_AGEMA_signal_5196), .A1_f (new_AGEMA_signal_5197), .B0_t (RoundKey[113]), .B0_f (new_AGEMA_signal_5198), .B1_t (new_AGEMA_signal_5199), .B1_f (new_AGEMA_signal_5200), .Z0_t (ciphertext_s0_t[113]), .Z0_f (ciphertext_s0_f[113]), .Z1_t (ciphertext_s1_t[113]), .Z1_f (ciphertext_s1_f[113]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1519 ( .A0_t (RoundInput[114]), .A0_f (new_AGEMA_signal_5204), .A1_t (new_AGEMA_signal_5205), .A1_f (new_AGEMA_signal_5206), .B0_t (RoundKey[114]), .B0_f (new_AGEMA_signal_5207), .B1_t (new_AGEMA_signal_5208), .B1_f (new_AGEMA_signal_5209), .Z0_t (ciphertext_s0_t[114]), .Z0_f (ciphertext_s0_f[114]), .Z1_t (ciphertext_s1_t[114]), .Z1_f (ciphertext_s1_f[114]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1520 ( .A0_t (RoundInput[115]), .A0_f (new_AGEMA_signal_5213), .A1_t (new_AGEMA_signal_5214), .A1_f (new_AGEMA_signal_5215), .B0_t (RoundKey[115]), .B0_f (new_AGEMA_signal_5216), .B1_t (new_AGEMA_signal_5217), .B1_f (new_AGEMA_signal_5218), .Z0_t (ciphertext_s0_t[115]), .Z0_f (ciphertext_s0_f[115]), .Z1_t (ciphertext_s1_t[115]), .Z1_f (ciphertext_s1_f[115]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1521 ( .A0_t (RoundInput[116]), .A0_f (new_AGEMA_signal_5222), .A1_t (new_AGEMA_signal_5223), .A1_f (new_AGEMA_signal_5224), .B0_t (RoundKey[116]), .B0_f (new_AGEMA_signal_5225), .B1_t (new_AGEMA_signal_5226), .B1_f (new_AGEMA_signal_5227), .Z0_t (ciphertext_s0_t[116]), .Z0_f (ciphertext_s0_f[116]), .Z1_t (ciphertext_s1_t[116]), .Z1_f (ciphertext_s1_f[116]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1522 ( .A0_t (RoundInput[117]), .A0_f (new_AGEMA_signal_5231), .A1_t (new_AGEMA_signal_5232), .A1_f (new_AGEMA_signal_5233), .B0_t (RoundKey[117]), .B0_f (new_AGEMA_signal_5234), .B1_t (new_AGEMA_signal_5235), .B1_f (new_AGEMA_signal_5236), .Z0_t (ciphertext_s0_t[117]), .Z0_f (ciphertext_s0_f[117]), .Z1_t (ciphertext_s1_t[117]), .Z1_f (ciphertext_s1_f[117]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1523 ( .A0_t (RoundInput[118]), .A0_f (new_AGEMA_signal_5240), .A1_t (new_AGEMA_signal_5241), .A1_f (new_AGEMA_signal_5242), .B0_t (RoundKey[118]), .B0_f (new_AGEMA_signal_5243), .B1_t (new_AGEMA_signal_5244), .B1_f (new_AGEMA_signal_5245), .Z0_t (ciphertext_s0_t[118]), .Z0_f (ciphertext_s0_f[118]), .Z1_t (ciphertext_s1_t[118]), .Z1_f (ciphertext_s1_f[118]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1524 ( .A0_t (RoundInput[119]), .A0_f (new_AGEMA_signal_5249), .A1_t (new_AGEMA_signal_5250), .A1_f (new_AGEMA_signal_5251), .B0_t (RoundKey[119]), .B0_f (new_AGEMA_signal_5252), .B1_t (new_AGEMA_signal_5253), .B1_f (new_AGEMA_signal_5254), .Z0_t (ciphertext_s0_t[119]), .Z0_f (ciphertext_s0_f[119]), .Z1_t (ciphertext_s1_t[119]), .Z1_f (ciphertext_s1_f[119]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1525 ( .A0_t (RoundInput[11]), .A0_f (new_AGEMA_signal_5258), .A1_t (new_AGEMA_signal_5259), .A1_f (new_AGEMA_signal_5260), .B0_t (RoundKey[11]), .B0_f (new_AGEMA_signal_5261), .B1_t (new_AGEMA_signal_5262), .B1_f (new_AGEMA_signal_5263), .Z0_t (ciphertext_s0_t[11]), .Z0_f (ciphertext_s0_f[11]), .Z1_t (ciphertext_s1_t[11]), .Z1_f (ciphertext_s1_f[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1526 ( .A0_t (RoundInput[120]), .A0_f (new_AGEMA_signal_5267), .A1_t (new_AGEMA_signal_5268), .A1_f (new_AGEMA_signal_5269), .B0_t (RoundKey[120]), .B0_f (new_AGEMA_signal_5270), .B1_t (new_AGEMA_signal_5271), .B1_f (new_AGEMA_signal_5272), .Z0_t (ciphertext_s0_t[120]), .Z0_f (ciphertext_s0_f[120]), .Z1_t (ciphertext_s1_t[120]), .Z1_f (ciphertext_s1_f[120]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1527 ( .A0_t (RoundInput[121]), .A0_f (new_AGEMA_signal_5276), .A1_t (new_AGEMA_signal_5277), .A1_f (new_AGEMA_signal_5278), .B0_t (RoundKey[121]), .B0_f (new_AGEMA_signal_5279), .B1_t (new_AGEMA_signal_5280), .B1_f (new_AGEMA_signal_5281), .Z0_t (ciphertext_s0_t[121]), .Z0_f (ciphertext_s0_f[121]), .Z1_t (ciphertext_s1_t[121]), .Z1_f (ciphertext_s1_f[121]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1528 ( .A0_t (RoundInput[122]), .A0_f (new_AGEMA_signal_5285), .A1_t (new_AGEMA_signal_5286), .A1_f (new_AGEMA_signal_5287), .B0_t (RoundKey[122]), .B0_f (new_AGEMA_signal_5288), .B1_t (new_AGEMA_signal_5289), .B1_f (new_AGEMA_signal_5290), .Z0_t (ciphertext_s0_t[122]), .Z0_f (ciphertext_s0_f[122]), .Z1_t (ciphertext_s1_t[122]), .Z1_f (ciphertext_s1_f[122]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1529 ( .A0_t (RoundInput[123]), .A0_f (new_AGEMA_signal_5294), .A1_t (new_AGEMA_signal_5295), .A1_f (new_AGEMA_signal_5296), .B0_t (RoundKey[123]), .B0_f (new_AGEMA_signal_5297), .B1_t (new_AGEMA_signal_5298), .B1_f (new_AGEMA_signal_5299), .Z0_t (ciphertext_s0_t[123]), .Z0_f (ciphertext_s0_f[123]), .Z1_t (ciphertext_s1_t[123]), .Z1_f (ciphertext_s1_f[123]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1530 ( .A0_t (RoundInput[124]), .A0_f (new_AGEMA_signal_5303), .A1_t (new_AGEMA_signal_5304), .A1_f (new_AGEMA_signal_5305), .B0_t (RoundKey[124]), .B0_f (new_AGEMA_signal_5306), .B1_t (new_AGEMA_signal_5307), .B1_f (new_AGEMA_signal_5308), .Z0_t (ciphertext_s0_t[124]), .Z0_f (ciphertext_s0_f[124]), .Z1_t (ciphertext_s1_t[124]), .Z1_f (ciphertext_s1_f[124]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1531 ( .A0_t (RoundInput[125]), .A0_f (new_AGEMA_signal_5312), .A1_t (new_AGEMA_signal_5313), .A1_f (new_AGEMA_signal_5314), .B0_t (RoundKey[125]), .B0_f (new_AGEMA_signal_5315), .B1_t (new_AGEMA_signal_5316), .B1_f (new_AGEMA_signal_5317), .Z0_t (ciphertext_s0_t[125]), .Z0_f (ciphertext_s0_f[125]), .Z1_t (ciphertext_s1_t[125]), .Z1_f (ciphertext_s1_f[125]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1532 ( .A0_t (RoundInput[126]), .A0_f (new_AGEMA_signal_5321), .A1_t (new_AGEMA_signal_5322), .A1_f (new_AGEMA_signal_5323), .B0_t (RoundKey[126]), .B0_f (new_AGEMA_signal_5324), .B1_t (new_AGEMA_signal_5325), .B1_f (new_AGEMA_signal_5326), .Z0_t (ciphertext_s0_t[126]), .Z0_f (ciphertext_s0_f[126]), .Z1_t (ciphertext_s1_t[126]), .Z1_f (ciphertext_s1_f[126]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1533 ( .A0_t (RoundInput[127]), .A0_f (new_AGEMA_signal_5330), .A1_t (new_AGEMA_signal_5331), .A1_f (new_AGEMA_signal_5332), .B0_t (RoundKey[127]), .B0_f (new_AGEMA_signal_5333), .B1_t (new_AGEMA_signal_5334), .B1_f (new_AGEMA_signal_5335), .Z0_t (ciphertext_s0_t[127]), .Z0_f (ciphertext_s0_f[127]), .Z1_t (ciphertext_s1_t[127]), .Z1_f (ciphertext_s1_f[127]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1534 ( .A0_t (RoundInput[12]), .A0_f (new_AGEMA_signal_5339), .A1_t (new_AGEMA_signal_5340), .A1_f (new_AGEMA_signal_5341), .B0_t (RoundKey[12]), .B0_f (new_AGEMA_signal_5342), .B1_t (new_AGEMA_signal_5343), .B1_f (new_AGEMA_signal_5344), .Z0_t (ciphertext_s0_t[12]), .Z0_f (ciphertext_s0_f[12]), .Z1_t (ciphertext_s1_t[12]), .Z1_f (ciphertext_s1_f[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1535 ( .A0_t (RoundInput[13]), .A0_f (new_AGEMA_signal_5348), .A1_t (new_AGEMA_signal_5349), .A1_f (new_AGEMA_signal_5350), .B0_t (RoundKey[13]), .B0_f (new_AGEMA_signal_5351), .B1_t (new_AGEMA_signal_5352), .B1_f (new_AGEMA_signal_5353), .Z0_t (ciphertext_s0_t[13]), .Z0_f (ciphertext_s0_f[13]), .Z1_t (ciphertext_s1_t[13]), .Z1_f (ciphertext_s1_f[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1536 ( .A0_t (RoundInput[14]), .A0_f (new_AGEMA_signal_5357), .A1_t (new_AGEMA_signal_5358), .A1_f (new_AGEMA_signal_5359), .B0_t (RoundKey[14]), .B0_f (new_AGEMA_signal_5360), .B1_t (new_AGEMA_signal_5361), .B1_f (new_AGEMA_signal_5362), .Z0_t (ciphertext_s0_t[14]), .Z0_f (ciphertext_s0_f[14]), .Z1_t (ciphertext_s1_t[14]), .Z1_f (ciphertext_s1_f[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1537 ( .A0_t (RoundInput[15]), .A0_f (new_AGEMA_signal_5366), .A1_t (new_AGEMA_signal_5367), .A1_f (new_AGEMA_signal_5368), .B0_t (RoundKey[15]), .B0_f (new_AGEMA_signal_5369), .B1_t (new_AGEMA_signal_5370), .B1_f (new_AGEMA_signal_5371), .Z0_t (ciphertext_s0_t[15]), .Z0_f (ciphertext_s0_f[15]), .Z1_t (ciphertext_s1_t[15]), .Z1_f (ciphertext_s1_f[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1538 ( .A0_t (RoundInput[16]), .A0_f (new_AGEMA_signal_5375), .A1_t (new_AGEMA_signal_5376), .A1_f (new_AGEMA_signal_5377), .B0_t (RoundKey[16]), .B0_f (new_AGEMA_signal_5378), .B1_t (new_AGEMA_signal_5379), .B1_f (new_AGEMA_signal_5380), .Z0_t (ciphertext_s0_t[16]), .Z0_f (ciphertext_s0_f[16]), .Z1_t (ciphertext_s1_t[16]), .Z1_f (ciphertext_s1_f[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1539 ( .A0_t (RoundInput[17]), .A0_f (new_AGEMA_signal_5384), .A1_t (new_AGEMA_signal_5385), .A1_f (new_AGEMA_signal_5386), .B0_t (RoundKey[17]), .B0_f (new_AGEMA_signal_5387), .B1_t (new_AGEMA_signal_5388), .B1_f (new_AGEMA_signal_5389), .Z0_t (ciphertext_s0_t[17]), .Z0_f (ciphertext_s0_f[17]), .Z1_t (ciphertext_s1_t[17]), .Z1_f (ciphertext_s1_f[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1540 ( .A0_t (RoundInput[18]), .A0_f (new_AGEMA_signal_5393), .A1_t (new_AGEMA_signal_5394), .A1_f (new_AGEMA_signal_5395), .B0_t (RoundKey[18]), .B0_f (new_AGEMA_signal_5396), .B1_t (new_AGEMA_signal_5397), .B1_f (new_AGEMA_signal_5398), .Z0_t (ciphertext_s0_t[18]), .Z0_f (ciphertext_s0_f[18]), .Z1_t (ciphertext_s1_t[18]), .Z1_f (ciphertext_s1_f[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1541 ( .A0_t (RoundInput[19]), .A0_f (new_AGEMA_signal_5402), .A1_t (new_AGEMA_signal_5403), .A1_f (new_AGEMA_signal_5404), .B0_t (RoundKey[19]), .B0_f (new_AGEMA_signal_5405), .B1_t (new_AGEMA_signal_5406), .B1_f (new_AGEMA_signal_5407), .Z0_t (ciphertext_s0_t[19]), .Z0_f (ciphertext_s0_f[19]), .Z1_t (ciphertext_s1_t[19]), .Z1_f (ciphertext_s1_f[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1542 ( .A0_t (RoundInput[1]), .A0_f (new_AGEMA_signal_5411), .A1_t (new_AGEMA_signal_5412), .A1_f (new_AGEMA_signal_5413), .B0_t (RoundKey[1]), .B0_f (new_AGEMA_signal_5414), .B1_t (new_AGEMA_signal_5415), .B1_f (new_AGEMA_signal_5416), .Z0_t (ciphertext_s0_t[1]), .Z0_f (ciphertext_s0_f[1]), .Z1_t (ciphertext_s1_t[1]), .Z1_f (ciphertext_s1_f[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1543 ( .A0_t (RoundInput[20]), .A0_f (new_AGEMA_signal_5420), .A1_t (new_AGEMA_signal_5421), .A1_f (new_AGEMA_signal_5422), .B0_t (RoundKey[20]), .B0_f (new_AGEMA_signal_5423), .B1_t (new_AGEMA_signal_5424), .B1_f (new_AGEMA_signal_5425), .Z0_t (ciphertext_s0_t[20]), .Z0_f (ciphertext_s0_f[20]), .Z1_t (ciphertext_s1_t[20]), .Z1_f (ciphertext_s1_f[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1544 ( .A0_t (RoundInput[21]), .A0_f (new_AGEMA_signal_5429), .A1_t (new_AGEMA_signal_5430), .A1_f (new_AGEMA_signal_5431), .B0_t (RoundKey[21]), .B0_f (new_AGEMA_signal_5432), .B1_t (new_AGEMA_signal_5433), .B1_f (new_AGEMA_signal_5434), .Z0_t (ciphertext_s0_t[21]), .Z0_f (ciphertext_s0_f[21]), .Z1_t (ciphertext_s1_t[21]), .Z1_f (ciphertext_s1_f[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1545 ( .A0_t (RoundInput[22]), .A0_f (new_AGEMA_signal_5438), .A1_t (new_AGEMA_signal_5439), .A1_f (new_AGEMA_signal_5440), .B0_t (RoundKey[22]), .B0_f (new_AGEMA_signal_5441), .B1_t (new_AGEMA_signal_5442), .B1_f (new_AGEMA_signal_5443), .Z0_t (ciphertext_s0_t[22]), .Z0_f (ciphertext_s0_f[22]), .Z1_t (ciphertext_s1_t[22]), .Z1_f (ciphertext_s1_f[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1546 ( .A0_t (RoundInput[23]), .A0_f (new_AGEMA_signal_5447), .A1_t (new_AGEMA_signal_5448), .A1_f (new_AGEMA_signal_5449), .B0_t (RoundKey[23]), .B0_f (new_AGEMA_signal_5450), .B1_t (new_AGEMA_signal_5451), .B1_f (new_AGEMA_signal_5452), .Z0_t (ciphertext_s0_t[23]), .Z0_f (ciphertext_s0_f[23]), .Z1_t (ciphertext_s1_t[23]), .Z1_f (ciphertext_s1_f[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1547 ( .A0_t (RoundInput[24]), .A0_f (new_AGEMA_signal_5456), .A1_t (new_AGEMA_signal_5457), .A1_f (new_AGEMA_signal_5458), .B0_t (RoundKey[24]), .B0_f (new_AGEMA_signal_5459), .B1_t (new_AGEMA_signal_5460), .B1_f (new_AGEMA_signal_5461), .Z0_t (ciphertext_s0_t[24]), .Z0_f (ciphertext_s0_f[24]), .Z1_t (ciphertext_s1_t[24]), .Z1_f (ciphertext_s1_f[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1548 ( .A0_t (RoundInput[25]), .A0_f (new_AGEMA_signal_5465), .A1_t (new_AGEMA_signal_5466), .A1_f (new_AGEMA_signal_5467), .B0_t (RoundKey[25]), .B0_f (new_AGEMA_signal_5468), .B1_t (new_AGEMA_signal_5469), .B1_f (new_AGEMA_signal_5470), .Z0_t (ciphertext_s0_t[25]), .Z0_f (ciphertext_s0_f[25]), .Z1_t (ciphertext_s1_t[25]), .Z1_f (ciphertext_s1_f[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1549 ( .A0_t (RoundInput[26]), .A0_f (new_AGEMA_signal_5474), .A1_t (new_AGEMA_signal_5475), .A1_f (new_AGEMA_signal_5476), .B0_t (RoundKey[26]), .B0_f (new_AGEMA_signal_5477), .B1_t (new_AGEMA_signal_5478), .B1_f (new_AGEMA_signal_5479), .Z0_t (ciphertext_s0_t[26]), .Z0_f (ciphertext_s0_f[26]), .Z1_t (ciphertext_s1_t[26]), .Z1_f (ciphertext_s1_f[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1550 ( .A0_t (RoundInput[27]), .A0_f (new_AGEMA_signal_5483), .A1_t (new_AGEMA_signal_5484), .A1_f (new_AGEMA_signal_5485), .B0_t (RoundKey[27]), .B0_f (new_AGEMA_signal_5486), .B1_t (new_AGEMA_signal_5487), .B1_f (new_AGEMA_signal_5488), .Z0_t (ciphertext_s0_t[27]), .Z0_f (ciphertext_s0_f[27]), .Z1_t (ciphertext_s1_t[27]), .Z1_f (ciphertext_s1_f[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1551 ( .A0_t (RoundInput[28]), .A0_f (new_AGEMA_signal_5492), .A1_t (new_AGEMA_signal_5493), .A1_f (new_AGEMA_signal_5494), .B0_t (RoundKey[28]), .B0_f (new_AGEMA_signal_5495), .B1_t (new_AGEMA_signal_5496), .B1_f (new_AGEMA_signal_5497), .Z0_t (ciphertext_s0_t[28]), .Z0_f (ciphertext_s0_f[28]), .Z1_t (ciphertext_s1_t[28]), .Z1_f (ciphertext_s1_f[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1552 ( .A0_t (RoundInput[29]), .A0_f (new_AGEMA_signal_5501), .A1_t (new_AGEMA_signal_5502), .A1_f (new_AGEMA_signal_5503), .B0_t (RoundKey[29]), .B0_f (new_AGEMA_signal_5504), .B1_t (new_AGEMA_signal_5505), .B1_f (new_AGEMA_signal_5506), .Z0_t (ciphertext_s0_t[29]), .Z0_f (ciphertext_s0_f[29]), .Z1_t (ciphertext_s1_t[29]), .Z1_f (ciphertext_s1_f[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1553 ( .A0_t (RoundInput[2]), .A0_f (new_AGEMA_signal_5510), .A1_t (new_AGEMA_signal_5511), .A1_f (new_AGEMA_signal_5512), .B0_t (RoundKey[2]), .B0_f (new_AGEMA_signal_5513), .B1_t (new_AGEMA_signal_5514), .B1_f (new_AGEMA_signal_5515), .Z0_t (ciphertext_s0_t[2]), .Z0_f (ciphertext_s0_f[2]), .Z1_t (ciphertext_s1_t[2]), .Z1_f (ciphertext_s1_f[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1554 ( .A0_t (RoundInput[30]), .A0_f (new_AGEMA_signal_5519), .A1_t (new_AGEMA_signal_5520), .A1_f (new_AGEMA_signal_5521), .B0_t (RoundKey[30]), .B0_f (new_AGEMA_signal_5522), .B1_t (new_AGEMA_signal_5523), .B1_f (new_AGEMA_signal_5524), .Z0_t (ciphertext_s0_t[30]), .Z0_f (ciphertext_s0_f[30]), .Z1_t (ciphertext_s1_t[30]), .Z1_f (ciphertext_s1_f[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1555 ( .A0_t (RoundInput[31]), .A0_f (new_AGEMA_signal_5528), .A1_t (new_AGEMA_signal_5529), .A1_f (new_AGEMA_signal_5530), .B0_t (RoundKey[31]), .B0_f (new_AGEMA_signal_5531), .B1_t (new_AGEMA_signal_5532), .B1_f (new_AGEMA_signal_5533), .Z0_t (ciphertext_s0_t[31]), .Z0_f (ciphertext_s0_f[31]), .Z1_t (ciphertext_s1_t[31]), .Z1_f (ciphertext_s1_f[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1556 ( .A0_t (RoundInput[32]), .A0_f (new_AGEMA_signal_5537), .A1_t (new_AGEMA_signal_5538), .A1_f (new_AGEMA_signal_5539), .B0_t (RoundKey[32]), .B0_f (new_AGEMA_signal_5540), .B1_t (new_AGEMA_signal_5541), .B1_f (new_AGEMA_signal_5542), .Z0_t (ciphertext_s0_t[32]), .Z0_f (ciphertext_s0_f[32]), .Z1_t (ciphertext_s1_t[32]), .Z1_f (ciphertext_s1_f[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1557 ( .A0_t (RoundInput[33]), .A0_f (new_AGEMA_signal_5546), .A1_t (new_AGEMA_signal_5547), .A1_f (new_AGEMA_signal_5548), .B0_t (RoundKey[33]), .B0_f (new_AGEMA_signal_5549), .B1_t (new_AGEMA_signal_5550), .B1_f (new_AGEMA_signal_5551), .Z0_t (ciphertext_s0_t[33]), .Z0_f (ciphertext_s0_f[33]), .Z1_t (ciphertext_s1_t[33]), .Z1_f (ciphertext_s1_f[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1558 ( .A0_t (RoundInput[34]), .A0_f (new_AGEMA_signal_5555), .A1_t (new_AGEMA_signal_5556), .A1_f (new_AGEMA_signal_5557), .B0_t (RoundKey[34]), .B0_f (new_AGEMA_signal_5558), .B1_t (new_AGEMA_signal_5559), .B1_f (new_AGEMA_signal_5560), .Z0_t (ciphertext_s0_t[34]), .Z0_f (ciphertext_s0_f[34]), .Z1_t (ciphertext_s1_t[34]), .Z1_f (ciphertext_s1_f[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1559 ( .A0_t (RoundInput[35]), .A0_f (new_AGEMA_signal_5564), .A1_t (new_AGEMA_signal_5565), .A1_f (new_AGEMA_signal_5566), .B0_t (RoundKey[35]), .B0_f (new_AGEMA_signal_5567), .B1_t (new_AGEMA_signal_5568), .B1_f (new_AGEMA_signal_5569), .Z0_t (ciphertext_s0_t[35]), .Z0_f (ciphertext_s0_f[35]), .Z1_t (ciphertext_s1_t[35]), .Z1_f (ciphertext_s1_f[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1560 ( .A0_t (RoundInput[36]), .A0_f (new_AGEMA_signal_5573), .A1_t (new_AGEMA_signal_5574), .A1_f (new_AGEMA_signal_5575), .B0_t (RoundKey[36]), .B0_f (new_AGEMA_signal_5576), .B1_t (new_AGEMA_signal_5577), .B1_f (new_AGEMA_signal_5578), .Z0_t (ciphertext_s0_t[36]), .Z0_f (ciphertext_s0_f[36]), .Z1_t (ciphertext_s1_t[36]), .Z1_f (ciphertext_s1_f[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1561 ( .A0_t (RoundInput[37]), .A0_f (new_AGEMA_signal_5582), .A1_t (new_AGEMA_signal_5583), .A1_f (new_AGEMA_signal_5584), .B0_t (RoundKey[37]), .B0_f (new_AGEMA_signal_5585), .B1_t (new_AGEMA_signal_5586), .B1_f (new_AGEMA_signal_5587), .Z0_t (ciphertext_s0_t[37]), .Z0_f (ciphertext_s0_f[37]), .Z1_t (ciphertext_s1_t[37]), .Z1_f (ciphertext_s1_f[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1562 ( .A0_t (RoundInput[38]), .A0_f (new_AGEMA_signal_5591), .A1_t (new_AGEMA_signal_5592), .A1_f (new_AGEMA_signal_5593), .B0_t (RoundKey[38]), .B0_f (new_AGEMA_signal_5594), .B1_t (new_AGEMA_signal_5595), .B1_f (new_AGEMA_signal_5596), .Z0_t (ciphertext_s0_t[38]), .Z0_f (ciphertext_s0_f[38]), .Z1_t (ciphertext_s1_t[38]), .Z1_f (ciphertext_s1_f[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1563 ( .A0_t (RoundInput[39]), .A0_f (new_AGEMA_signal_5600), .A1_t (new_AGEMA_signal_5601), .A1_f (new_AGEMA_signal_5602), .B0_t (RoundKey[39]), .B0_f (new_AGEMA_signal_5603), .B1_t (new_AGEMA_signal_5604), .B1_f (new_AGEMA_signal_5605), .Z0_t (ciphertext_s0_t[39]), .Z0_f (ciphertext_s0_f[39]), .Z1_t (ciphertext_s1_t[39]), .Z1_f (ciphertext_s1_f[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1564 ( .A0_t (RoundInput[3]), .A0_f (new_AGEMA_signal_5609), .A1_t (new_AGEMA_signal_5610), .A1_f (new_AGEMA_signal_5611), .B0_t (RoundKey[3]), .B0_f (new_AGEMA_signal_5612), .B1_t (new_AGEMA_signal_5613), .B1_f (new_AGEMA_signal_5614), .Z0_t (ciphertext_s0_t[3]), .Z0_f (ciphertext_s0_f[3]), .Z1_t (ciphertext_s1_t[3]), .Z1_f (ciphertext_s1_f[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1565 ( .A0_t (RoundInput[40]), .A0_f (new_AGEMA_signal_5618), .A1_t (new_AGEMA_signal_5619), .A1_f (new_AGEMA_signal_5620), .B0_t (RoundKey[40]), .B0_f (new_AGEMA_signal_5621), .B1_t (new_AGEMA_signal_5622), .B1_f (new_AGEMA_signal_5623), .Z0_t (ciphertext_s0_t[40]), .Z0_f (ciphertext_s0_f[40]), .Z1_t (ciphertext_s1_t[40]), .Z1_f (ciphertext_s1_f[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1566 ( .A0_t (RoundInput[41]), .A0_f (new_AGEMA_signal_5627), .A1_t (new_AGEMA_signal_5628), .A1_f (new_AGEMA_signal_5629), .B0_t (RoundKey[41]), .B0_f (new_AGEMA_signal_5630), .B1_t (new_AGEMA_signal_5631), .B1_f (new_AGEMA_signal_5632), .Z0_t (ciphertext_s0_t[41]), .Z0_f (ciphertext_s0_f[41]), .Z1_t (ciphertext_s1_t[41]), .Z1_f (ciphertext_s1_f[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1567 ( .A0_t (RoundInput[42]), .A0_f (new_AGEMA_signal_5636), .A1_t (new_AGEMA_signal_5637), .A1_f (new_AGEMA_signal_5638), .B0_t (RoundKey[42]), .B0_f (new_AGEMA_signal_5639), .B1_t (new_AGEMA_signal_5640), .B1_f (new_AGEMA_signal_5641), .Z0_t (ciphertext_s0_t[42]), .Z0_f (ciphertext_s0_f[42]), .Z1_t (ciphertext_s1_t[42]), .Z1_f (ciphertext_s1_f[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1568 ( .A0_t (RoundInput[43]), .A0_f (new_AGEMA_signal_5645), .A1_t (new_AGEMA_signal_5646), .A1_f (new_AGEMA_signal_5647), .B0_t (RoundKey[43]), .B0_f (new_AGEMA_signal_5648), .B1_t (new_AGEMA_signal_5649), .B1_f (new_AGEMA_signal_5650), .Z0_t (ciphertext_s0_t[43]), .Z0_f (ciphertext_s0_f[43]), .Z1_t (ciphertext_s1_t[43]), .Z1_f (ciphertext_s1_f[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1569 ( .A0_t (RoundInput[44]), .A0_f (new_AGEMA_signal_5654), .A1_t (new_AGEMA_signal_5655), .A1_f (new_AGEMA_signal_5656), .B0_t (RoundKey[44]), .B0_f (new_AGEMA_signal_5657), .B1_t (new_AGEMA_signal_5658), .B1_f (new_AGEMA_signal_5659), .Z0_t (ciphertext_s0_t[44]), .Z0_f (ciphertext_s0_f[44]), .Z1_t (ciphertext_s1_t[44]), .Z1_f (ciphertext_s1_f[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1570 ( .A0_t (RoundInput[45]), .A0_f (new_AGEMA_signal_5663), .A1_t (new_AGEMA_signal_5664), .A1_f (new_AGEMA_signal_5665), .B0_t (RoundKey[45]), .B0_f (new_AGEMA_signal_5666), .B1_t (new_AGEMA_signal_5667), .B1_f (new_AGEMA_signal_5668), .Z0_t (ciphertext_s0_t[45]), .Z0_f (ciphertext_s0_f[45]), .Z1_t (ciphertext_s1_t[45]), .Z1_f (ciphertext_s1_f[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1571 ( .A0_t (RoundInput[46]), .A0_f (new_AGEMA_signal_5672), .A1_t (new_AGEMA_signal_5673), .A1_f (new_AGEMA_signal_5674), .B0_t (RoundKey[46]), .B0_f (new_AGEMA_signal_5675), .B1_t (new_AGEMA_signal_5676), .B1_f (new_AGEMA_signal_5677), .Z0_t (ciphertext_s0_t[46]), .Z0_f (ciphertext_s0_f[46]), .Z1_t (ciphertext_s1_t[46]), .Z1_f (ciphertext_s1_f[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1572 ( .A0_t (RoundInput[47]), .A0_f (new_AGEMA_signal_5681), .A1_t (new_AGEMA_signal_5682), .A1_f (new_AGEMA_signal_5683), .B0_t (RoundKey[47]), .B0_f (new_AGEMA_signal_5684), .B1_t (new_AGEMA_signal_5685), .B1_f (new_AGEMA_signal_5686), .Z0_t (ciphertext_s0_t[47]), .Z0_f (ciphertext_s0_f[47]), .Z1_t (ciphertext_s1_t[47]), .Z1_f (ciphertext_s1_f[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1573 ( .A0_t (RoundInput[48]), .A0_f (new_AGEMA_signal_5690), .A1_t (new_AGEMA_signal_5691), .A1_f (new_AGEMA_signal_5692), .B0_t (RoundKey[48]), .B0_f (new_AGEMA_signal_5693), .B1_t (new_AGEMA_signal_5694), .B1_f (new_AGEMA_signal_5695), .Z0_t (ciphertext_s0_t[48]), .Z0_f (ciphertext_s0_f[48]), .Z1_t (ciphertext_s1_t[48]), .Z1_f (ciphertext_s1_f[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1574 ( .A0_t (RoundInput[49]), .A0_f (new_AGEMA_signal_5699), .A1_t (new_AGEMA_signal_5700), .A1_f (new_AGEMA_signal_5701), .B0_t (RoundKey[49]), .B0_f (new_AGEMA_signal_5702), .B1_t (new_AGEMA_signal_5703), .B1_f (new_AGEMA_signal_5704), .Z0_t (ciphertext_s0_t[49]), .Z0_f (ciphertext_s0_f[49]), .Z1_t (ciphertext_s1_t[49]), .Z1_f (ciphertext_s1_f[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1575 ( .A0_t (RoundInput[4]), .A0_f (new_AGEMA_signal_5708), .A1_t (new_AGEMA_signal_5709), .A1_f (new_AGEMA_signal_5710), .B0_t (RoundKey[4]), .B0_f (new_AGEMA_signal_5711), .B1_t (new_AGEMA_signal_5712), .B1_f (new_AGEMA_signal_5713), .Z0_t (ciphertext_s0_t[4]), .Z0_f (ciphertext_s0_f[4]), .Z1_t (ciphertext_s1_t[4]), .Z1_f (ciphertext_s1_f[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1576 ( .A0_t (RoundInput[50]), .A0_f (new_AGEMA_signal_5717), .A1_t (new_AGEMA_signal_5718), .A1_f (new_AGEMA_signal_5719), .B0_t (RoundKey[50]), .B0_f (new_AGEMA_signal_5720), .B1_t (new_AGEMA_signal_5721), .B1_f (new_AGEMA_signal_5722), .Z0_t (ciphertext_s0_t[50]), .Z0_f (ciphertext_s0_f[50]), .Z1_t (ciphertext_s1_t[50]), .Z1_f (ciphertext_s1_f[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1577 ( .A0_t (RoundInput[51]), .A0_f (new_AGEMA_signal_5726), .A1_t (new_AGEMA_signal_5727), .A1_f (new_AGEMA_signal_5728), .B0_t (RoundKey[51]), .B0_f (new_AGEMA_signal_5729), .B1_t (new_AGEMA_signal_5730), .B1_f (new_AGEMA_signal_5731), .Z0_t (ciphertext_s0_t[51]), .Z0_f (ciphertext_s0_f[51]), .Z1_t (ciphertext_s1_t[51]), .Z1_f (ciphertext_s1_f[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1578 ( .A0_t (RoundInput[52]), .A0_f (new_AGEMA_signal_5735), .A1_t (new_AGEMA_signal_5736), .A1_f (new_AGEMA_signal_5737), .B0_t (RoundKey[52]), .B0_f (new_AGEMA_signal_5738), .B1_t (new_AGEMA_signal_5739), .B1_f (new_AGEMA_signal_5740), .Z0_t (ciphertext_s0_t[52]), .Z0_f (ciphertext_s0_f[52]), .Z1_t (ciphertext_s1_t[52]), .Z1_f (ciphertext_s1_f[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1579 ( .A0_t (RoundInput[53]), .A0_f (new_AGEMA_signal_5744), .A1_t (new_AGEMA_signal_5745), .A1_f (new_AGEMA_signal_5746), .B0_t (RoundKey[53]), .B0_f (new_AGEMA_signal_5747), .B1_t (new_AGEMA_signal_5748), .B1_f (new_AGEMA_signal_5749), .Z0_t (ciphertext_s0_t[53]), .Z0_f (ciphertext_s0_f[53]), .Z1_t (ciphertext_s1_t[53]), .Z1_f (ciphertext_s1_f[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1580 ( .A0_t (RoundInput[54]), .A0_f (new_AGEMA_signal_5753), .A1_t (new_AGEMA_signal_5754), .A1_f (new_AGEMA_signal_5755), .B0_t (RoundKey[54]), .B0_f (new_AGEMA_signal_5756), .B1_t (new_AGEMA_signal_5757), .B1_f (new_AGEMA_signal_5758), .Z0_t (ciphertext_s0_t[54]), .Z0_f (ciphertext_s0_f[54]), .Z1_t (ciphertext_s1_t[54]), .Z1_f (ciphertext_s1_f[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1581 ( .A0_t (RoundInput[55]), .A0_f (new_AGEMA_signal_5762), .A1_t (new_AGEMA_signal_5763), .A1_f (new_AGEMA_signal_5764), .B0_t (RoundKey[55]), .B0_f (new_AGEMA_signal_5765), .B1_t (new_AGEMA_signal_5766), .B1_f (new_AGEMA_signal_5767), .Z0_t (ciphertext_s0_t[55]), .Z0_f (ciphertext_s0_f[55]), .Z1_t (ciphertext_s1_t[55]), .Z1_f (ciphertext_s1_f[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1582 ( .A0_t (RoundInput[56]), .A0_f (new_AGEMA_signal_5771), .A1_t (new_AGEMA_signal_5772), .A1_f (new_AGEMA_signal_5773), .B0_t (RoundKey[56]), .B0_f (new_AGEMA_signal_5774), .B1_t (new_AGEMA_signal_5775), .B1_f (new_AGEMA_signal_5776), .Z0_t (ciphertext_s0_t[56]), .Z0_f (ciphertext_s0_f[56]), .Z1_t (ciphertext_s1_t[56]), .Z1_f (ciphertext_s1_f[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1583 ( .A0_t (RoundInput[57]), .A0_f (new_AGEMA_signal_5780), .A1_t (new_AGEMA_signal_5781), .A1_f (new_AGEMA_signal_5782), .B0_t (RoundKey[57]), .B0_f (new_AGEMA_signal_5783), .B1_t (new_AGEMA_signal_5784), .B1_f (new_AGEMA_signal_5785), .Z0_t (ciphertext_s0_t[57]), .Z0_f (ciphertext_s0_f[57]), .Z1_t (ciphertext_s1_t[57]), .Z1_f (ciphertext_s1_f[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1584 ( .A0_t (RoundInput[58]), .A0_f (new_AGEMA_signal_5789), .A1_t (new_AGEMA_signal_5790), .A1_f (new_AGEMA_signal_5791), .B0_t (RoundKey[58]), .B0_f (new_AGEMA_signal_5792), .B1_t (new_AGEMA_signal_5793), .B1_f (new_AGEMA_signal_5794), .Z0_t (ciphertext_s0_t[58]), .Z0_f (ciphertext_s0_f[58]), .Z1_t (ciphertext_s1_t[58]), .Z1_f (ciphertext_s1_f[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1585 ( .A0_t (RoundInput[59]), .A0_f (new_AGEMA_signal_5798), .A1_t (new_AGEMA_signal_5799), .A1_f (new_AGEMA_signal_5800), .B0_t (RoundKey[59]), .B0_f (new_AGEMA_signal_5801), .B1_t (new_AGEMA_signal_5802), .B1_f (new_AGEMA_signal_5803), .Z0_t (ciphertext_s0_t[59]), .Z0_f (ciphertext_s0_f[59]), .Z1_t (ciphertext_s1_t[59]), .Z1_f (ciphertext_s1_f[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1586 ( .A0_t (RoundInput[5]), .A0_f (new_AGEMA_signal_5807), .A1_t (new_AGEMA_signal_5808), .A1_f (new_AGEMA_signal_5809), .B0_t (RoundKey[5]), .B0_f (new_AGEMA_signal_5810), .B1_t (new_AGEMA_signal_5811), .B1_f (new_AGEMA_signal_5812), .Z0_t (ciphertext_s0_t[5]), .Z0_f (ciphertext_s0_f[5]), .Z1_t (ciphertext_s1_t[5]), .Z1_f (ciphertext_s1_f[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1587 ( .A0_t (RoundInput[60]), .A0_f (new_AGEMA_signal_5816), .A1_t (new_AGEMA_signal_5817), .A1_f (new_AGEMA_signal_5818), .B0_t (RoundKey[60]), .B0_f (new_AGEMA_signal_5819), .B1_t (new_AGEMA_signal_5820), .B1_f (new_AGEMA_signal_5821), .Z0_t (ciphertext_s0_t[60]), .Z0_f (ciphertext_s0_f[60]), .Z1_t (ciphertext_s1_t[60]), .Z1_f (ciphertext_s1_f[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1588 ( .A0_t (RoundInput[61]), .A0_f (new_AGEMA_signal_5825), .A1_t (new_AGEMA_signal_5826), .A1_f (new_AGEMA_signal_5827), .B0_t (RoundKey[61]), .B0_f (new_AGEMA_signal_5828), .B1_t (new_AGEMA_signal_5829), .B1_f (new_AGEMA_signal_5830), .Z0_t (ciphertext_s0_t[61]), .Z0_f (ciphertext_s0_f[61]), .Z1_t (ciphertext_s1_t[61]), .Z1_f (ciphertext_s1_f[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1589 ( .A0_t (RoundInput[62]), .A0_f (new_AGEMA_signal_5834), .A1_t (new_AGEMA_signal_5835), .A1_f (new_AGEMA_signal_5836), .B0_t (RoundKey[62]), .B0_f (new_AGEMA_signal_5837), .B1_t (new_AGEMA_signal_5838), .B1_f (new_AGEMA_signal_5839), .Z0_t (ciphertext_s0_t[62]), .Z0_f (ciphertext_s0_f[62]), .Z1_t (ciphertext_s1_t[62]), .Z1_f (ciphertext_s1_f[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1590 ( .A0_t (RoundInput[63]), .A0_f (new_AGEMA_signal_5843), .A1_t (new_AGEMA_signal_5844), .A1_f (new_AGEMA_signal_5845), .B0_t (RoundKey[63]), .B0_f (new_AGEMA_signal_5846), .B1_t (new_AGEMA_signal_5847), .B1_f (new_AGEMA_signal_5848), .Z0_t (ciphertext_s0_t[63]), .Z0_f (ciphertext_s0_f[63]), .Z1_t (ciphertext_s1_t[63]), .Z1_f (ciphertext_s1_f[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1591 ( .A0_t (RoundInput[64]), .A0_f (new_AGEMA_signal_5852), .A1_t (new_AGEMA_signal_5853), .A1_f (new_AGEMA_signal_5854), .B0_t (RoundKey[64]), .B0_f (new_AGEMA_signal_5855), .B1_t (new_AGEMA_signal_5856), .B1_f (new_AGEMA_signal_5857), .Z0_t (ciphertext_s0_t[64]), .Z0_f (ciphertext_s0_f[64]), .Z1_t (ciphertext_s1_t[64]), .Z1_f (ciphertext_s1_f[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1592 ( .A0_t (RoundInput[65]), .A0_f (new_AGEMA_signal_5861), .A1_t (new_AGEMA_signal_5862), .A1_f (new_AGEMA_signal_5863), .B0_t (RoundKey[65]), .B0_f (new_AGEMA_signal_5864), .B1_t (new_AGEMA_signal_5865), .B1_f (new_AGEMA_signal_5866), .Z0_t (ciphertext_s0_t[65]), .Z0_f (ciphertext_s0_f[65]), .Z1_t (ciphertext_s1_t[65]), .Z1_f (ciphertext_s1_f[65]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1593 ( .A0_t (RoundInput[66]), .A0_f (new_AGEMA_signal_5870), .A1_t (new_AGEMA_signal_5871), .A1_f (new_AGEMA_signal_5872), .B0_t (RoundKey[66]), .B0_f (new_AGEMA_signal_5873), .B1_t (new_AGEMA_signal_5874), .B1_f (new_AGEMA_signal_5875), .Z0_t (ciphertext_s0_t[66]), .Z0_f (ciphertext_s0_f[66]), .Z1_t (ciphertext_s1_t[66]), .Z1_f (ciphertext_s1_f[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1594 ( .A0_t (RoundInput[67]), .A0_f (new_AGEMA_signal_5879), .A1_t (new_AGEMA_signal_5880), .A1_f (new_AGEMA_signal_5881), .B0_t (RoundKey[67]), .B0_f (new_AGEMA_signal_5882), .B1_t (new_AGEMA_signal_5883), .B1_f (new_AGEMA_signal_5884), .Z0_t (ciphertext_s0_t[67]), .Z0_f (ciphertext_s0_f[67]), .Z1_t (ciphertext_s1_t[67]), .Z1_f (ciphertext_s1_f[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1595 ( .A0_t (RoundInput[68]), .A0_f (new_AGEMA_signal_5888), .A1_t (new_AGEMA_signal_5889), .A1_f (new_AGEMA_signal_5890), .B0_t (RoundKey[68]), .B0_f (new_AGEMA_signal_5891), .B1_t (new_AGEMA_signal_5892), .B1_f (new_AGEMA_signal_5893), .Z0_t (ciphertext_s0_t[68]), .Z0_f (ciphertext_s0_f[68]), .Z1_t (ciphertext_s1_t[68]), .Z1_f (ciphertext_s1_f[68]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1596 ( .A0_t (RoundInput[69]), .A0_f (new_AGEMA_signal_5897), .A1_t (new_AGEMA_signal_5898), .A1_f (new_AGEMA_signal_5899), .B0_t (RoundKey[69]), .B0_f (new_AGEMA_signal_5900), .B1_t (new_AGEMA_signal_5901), .B1_f (new_AGEMA_signal_5902), .Z0_t (ciphertext_s0_t[69]), .Z0_f (ciphertext_s0_f[69]), .Z1_t (ciphertext_s1_t[69]), .Z1_f (ciphertext_s1_f[69]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1597 ( .A0_t (RoundInput[6]), .A0_f (new_AGEMA_signal_5906), .A1_t (new_AGEMA_signal_5907), .A1_f (new_AGEMA_signal_5908), .B0_t (RoundKey[6]), .B0_f (new_AGEMA_signal_5909), .B1_t (new_AGEMA_signal_5910), .B1_f (new_AGEMA_signal_5911), .Z0_t (ciphertext_s0_t[6]), .Z0_f (ciphertext_s0_f[6]), .Z1_t (ciphertext_s1_t[6]), .Z1_f (ciphertext_s1_f[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1598 ( .A0_t (RoundInput[70]), .A0_f (new_AGEMA_signal_5915), .A1_t (new_AGEMA_signal_5916), .A1_f (new_AGEMA_signal_5917), .B0_t (RoundKey[70]), .B0_f (new_AGEMA_signal_5918), .B1_t (new_AGEMA_signal_5919), .B1_f (new_AGEMA_signal_5920), .Z0_t (ciphertext_s0_t[70]), .Z0_f (ciphertext_s0_f[70]), .Z1_t (ciphertext_s1_t[70]), .Z1_f (ciphertext_s1_f[70]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1599 ( .A0_t (RoundInput[71]), .A0_f (new_AGEMA_signal_5924), .A1_t (new_AGEMA_signal_5925), .A1_f (new_AGEMA_signal_5926), .B0_t (RoundKey[71]), .B0_f (new_AGEMA_signal_5927), .B1_t (new_AGEMA_signal_5928), .B1_f (new_AGEMA_signal_5929), .Z0_t (ciphertext_s0_t[71]), .Z0_f (ciphertext_s0_f[71]), .Z1_t (ciphertext_s1_t[71]), .Z1_f (ciphertext_s1_f[71]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1600 ( .A0_t (RoundInput[72]), .A0_f (new_AGEMA_signal_5933), .A1_t (new_AGEMA_signal_5934), .A1_f (new_AGEMA_signal_5935), .B0_t (RoundKey[72]), .B0_f (new_AGEMA_signal_5936), .B1_t (new_AGEMA_signal_5937), .B1_f (new_AGEMA_signal_5938), .Z0_t (ciphertext_s0_t[72]), .Z0_f (ciphertext_s0_f[72]), .Z1_t (ciphertext_s1_t[72]), .Z1_f (ciphertext_s1_f[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1601 ( .A0_t (RoundInput[73]), .A0_f (new_AGEMA_signal_5942), .A1_t (new_AGEMA_signal_5943), .A1_f (new_AGEMA_signal_5944), .B0_t (RoundKey[73]), .B0_f (new_AGEMA_signal_5945), .B1_t (new_AGEMA_signal_5946), .B1_f (new_AGEMA_signal_5947), .Z0_t (ciphertext_s0_t[73]), .Z0_f (ciphertext_s0_f[73]), .Z1_t (ciphertext_s1_t[73]), .Z1_f (ciphertext_s1_f[73]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1602 ( .A0_t (RoundInput[74]), .A0_f (new_AGEMA_signal_5951), .A1_t (new_AGEMA_signal_5952), .A1_f (new_AGEMA_signal_5953), .B0_t (RoundKey[74]), .B0_f (new_AGEMA_signal_5954), .B1_t (new_AGEMA_signal_5955), .B1_f (new_AGEMA_signal_5956), .Z0_t (ciphertext_s0_t[74]), .Z0_f (ciphertext_s0_f[74]), .Z1_t (ciphertext_s1_t[74]), .Z1_f (ciphertext_s1_f[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1603 ( .A0_t (RoundInput[75]), .A0_f (new_AGEMA_signal_5960), .A1_t (new_AGEMA_signal_5961), .A1_f (new_AGEMA_signal_5962), .B0_t (RoundKey[75]), .B0_f (new_AGEMA_signal_5963), .B1_t (new_AGEMA_signal_5964), .B1_f (new_AGEMA_signal_5965), .Z0_t (ciphertext_s0_t[75]), .Z0_f (ciphertext_s0_f[75]), .Z1_t (ciphertext_s1_t[75]), .Z1_f (ciphertext_s1_f[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1604 ( .A0_t (RoundInput[76]), .A0_f (new_AGEMA_signal_5969), .A1_t (new_AGEMA_signal_5970), .A1_f (new_AGEMA_signal_5971), .B0_t (RoundKey[76]), .B0_f (new_AGEMA_signal_5972), .B1_t (new_AGEMA_signal_5973), .B1_f (new_AGEMA_signal_5974), .Z0_t (ciphertext_s0_t[76]), .Z0_f (ciphertext_s0_f[76]), .Z1_t (ciphertext_s1_t[76]), .Z1_f (ciphertext_s1_f[76]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1605 ( .A0_t (RoundInput[77]), .A0_f (new_AGEMA_signal_5978), .A1_t (new_AGEMA_signal_5979), .A1_f (new_AGEMA_signal_5980), .B0_t (RoundKey[77]), .B0_f (new_AGEMA_signal_5981), .B1_t (new_AGEMA_signal_5982), .B1_f (new_AGEMA_signal_5983), .Z0_t (ciphertext_s0_t[77]), .Z0_f (ciphertext_s0_f[77]), .Z1_t (ciphertext_s1_t[77]), .Z1_f (ciphertext_s1_f[77]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1606 ( .A0_t (RoundInput[78]), .A0_f (new_AGEMA_signal_5987), .A1_t (new_AGEMA_signal_5988), .A1_f (new_AGEMA_signal_5989), .B0_t (RoundKey[78]), .B0_f (new_AGEMA_signal_5990), .B1_t (new_AGEMA_signal_5991), .B1_f (new_AGEMA_signal_5992), .Z0_t (ciphertext_s0_t[78]), .Z0_f (ciphertext_s0_f[78]), .Z1_t (ciphertext_s1_t[78]), .Z1_f (ciphertext_s1_f[78]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1607 ( .A0_t (RoundInput[79]), .A0_f (new_AGEMA_signal_5996), .A1_t (new_AGEMA_signal_5997), .A1_f (new_AGEMA_signal_5998), .B0_t (RoundKey[79]), .B0_f (new_AGEMA_signal_5999), .B1_t (new_AGEMA_signal_6000), .B1_f (new_AGEMA_signal_6001), .Z0_t (ciphertext_s0_t[79]), .Z0_f (ciphertext_s0_f[79]), .Z1_t (ciphertext_s1_t[79]), .Z1_f (ciphertext_s1_f[79]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1608 ( .A0_t (RoundInput[7]), .A0_f (new_AGEMA_signal_6005), .A1_t (new_AGEMA_signal_6006), .A1_f (new_AGEMA_signal_6007), .B0_t (RoundKey[7]), .B0_f (new_AGEMA_signal_6008), .B1_t (new_AGEMA_signal_6009), .B1_f (new_AGEMA_signal_6010), .Z0_t (ciphertext_s0_t[7]), .Z0_f (ciphertext_s0_f[7]), .Z1_t (ciphertext_s1_t[7]), .Z1_f (ciphertext_s1_f[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1609 ( .A0_t (RoundInput[80]), .A0_f (new_AGEMA_signal_6014), .A1_t (new_AGEMA_signal_6015), .A1_f (new_AGEMA_signal_6016), .B0_t (RoundKey[80]), .B0_f (new_AGEMA_signal_6017), .B1_t (new_AGEMA_signal_6018), .B1_f (new_AGEMA_signal_6019), .Z0_t (ciphertext_s0_t[80]), .Z0_f (ciphertext_s0_f[80]), .Z1_t (ciphertext_s1_t[80]), .Z1_f (ciphertext_s1_f[80]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1610 ( .A0_t (RoundInput[81]), .A0_f (new_AGEMA_signal_6023), .A1_t (new_AGEMA_signal_6024), .A1_f (new_AGEMA_signal_6025), .B0_t (RoundKey[81]), .B0_f (new_AGEMA_signal_6026), .B1_t (new_AGEMA_signal_6027), .B1_f (new_AGEMA_signal_6028), .Z0_t (ciphertext_s0_t[81]), .Z0_f (ciphertext_s0_f[81]), .Z1_t (ciphertext_s1_t[81]), .Z1_f (ciphertext_s1_f[81]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1611 ( .A0_t (RoundInput[82]), .A0_f (new_AGEMA_signal_6032), .A1_t (new_AGEMA_signal_6033), .A1_f (new_AGEMA_signal_6034), .B0_t (RoundKey[82]), .B0_f (new_AGEMA_signal_6035), .B1_t (new_AGEMA_signal_6036), .B1_f (new_AGEMA_signal_6037), .Z0_t (ciphertext_s0_t[82]), .Z0_f (ciphertext_s0_f[82]), .Z1_t (ciphertext_s1_t[82]), .Z1_f (ciphertext_s1_f[82]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1612 ( .A0_t (RoundInput[83]), .A0_f (new_AGEMA_signal_6041), .A1_t (new_AGEMA_signal_6042), .A1_f (new_AGEMA_signal_6043), .B0_t (RoundKey[83]), .B0_f (new_AGEMA_signal_6044), .B1_t (new_AGEMA_signal_6045), .B1_f (new_AGEMA_signal_6046), .Z0_t (ciphertext_s0_t[83]), .Z0_f (ciphertext_s0_f[83]), .Z1_t (ciphertext_s1_t[83]), .Z1_f (ciphertext_s1_f[83]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1613 ( .A0_t (RoundInput[84]), .A0_f (new_AGEMA_signal_6050), .A1_t (new_AGEMA_signal_6051), .A1_f (new_AGEMA_signal_6052), .B0_t (RoundKey[84]), .B0_f (new_AGEMA_signal_6053), .B1_t (new_AGEMA_signal_6054), .B1_f (new_AGEMA_signal_6055), .Z0_t (ciphertext_s0_t[84]), .Z0_f (ciphertext_s0_f[84]), .Z1_t (ciphertext_s1_t[84]), .Z1_f (ciphertext_s1_f[84]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1614 ( .A0_t (RoundInput[85]), .A0_f (new_AGEMA_signal_6059), .A1_t (new_AGEMA_signal_6060), .A1_f (new_AGEMA_signal_6061), .B0_t (RoundKey[85]), .B0_f (new_AGEMA_signal_6062), .B1_t (new_AGEMA_signal_6063), .B1_f (new_AGEMA_signal_6064), .Z0_t (ciphertext_s0_t[85]), .Z0_f (ciphertext_s0_f[85]), .Z1_t (ciphertext_s1_t[85]), .Z1_f (ciphertext_s1_f[85]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1615 ( .A0_t (RoundInput[86]), .A0_f (new_AGEMA_signal_6068), .A1_t (new_AGEMA_signal_6069), .A1_f (new_AGEMA_signal_6070), .B0_t (RoundKey[86]), .B0_f (new_AGEMA_signal_6071), .B1_t (new_AGEMA_signal_6072), .B1_f (new_AGEMA_signal_6073), .Z0_t (ciphertext_s0_t[86]), .Z0_f (ciphertext_s0_f[86]), .Z1_t (ciphertext_s1_t[86]), .Z1_f (ciphertext_s1_f[86]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1616 ( .A0_t (RoundInput[87]), .A0_f (new_AGEMA_signal_6077), .A1_t (new_AGEMA_signal_6078), .A1_f (new_AGEMA_signal_6079), .B0_t (RoundKey[87]), .B0_f (new_AGEMA_signal_6080), .B1_t (new_AGEMA_signal_6081), .B1_f (new_AGEMA_signal_6082), .Z0_t (ciphertext_s0_t[87]), .Z0_f (ciphertext_s0_f[87]), .Z1_t (ciphertext_s1_t[87]), .Z1_f (ciphertext_s1_f[87]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1617 ( .A0_t (RoundInput[88]), .A0_f (new_AGEMA_signal_6086), .A1_t (new_AGEMA_signal_6087), .A1_f (new_AGEMA_signal_6088), .B0_t (RoundKey[88]), .B0_f (new_AGEMA_signal_6089), .B1_t (new_AGEMA_signal_6090), .B1_f (new_AGEMA_signal_6091), .Z0_t (ciphertext_s0_t[88]), .Z0_f (ciphertext_s0_f[88]), .Z1_t (ciphertext_s1_t[88]), .Z1_f (ciphertext_s1_f[88]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1618 ( .A0_t (RoundInput[89]), .A0_f (new_AGEMA_signal_6095), .A1_t (new_AGEMA_signal_6096), .A1_f (new_AGEMA_signal_6097), .B0_t (RoundKey[89]), .B0_f (new_AGEMA_signal_6098), .B1_t (new_AGEMA_signal_6099), .B1_f (new_AGEMA_signal_6100), .Z0_t (ciphertext_s0_t[89]), .Z0_f (ciphertext_s0_f[89]), .Z1_t (ciphertext_s1_t[89]), .Z1_f (ciphertext_s1_f[89]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1619 ( .A0_t (RoundInput[8]), .A0_f (new_AGEMA_signal_6104), .A1_t (new_AGEMA_signal_6105), .A1_f (new_AGEMA_signal_6106), .B0_t (RoundKey[8]), .B0_f (new_AGEMA_signal_6107), .B1_t (new_AGEMA_signal_6108), .B1_f (new_AGEMA_signal_6109), .Z0_t (ciphertext_s0_t[8]), .Z0_f (ciphertext_s0_f[8]), .Z1_t (ciphertext_s1_t[8]), .Z1_f (ciphertext_s1_f[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1620 ( .A0_t (RoundInput[90]), .A0_f (new_AGEMA_signal_6113), .A1_t (new_AGEMA_signal_6114), .A1_f (new_AGEMA_signal_6115), .B0_t (RoundKey[90]), .B0_f (new_AGEMA_signal_6116), .B1_t (new_AGEMA_signal_6117), .B1_f (new_AGEMA_signal_6118), .Z0_t (ciphertext_s0_t[90]), .Z0_f (ciphertext_s0_f[90]), .Z1_t (ciphertext_s1_t[90]), .Z1_f (ciphertext_s1_f[90]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1621 ( .A0_t (RoundInput[91]), .A0_f (new_AGEMA_signal_6122), .A1_t (new_AGEMA_signal_6123), .A1_f (new_AGEMA_signal_6124), .B0_t (RoundKey[91]), .B0_f (new_AGEMA_signal_6125), .B1_t (new_AGEMA_signal_6126), .B1_f (new_AGEMA_signal_6127), .Z0_t (ciphertext_s0_t[91]), .Z0_f (ciphertext_s0_f[91]), .Z1_t (ciphertext_s1_t[91]), .Z1_f (ciphertext_s1_f[91]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1622 ( .A0_t (RoundInput[92]), .A0_f (new_AGEMA_signal_6131), .A1_t (new_AGEMA_signal_6132), .A1_f (new_AGEMA_signal_6133), .B0_t (RoundKey[92]), .B0_f (new_AGEMA_signal_6134), .B1_t (new_AGEMA_signal_6135), .B1_f (new_AGEMA_signal_6136), .Z0_t (ciphertext_s0_t[92]), .Z0_f (ciphertext_s0_f[92]), .Z1_t (ciphertext_s1_t[92]), .Z1_f (ciphertext_s1_f[92]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1623 ( .A0_t (RoundInput[93]), .A0_f (new_AGEMA_signal_6140), .A1_t (new_AGEMA_signal_6141), .A1_f (new_AGEMA_signal_6142), .B0_t (RoundKey[93]), .B0_f (new_AGEMA_signal_6143), .B1_t (new_AGEMA_signal_6144), .B1_f (new_AGEMA_signal_6145), .Z0_t (ciphertext_s0_t[93]), .Z0_f (ciphertext_s0_f[93]), .Z1_t (ciphertext_s1_t[93]), .Z1_f (ciphertext_s1_f[93]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1624 ( .A0_t (RoundInput[94]), .A0_f (new_AGEMA_signal_6149), .A1_t (new_AGEMA_signal_6150), .A1_f (new_AGEMA_signal_6151), .B0_t (RoundKey[94]), .B0_f (new_AGEMA_signal_6152), .B1_t (new_AGEMA_signal_6153), .B1_f (new_AGEMA_signal_6154), .Z0_t (ciphertext_s0_t[94]), .Z0_f (ciphertext_s0_f[94]), .Z1_t (ciphertext_s1_t[94]), .Z1_f (ciphertext_s1_f[94]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1625 ( .A0_t (RoundInput[95]), .A0_f (new_AGEMA_signal_6158), .A1_t (new_AGEMA_signal_6159), .A1_f (new_AGEMA_signal_6160), .B0_t (RoundKey[95]), .B0_f (new_AGEMA_signal_6161), .B1_t (new_AGEMA_signal_6162), .B1_f (new_AGEMA_signal_6163), .Z0_t (ciphertext_s0_t[95]), .Z0_f (ciphertext_s0_f[95]), .Z1_t (ciphertext_s1_t[95]), .Z1_f (ciphertext_s1_f[95]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1626 ( .A0_t (RoundInput[96]), .A0_f (new_AGEMA_signal_6167), .A1_t (new_AGEMA_signal_6168), .A1_f (new_AGEMA_signal_6169), .B0_t (RoundKey[96]), .B0_f (new_AGEMA_signal_6170), .B1_t (new_AGEMA_signal_6171), .B1_f (new_AGEMA_signal_6172), .Z0_t (ciphertext_s0_t[96]), .Z0_f (ciphertext_s0_f[96]), .Z1_t (ciphertext_s1_t[96]), .Z1_f (ciphertext_s1_f[96]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1627 ( .A0_t (RoundInput[97]), .A0_f (new_AGEMA_signal_6176), .A1_t (new_AGEMA_signal_6177), .A1_f (new_AGEMA_signal_6178), .B0_t (RoundKey[97]), .B0_f (new_AGEMA_signal_6179), .B1_t (new_AGEMA_signal_6180), .B1_f (new_AGEMA_signal_6181), .Z0_t (ciphertext_s0_t[97]), .Z0_f (ciphertext_s0_f[97]), .Z1_t (ciphertext_s1_t[97]), .Z1_f (ciphertext_s1_f[97]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1628 ( .A0_t (RoundInput[98]), .A0_f (new_AGEMA_signal_6185), .A1_t (new_AGEMA_signal_6186), .A1_f (new_AGEMA_signal_6187), .B0_t (RoundKey[98]), .B0_f (new_AGEMA_signal_6188), .B1_t (new_AGEMA_signal_6189), .B1_f (new_AGEMA_signal_6190), .Z0_t (ciphertext_s0_t[98]), .Z0_f (ciphertext_s0_f[98]), .Z1_t (ciphertext_s1_t[98]), .Z1_f (ciphertext_s1_f[98]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1629 ( .A0_t (RoundInput[99]), .A0_f (new_AGEMA_signal_6194), .A1_t (new_AGEMA_signal_6195), .A1_f (new_AGEMA_signal_6196), .B0_t (RoundKey[99]), .B0_f (new_AGEMA_signal_6197), .B1_t (new_AGEMA_signal_6198), .B1_f (new_AGEMA_signal_6199), .Z0_t (ciphertext_s0_t[99]), .Z0_f (ciphertext_s0_f[99]), .Z1_t (ciphertext_s1_t[99]), .Z1_f (ciphertext_s1_f[99]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1630 ( .A0_t (RoundInput[9]), .A0_f (new_AGEMA_signal_6203), .A1_t (new_AGEMA_signal_6204), .A1_f (new_AGEMA_signal_6205), .B0_t (RoundKey[9]), .B0_f (new_AGEMA_signal_6206), .B1_t (new_AGEMA_signal_6207), .B1_f (new_AGEMA_signal_6208), .Z0_t (ciphertext_s0_t[9]), .Z0_f (ciphertext_s0_f[9]), .Z1_t (ciphertext_s1_t[9]), .Z1_f (ciphertext_s1_f[9]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1631 ( .A0_t (RoundCounter[3]), .A0_f (new_AGEMA_signal_5055), .B0_t (n851), .B0_f (new_AGEMA_signal_5057), .Z0_t (n852), .Z0_f (new_AGEMA_signal_6343) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1632 ( .A0_t (RoundCounter[0]), .A0_f (new_AGEMA_signal_5054), .B0_t (n852), .B0_f (new_AGEMA_signal_6343), .Z0_t (done_t), .Z0_f (done_f) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1634 ( .A0_t (RoundCounter[1]), .A0_f (new_AGEMA_signal_5051), .B0_t (RoundCounter[2]), .B0_f (new_AGEMA_signal_5052), .Z0_t (n856), .Z0_f (new_AGEMA_signal_6212) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1635 ( .A0_t (n853), .A0_f (new_AGEMA_signal_5058), .B0_t (n856), .B0_f (new_AGEMA_signal_6212), .Z0_t (n283), .Z0_f (new_AGEMA_signal_6344) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1637 ( .A0_t (n855), .A0_f (new_AGEMA_signal_5056), .B0_t (n856), .B0_f (new_AGEMA_signal_6212), .Z0_t (n285), .Z0_f (new_AGEMA_signal_6345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_0_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[0]), .A0_f (new_AGEMA_signal_17246), .A1_t (new_AGEMA_signal_17247), .A1_f (new_AGEMA_signal_17248), .B0_t (plaintext_s0_t[0]), .B0_f (plaintext_s0_f[0]), .B1_t (plaintext_s1_t[0]), .B1_f (plaintext_s1_f[0]), .Z0_t (RoundReg_Inst_ff_SDE_0_MUX_inst_X), .Z0_f (new_AGEMA_signal_17906), .Z1_t (new_AGEMA_signal_17907), .Z1_f (new_AGEMA_signal_17908) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_0_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_0_MUX_inst_X), .B0_f (new_AGEMA_signal_17906), .B1_t (new_AGEMA_signal_17907), .B1_f (new_AGEMA_signal_17908), .Z0_t (RoundReg_Inst_ff_SDE_0_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18404), .Z1_t (new_AGEMA_signal_18405), .Z1_f (new_AGEMA_signal_18406) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_0_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_0_MUX_inst_Y), .A0_f (new_AGEMA_signal_18404), .A1_t (new_AGEMA_signal_18405), .A1_f (new_AGEMA_signal_18406), .B0_t (RoundOutput[0]), .B0_f (new_AGEMA_signal_17246), .B1_t (new_AGEMA_signal_17247), .B1_f (new_AGEMA_signal_17248), .Z0_t (RoundInput[0]), .Z0_f (new_AGEMA_signal_5060), .Z1_t (new_AGEMA_signal_5061), .Z1_f (new_AGEMA_signal_5062) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_1_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[1]), .A0_f (new_AGEMA_signal_17801), .A1_t (new_AGEMA_signal_17802), .A1_f (new_AGEMA_signal_17803), .B0_t (plaintext_s0_t[1]), .B0_f (plaintext_s0_f[1]), .B1_t (plaintext_s1_t[1]), .B1_f (plaintext_s1_f[1]), .Z0_t (RoundReg_Inst_ff_SDE_1_MUX_inst_X), .Z0_f (new_AGEMA_signal_18410), .Z1_t (new_AGEMA_signal_18411), .Z1_f (new_AGEMA_signal_18412) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_1_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_1_MUX_inst_X), .B0_f (new_AGEMA_signal_18410), .B1_t (new_AGEMA_signal_18411), .B1_f (new_AGEMA_signal_18412), .Z0_t (RoundReg_Inst_ff_SDE_1_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18932), .Z1_t (new_AGEMA_signal_18933), .Z1_f (new_AGEMA_signal_18934) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_1_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_1_MUX_inst_Y), .A0_f (new_AGEMA_signal_18932), .A1_t (new_AGEMA_signal_18933), .A1_f (new_AGEMA_signal_18934), .B0_t (RoundOutput[1]), .B0_f (new_AGEMA_signal_17801), .B1_t (new_AGEMA_signal_17802), .B1_f (new_AGEMA_signal_17803), .Z0_t (RoundInput[1]), .Z0_f (new_AGEMA_signal_5411), .Z1_t (new_AGEMA_signal_5412), .Z1_f (new_AGEMA_signal_5413) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_2_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[2]), .A0_f (new_AGEMA_signal_17396), .A1_t (new_AGEMA_signal_17397), .A1_f (new_AGEMA_signal_17398), .B0_t (plaintext_s0_t[2]), .B0_f (plaintext_s0_f[2]), .B1_t (plaintext_s1_t[2]), .B1_f (plaintext_s1_f[2]), .Z0_t (RoundReg_Inst_ff_SDE_2_MUX_inst_X), .Z0_f (new_AGEMA_signal_17912), .Z1_t (new_AGEMA_signal_17913), .Z1_f (new_AGEMA_signal_17914) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_2_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_2_MUX_inst_X), .B0_f (new_AGEMA_signal_17912), .B1_t (new_AGEMA_signal_17913), .B1_f (new_AGEMA_signal_17914), .Z0_t (RoundReg_Inst_ff_SDE_2_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18413), .Z1_t (new_AGEMA_signal_18414), .Z1_f (new_AGEMA_signal_18415) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_2_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_2_MUX_inst_Y), .A0_f (new_AGEMA_signal_18413), .A1_t (new_AGEMA_signal_18414), .A1_f (new_AGEMA_signal_18415), .B0_t (RoundOutput[2]), .B0_f (new_AGEMA_signal_17396), .B1_t (new_AGEMA_signal_17397), .B1_f (new_AGEMA_signal_17398), .Z0_t (RoundInput[2]), .Z0_f (new_AGEMA_signal_5510), .Z1_t (new_AGEMA_signal_5511), .Z1_f (new_AGEMA_signal_5512) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_3_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[3]), .A0_f (new_AGEMA_signal_17825), .A1_t (new_AGEMA_signal_17826), .A1_f (new_AGEMA_signal_17827), .B0_t (plaintext_s0_t[3]), .B0_f (plaintext_s0_f[3]), .B1_t (plaintext_s1_t[3]), .B1_f (plaintext_s1_f[3]), .Z0_t (RoundReg_Inst_ff_SDE_3_MUX_inst_X), .Z0_f (new_AGEMA_signal_18419), .Z1_t (new_AGEMA_signal_18420), .Z1_f (new_AGEMA_signal_18421) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_3_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_3_MUX_inst_X), .B0_f (new_AGEMA_signal_18419), .B1_t (new_AGEMA_signal_18420), .B1_f (new_AGEMA_signal_18421), .Z0_t (RoundReg_Inst_ff_SDE_3_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18935), .Z1_t (new_AGEMA_signal_18936), .Z1_f (new_AGEMA_signal_18937) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_3_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_3_MUX_inst_Y), .A0_f (new_AGEMA_signal_18935), .A1_t (new_AGEMA_signal_18936), .A1_f (new_AGEMA_signal_18937), .B0_t (RoundOutput[3]), .B0_f (new_AGEMA_signal_17825), .B1_t (new_AGEMA_signal_17826), .B1_f (new_AGEMA_signal_17827), .Z0_t (RoundInput[3]), .Z0_f (new_AGEMA_signal_5609), .Z1_t (new_AGEMA_signal_5610), .Z1_f (new_AGEMA_signal_5611) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_4_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[4]), .A0_f (new_AGEMA_signal_17840), .A1_t (new_AGEMA_signal_17841), .A1_f (new_AGEMA_signal_17842), .B0_t (plaintext_s0_t[4]), .B0_f (plaintext_s0_f[4]), .B1_t (plaintext_s1_t[4]), .B1_f (plaintext_s1_f[4]), .Z0_t (RoundReg_Inst_ff_SDE_4_MUX_inst_X), .Z0_f (new_AGEMA_signal_18425), .Z1_t (new_AGEMA_signal_18426), .Z1_f (new_AGEMA_signal_18427) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_4_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_4_MUX_inst_X), .B0_f (new_AGEMA_signal_18425), .B1_t (new_AGEMA_signal_18426), .B1_f (new_AGEMA_signal_18427), .Z0_t (RoundReg_Inst_ff_SDE_4_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18938), .Z1_t (new_AGEMA_signal_18939), .Z1_f (new_AGEMA_signal_18940) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_4_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_4_MUX_inst_Y), .A0_f (new_AGEMA_signal_18938), .A1_t (new_AGEMA_signal_18939), .A1_f (new_AGEMA_signal_18940), .B0_t (RoundOutput[4]), .B0_f (new_AGEMA_signal_17840), .B1_t (new_AGEMA_signal_17841), .B1_f (new_AGEMA_signal_17842), .Z0_t (RoundInput[4]), .Z0_f (new_AGEMA_signal_5708), .Z1_t (new_AGEMA_signal_5709), .Z1_f (new_AGEMA_signal_5710) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_5_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[5]), .A0_f (new_AGEMA_signal_17495), .A1_t (new_AGEMA_signal_17496), .A1_f (new_AGEMA_signal_17497), .B0_t (plaintext_s0_t[5]), .B0_f (plaintext_s0_f[5]), .B1_t (plaintext_s1_t[5]), .B1_f (plaintext_s1_f[5]), .Z0_t (RoundReg_Inst_ff_SDE_5_MUX_inst_X), .Z0_f (new_AGEMA_signal_17918), .Z1_t (new_AGEMA_signal_17919), .Z1_f (new_AGEMA_signal_17920) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_5_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_5_MUX_inst_X), .B0_f (new_AGEMA_signal_17918), .B1_t (new_AGEMA_signal_17919), .B1_f (new_AGEMA_signal_17920), .Z0_t (RoundReg_Inst_ff_SDE_5_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18428), .Z1_t (new_AGEMA_signal_18429), .Z1_f (new_AGEMA_signal_18430) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_5_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_5_MUX_inst_Y), .A0_f (new_AGEMA_signal_18428), .A1_t (new_AGEMA_signal_18429), .A1_f (new_AGEMA_signal_18430), .B0_t (RoundOutput[5]), .B0_f (new_AGEMA_signal_17495), .B1_t (new_AGEMA_signal_17496), .B1_f (new_AGEMA_signal_17497), .Z0_t (RoundInput[5]), .Z0_f (new_AGEMA_signal_5807), .Z1_t (new_AGEMA_signal_5808), .Z1_f (new_AGEMA_signal_5809) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_6_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[6]), .A0_f (new_AGEMA_signal_17528), .A1_t (new_AGEMA_signal_17529), .A1_f (new_AGEMA_signal_17530), .B0_t (plaintext_s0_t[6]), .B0_f (plaintext_s0_f[6]), .B1_t (plaintext_s1_t[6]), .B1_f (plaintext_s1_f[6]), .Z0_t (RoundReg_Inst_ff_SDE_6_MUX_inst_X), .Z0_f (new_AGEMA_signal_17924), .Z1_t (new_AGEMA_signal_17925), .Z1_f (new_AGEMA_signal_17926) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_6_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_6_MUX_inst_X), .B0_f (new_AGEMA_signal_17924), .B1_t (new_AGEMA_signal_17925), .B1_f (new_AGEMA_signal_17926), .Z0_t (RoundReg_Inst_ff_SDE_6_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18431), .Z1_t (new_AGEMA_signal_18432), .Z1_f (new_AGEMA_signal_18433) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_6_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_6_MUX_inst_Y), .A0_f (new_AGEMA_signal_18431), .A1_t (new_AGEMA_signal_18432), .A1_f (new_AGEMA_signal_18433), .B0_t (RoundOutput[6]), .B0_f (new_AGEMA_signal_17528), .B1_t (new_AGEMA_signal_17529), .B1_f (new_AGEMA_signal_17530), .Z0_t (RoundInput[6]), .Z0_f (new_AGEMA_signal_5906), .Z1_t (new_AGEMA_signal_5907), .Z1_f (new_AGEMA_signal_5908) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_7_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[7]), .A0_f (new_AGEMA_signal_17561), .A1_t (new_AGEMA_signal_17562), .A1_f (new_AGEMA_signal_17563), .B0_t (plaintext_s0_t[7]), .B0_f (plaintext_s0_f[7]), .B1_t (plaintext_s1_t[7]), .B1_f (plaintext_s1_f[7]), .Z0_t (RoundReg_Inst_ff_SDE_7_MUX_inst_X), .Z0_f (new_AGEMA_signal_17930), .Z1_t (new_AGEMA_signal_17931), .Z1_f (new_AGEMA_signal_17932) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_7_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_7_MUX_inst_X), .B0_f (new_AGEMA_signal_17930), .B1_t (new_AGEMA_signal_17931), .B1_f (new_AGEMA_signal_17932), .Z0_t (RoundReg_Inst_ff_SDE_7_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18434), .Z1_t (new_AGEMA_signal_18435), .Z1_f (new_AGEMA_signal_18436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_7_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_7_MUX_inst_Y), .A0_f (new_AGEMA_signal_18434), .A1_t (new_AGEMA_signal_18435), .A1_f (new_AGEMA_signal_18436), .B0_t (RoundOutput[7]), .B0_f (new_AGEMA_signal_17561), .B1_t (new_AGEMA_signal_17562), .B1_f (new_AGEMA_signal_17563), .Z0_t (RoundInput[7]), .Z0_f (new_AGEMA_signal_6005), .Z1_t (new_AGEMA_signal_6006), .Z1_f (new_AGEMA_signal_6007) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_8_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[8]), .A0_f (new_AGEMA_signal_17594), .A1_t (new_AGEMA_signal_17595), .A1_f (new_AGEMA_signal_17596), .B0_t (plaintext_s0_t[8]), .B0_f (plaintext_s0_f[8]), .B1_t (plaintext_s1_t[8]), .B1_f (plaintext_s1_f[8]), .Z0_t (RoundReg_Inst_ff_SDE_8_MUX_inst_X), .Z0_f (new_AGEMA_signal_17936), .Z1_t (new_AGEMA_signal_17937), .Z1_f (new_AGEMA_signal_17938) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_8_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_8_MUX_inst_X), .B0_f (new_AGEMA_signal_17936), .B1_t (new_AGEMA_signal_17937), .B1_f (new_AGEMA_signal_17938), .Z0_t (RoundReg_Inst_ff_SDE_8_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18437), .Z1_t (new_AGEMA_signal_18438), .Z1_f (new_AGEMA_signal_18439) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_8_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_8_MUX_inst_Y), .A0_f (new_AGEMA_signal_18437), .A1_t (new_AGEMA_signal_18438), .A1_f (new_AGEMA_signal_18439), .B0_t (RoundOutput[8]), .B0_f (new_AGEMA_signal_17594), .B1_t (new_AGEMA_signal_17595), .B1_f (new_AGEMA_signal_17596), .Z0_t (RoundInput[8]), .Z0_f (new_AGEMA_signal_6104), .Z1_t (new_AGEMA_signal_6105), .Z1_f (new_AGEMA_signal_6106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_9_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[9]), .A0_f (new_AGEMA_signal_17900), .A1_t (new_AGEMA_signal_17901), .A1_f (new_AGEMA_signal_17902), .B0_t (plaintext_s0_t[9]), .B0_f (plaintext_s0_f[9]), .B1_t (plaintext_s1_t[9]), .B1_f (plaintext_s1_f[9]), .Z0_t (RoundReg_Inst_ff_SDE_9_MUX_inst_X), .Z0_f (new_AGEMA_signal_18443), .Z1_t (new_AGEMA_signal_18444), .Z1_f (new_AGEMA_signal_18445) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_9_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_9_MUX_inst_X), .B0_f (new_AGEMA_signal_18443), .B1_t (new_AGEMA_signal_18444), .B1_f (new_AGEMA_signal_18445), .Z0_t (RoundReg_Inst_ff_SDE_9_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18941), .Z1_t (new_AGEMA_signal_18942), .Z1_f (new_AGEMA_signal_18943) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_9_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_9_MUX_inst_Y), .A0_f (new_AGEMA_signal_18941), .A1_t (new_AGEMA_signal_18942), .A1_f (new_AGEMA_signal_18943), .B0_t (RoundOutput[9]), .B0_f (new_AGEMA_signal_17900), .B1_t (new_AGEMA_signal_17901), .B1_f (new_AGEMA_signal_17902), .Z0_t (RoundInput[9]), .Z0_f (new_AGEMA_signal_6203), .Z1_t (new_AGEMA_signal_6204), .Z1_f (new_AGEMA_signal_6205) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_10_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[10]), .A0_f (new_AGEMA_signal_17279), .A1_t (new_AGEMA_signal_17280), .A1_f (new_AGEMA_signal_17281), .B0_t (plaintext_s0_t[10]), .B0_f (plaintext_s0_f[10]), .B1_t (plaintext_s1_t[10]), .B1_f (plaintext_s1_f[10]), .Z0_t (RoundReg_Inst_ff_SDE_10_MUX_inst_X), .Z0_f (new_AGEMA_signal_17942), .Z1_t (new_AGEMA_signal_17943), .Z1_f (new_AGEMA_signal_17944) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_10_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_10_MUX_inst_X), .B0_f (new_AGEMA_signal_17942), .B1_t (new_AGEMA_signal_17943), .B1_f (new_AGEMA_signal_17944), .Z0_t (RoundReg_Inst_ff_SDE_10_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18446), .Z1_t (new_AGEMA_signal_18447), .Z1_f (new_AGEMA_signal_18448) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_10_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_10_MUX_inst_Y), .A0_f (new_AGEMA_signal_18446), .A1_t (new_AGEMA_signal_18447), .A1_f (new_AGEMA_signal_18448), .B0_t (RoundOutput[10]), .B0_f (new_AGEMA_signal_17279), .B1_t (new_AGEMA_signal_17280), .B1_f (new_AGEMA_signal_17281), .Z0_t (RoundInput[10]), .Z0_f (new_AGEMA_signal_5159), .Z1_t (new_AGEMA_signal_5160), .Z1_f (new_AGEMA_signal_5161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_11_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[11]), .A0_f (new_AGEMA_signal_17780), .A1_t (new_AGEMA_signal_17781), .A1_f (new_AGEMA_signal_17782), .B0_t (plaintext_s0_t[11]), .B0_f (plaintext_s0_f[11]), .B1_t (plaintext_s1_t[11]), .B1_f (plaintext_s1_f[11]), .Z0_t (RoundReg_Inst_ff_SDE_11_MUX_inst_X), .Z0_f (new_AGEMA_signal_18452), .Z1_t (new_AGEMA_signal_18453), .Z1_f (new_AGEMA_signal_18454) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_11_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_11_MUX_inst_X), .B0_f (new_AGEMA_signal_18452), .B1_t (new_AGEMA_signal_18453), .B1_f (new_AGEMA_signal_18454), .Z0_t (RoundReg_Inst_ff_SDE_11_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18944), .Z1_t (new_AGEMA_signal_18945), .Z1_f (new_AGEMA_signal_18946) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_11_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_11_MUX_inst_Y), .A0_f (new_AGEMA_signal_18944), .A1_t (new_AGEMA_signal_18945), .A1_f (new_AGEMA_signal_18946), .B0_t (RoundOutput[11]), .B0_f (new_AGEMA_signal_17780), .B1_t (new_AGEMA_signal_17781), .B1_f (new_AGEMA_signal_17782), .Z0_t (RoundInput[11]), .Z0_f (new_AGEMA_signal_5258), .Z1_t (new_AGEMA_signal_5259), .Z1_f (new_AGEMA_signal_5260) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_12_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[12]), .A0_f (new_AGEMA_signal_17792), .A1_t (new_AGEMA_signal_17793), .A1_f (new_AGEMA_signal_17794), .B0_t (plaintext_s0_t[12]), .B0_f (plaintext_s0_f[12]), .B1_t (plaintext_s1_t[12]), .B1_f (plaintext_s1_f[12]), .Z0_t (RoundReg_Inst_ff_SDE_12_MUX_inst_X), .Z0_f (new_AGEMA_signal_18458), .Z1_t (new_AGEMA_signal_18459), .Z1_f (new_AGEMA_signal_18460) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_12_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_12_MUX_inst_X), .B0_f (new_AGEMA_signal_18458), .B1_t (new_AGEMA_signal_18459), .B1_f (new_AGEMA_signal_18460), .Z0_t (RoundReg_Inst_ff_SDE_12_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18947), .Z1_t (new_AGEMA_signal_18948), .Z1_f (new_AGEMA_signal_18949) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_12_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_12_MUX_inst_Y), .A0_f (new_AGEMA_signal_18947), .A1_t (new_AGEMA_signal_18948), .A1_f (new_AGEMA_signal_18949), .B0_t (RoundOutput[12]), .B0_f (new_AGEMA_signal_17792), .B1_t (new_AGEMA_signal_17793), .B1_f (new_AGEMA_signal_17794), .Z0_t (RoundInput[12]), .Z0_f (new_AGEMA_signal_5339), .Z1_t (new_AGEMA_signal_5340), .Z1_f (new_AGEMA_signal_5341) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_13_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[13]), .A0_f (new_AGEMA_signal_17342), .A1_t (new_AGEMA_signal_17343), .A1_f (new_AGEMA_signal_17344), .B0_t (plaintext_s0_t[13]), .B0_f (plaintext_s0_f[13]), .B1_t (plaintext_s1_t[13]), .B1_f (plaintext_s1_f[13]), .Z0_t (RoundReg_Inst_ff_SDE_13_MUX_inst_X), .Z0_f (new_AGEMA_signal_17948), .Z1_t (new_AGEMA_signal_17949), .Z1_f (new_AGEMA_signal_17950) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_13_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_13_MUX_inst_X), .B0_f (new_AGEMA_signal_17948), .B1_t (new_AGEMA_signal_17949), .B1_f (new_AGEMA_signal_17950), .Z0_t (RoundReg_Inst_ff_SDE_13_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18461), .Z1_t (new_AGEMA_signal_18462), .Z1_f (new_AGEMA_signal_18463) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_13_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_13_MUX_inst_Y), .A0_f (new_AGEMA_signal_18461), .A1_t (new_AGEMA_signal_18462), .A1_f (new_AGEMA_signal_18463), .B0_t (RoundOutput[13]), .B0_f (new_AGEMA_signal_17342), .B1_t (new_AGEMA_signal_17343), .B1_f (new_AGEMA_signal_17344), .Z0_t (RoundInput[13]), .Z0_f (new_AGEMA_signal_5348), .Z1_t (new_AGEMA_signal_5349), .Z1_f (new_AGEMA_signal_5350) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_14_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[14]), .A0_f (new_AGEMA_signal_17345), .A1_t (new_AGEMA_signal_17346), .A1_f (new_AGEMA_signal_17347), .B0_t (plaintext_s0_t[14]), .B0_f (plaintext_s0_f[14]), .B1_t (plaintext_s1_t[14]), .B1_f (plaintext_s1_f[14]), .Z0_t (RoundReg_Inst_ff_SDE_14_MUX_inst_X), .Z0_f (new_AGEMA_signal_17954), .Z1_t (new_AGEMA_signal_17955), .Z1_f (new_AGEMA_signal_17956) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_14_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_14_MUX_inst_X), .B0_f (new_AGEMA_signal_17954), .B1_t (new_AGEMA_signal_17955), .B1_f (new_AGEMA_signal_17956), .Z0_t (RoundReg_Inst_ff_SDE_14_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18464), .Z1_t (new_AGEMA_signal_18465), .Z1_f (new_AGEMA_signal_18466) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_14_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_14_MUX_inst_Y), .A0_f (new_AGEMA_signal_18464), .A1_t (new_AGEMA_signal_18465), .A1_f (new_AGEMA_signal_18466), .B0_t (RoundOutput[14]), .B0_f (new_AGEMA_signal_17345), .B1_t (new_AGEMA_signal_17346), .B1_f (new_AGEMA_signal_17347), .Z0_t (RoundInput[14]), .Z0_f (new_AGEMA_signal_5357), .Z1_t (new_AGEMA_signal_5358), .Z1_f (new_AGEMA_signal_5359) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_15_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[15]), .A0_f (new_AGEMA_signal_17348), .A1_t (new_AGEMA_signal_17349), .A1_f (new_AGEMA_signal_17350), .B0_t (plaintext_s0_t[15]), .B0_f (plaintext_s0_f[15]), .B1_t (plaintext_s1_t[15]), .B1_f (plaintext_s1_f[15]), .Z0_t (RoundReg_Inst_ff_SDE_15_MUX_inst_X), .Z0_f (new_AGEMA_signal_17960), .Z1_t (new_AGEMA_signal_17961), .Z1_f (new_AGEMA_signal_17962) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_15_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_15_MUX_inst_X), .B0_f (new_AGEMA_signal_17960), .B1_t (new_AGEMA_signal_17961), .B1_f (new_AGEMA_signal_17962), .Z0_t (RoundReg_Inst_ff_SDE_15_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18467), .Z1_t (new_AGEMA_signal_18468), .Z1_f (new_AGEMA_signal_18469) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_15_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_15_MUX_inst_Y), .A0_f (new_AGEMA_signal_18467), .A1_t (new_AGEMA_signal_18468), .A1_f (new_AGEMA_signal_18469), .B0_t (RoundOutput[15]), .B0_f (new_AGEMA_signal_17348), .B1_t (new_AGEMA_signal_17349), .B1_f (new_AGEMA_signal_17350), .Z0_t (RoundInput[15]), .Z0_f (new_AGEMA_signal_5366), .Z1_t (new_AGEMA_signal_5367), .Z1_f (new_AGEMA_signal_5368) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_16_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[16]), .A0_f (new_AGEMA_signal_17351), .A1_t (new_AGEMA_signal_17352), .A1_f (new_AGEMA_signal_17353), .B0_t (plaintext_s0_t[16]), .B0_f (plaintext_s0_f[16]), .B1_t (plaintext_s1_t[16]), .B1_f (plaintext_s1_f[16]), .Z0_t (RoundReg_Inst_ff_SDE_16_MUX_inst_X), .Z0_f (new_AGEMA_signal_17966), .Z1_t (new_AGEMA_signal_17967), .Z1_f (new_AGEMA_signal_17968) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_16_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_16_MUX_inst_X), .B0_f (new_AGEMA_signal_17966), .B1_t (new_AGEMA_signal_17967), .B1_f (new_AGEMA_signal_17968), .Z0_t (RoundReg_Inst_ff_SDE_16_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18470), .Z1_t (new_AGEMA_signal_18471), .Z1_f (new_AGEMA_signal_18472) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_16_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_16_MUX_inst_Y), .A0_f (new_AGEMA_signal_18470), .A1_t (new_AGEMA_signal_18471), .A1_f (new_AGEMA_signal_18472), .B0_t (RoundOutput[16]), .B0_f (new_AGEMA_signal_17351), .B1_t (new_AGEMA_signal_17352), .B1_f (new_AGEMA_signal_17353), .Z0_t (RoundInput[16]), .Z0_f (new_AGEMA_signal_5375), .Z1_t (new_AGEMA_signal_5376), .Z1_f (new_AGEMA_signal_5377) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_17_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[17]), .A0_f (new_AGEMA_signal_17795), .A1_t (new_AGEMA_signal_17796), .A1_f (new_AGEMA_signal_17797), .B0_t (plaintext_s0_t[17]), .B0_f (plaintext_s0_f[17]), .B1_t (plaintext_s1_t[17]), .B1_f (plaintext_s1_f[17]), .Z0_t (RoundReg_Inst_ff_SDE_17_MUX_inst_X), .Z0_f (new_AGEMA_signal_18476), .Z1_t (new_AGEMA_signal_18477), .Z1_f (new_AGEMA_signal_18478) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_17_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_17_MUX_inst_X), .B0_f (new_AGEMA_signal_18476), .B1_t (new_AGEMA_signal_18477), .B1_f (new_AGEMA_signal_18478), .Z0_t (RoundReg_Inst_ff_SDE_17_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18950), .Z1_t (new_AGEMA_signal_18951), .Z1_f (new_AGEMA_signal_18952) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_17_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_17_MUX_inst_Y), .A0_f (new_AGEMA_signal_18950), .A1_t (new_AGEMA_signal_18951), .A1_f (new_AGEMA_signal_18952), .B0_t (RoundOutput[17]), .B0_f (new_AGEMA_signal_17795), .B1_t (new_AGEMA_signal_17796), .B1_f (new_AGEMA_signal_17797), .Z0_t (RoundInput[17]), .Z0_f (new_AGEMA_signal_5384), .Z1_t (new_AGEMA_signal_5385), .Z1_f (new_AGEMA_signal_5386) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_18_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[18]), .A0_f (new_AGEMA_signal_17357), .A1_t (new_AGEMA_signal_17358), .A1_f (new_AGEMA_signal_17359), .B0_t (plaintext_s0_t[18]), .B0_f (plaintext_s0_f[18]), .B1_t (plaintext_s1_t[18]), .B1_f (plaintext_s1_f[18]), .Z0_t (RoundReg_Inst_ff_SDE_18_MUX_inst_X), .Z0_f (new_AGEMA_signal_17972), .Z1_t (new_AGEMA_signal_17973), .Z1_f (new_AGEMA_signal_17974) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_18_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_18_MUX_inst_X), .B0_f (new_AGEMA_signal_17972), .B1_t (new_AGEMA_signal_17973), .B1_f (new_AGEMA_signal_17974), .Z0_t (RoundReg_Inst_ff_SDE_18_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18479), .Z1_t (new_AGEMA_signal_18480), .Z1_f (new_AGEMA_signal_18481) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_18_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_18_MUX_inst_Y), .A0_f (new_AGEMA_signal_18479), .A1_t (new_AGEMA_signal_18480), .A1_f (new_AGEMA_signal_18481), .B0_t (RoundOutput[18]), .B0_f (new_AGEMA_signal_17357), .B1_t (new_AGEMA_signal_17358), .B1_f (new_AGEMA_signal_17359), .Z0_t (RoundInput[18]), .Z0_f (new_AGEMA_signal_5393), .Z1_t (new_AGEMA_signal_5394), .Z1_f (new_AGEMA_signal_5395) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_19_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[19]), .A0_f (new_AGEMA_signal_17798), .A1_t (new_AGEMA_signal_17799), .A1_f (new_AGEMA_signal_17800), .B0_t (plaintext_s0_t[19]), .B0_f (plaintext_s0_f[19]), .B1_t (plaintext_s1_t[19]), .B1_f (plaintext_s1_f[19]), .Z0_t (RoundReg_Inst_ff_SDE_19_MUX_inst_X), .Z0_f (new_AGEMA_signal_18485), .Z1_t (new_AGEMA_signal_18486), .Z1_f (new_AGEMA_signal_18487) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_19_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_19_MUX_inst_X), .B0_f (new_AGEMA_signal_18485), .B1_t (new_AGEMA_signal_18486), .B1_f (new_AGEMA_signal_18487), .Z0_t (RoundReg_Inst_ff_SDE_19_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18953), .Z1_t (new_AGEMA_signal_18954), .Z1_f (new_AGEMA_signal_18955) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_19_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_19_MUX_inst_Y), .A0_f (new_AGEMA_signal_18953), .A1_t (new_AGEMA_signal_18954), .A1_f (new_AGEMA_signal_18955), .B0_t (RoundOutput[19]), .B0_f (new_AGEMA_signal_17798), .B1_t (new_AGEMA_signal_17799), .B1_f (new_AGEMA_signal_17800), .Z0_t (RoundInput[19]), .Z0_f (new_AGEMA_signal_5402), .Z1_t (new_AGEMA_signal_5403), .Z1_f (new_AGEMA_signal_5404) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_20_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[20]), .A0_f (new_AGEMA_signal_17804), .A1_t (new_AGEMA_signal_17805), .A1_f (new_AGEMA_signal_17806), .B0_t (plaintext_s0_t[20]), .B0_f (plaintext_s0_f[20]), .B1_t (plaintext_s1_t[20]), .B1_f (plaintext_s1_f[20]), .Z0_t (RoundReg_Inst_ff_SDE_20_MUX_inst_X), .Z0_f (new_AGEMA_signal_18491), .Z1_t (new_AGEMA_signal_18492), .Z1_f (new_AGEMA_signal_18493) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_20_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_20_MUX_inst_X), .B0_f (new_AGEMA_signal_18491), .B1_t (new_AGEMA_signal_18492), .B1_f (new_AGEMA_signal_18493), .Z0_t (RoundReg_Inst_ff_SDE_20_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18956), .Z1_t (new_AGEMA_signal_18957), .Z1_f (new_AGEMA_signal_18958) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_20_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_20_MUX_inst_Y), .A0_f (new_AGEMA_signal_18956), .A1_t (new_AGEMA_signal_18957), .A1_f (new_AGEMA_signal_18958), .B0_t (RoundOutput[20]), .B0_f (new_AGEMA_signal_17804), .B1_t (new_AGEMA_signal_17805), .B1_f (new_AGEMA_signal_17806), .Z0_t (RoundInput[20]), .Z0_f (new_AGEMA_signal_5420), .Z1_t (new_AGEMA_signal_5421), .Z1_f (new_AGEMA_signal_5422) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_21_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[21]), .A0_f (new_AGEMA_signal_17369), .A1_t (new_AGEMA_signal_17370), .A1_f (new_AGEMA_signal_17371), .B0_t (plaintext_s0_t[21]), .B0_f (plaintext_s0_f[21]), .B1_t (plaintext_s1_t[21]), .B1_f (plaintext_s1_f[21]), .Z0_t (RoundReg_Inst_ff_SDE_21_MUX_inst_X), .Z0_f (new_AGEMA_signal_17978), .Z1_t (new_AGEMA_signal_17979), .Z1_f (new_AGEMA_signal_17980) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_21_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_21_MUX_inst_X), .B0_f (new_AGEMA_signal_17978), .B1_t (new_AGEMA_signal_17979), .B1_f (new_AGEMA_signal_17980), .Z0_t (RoundReg_Inst_ff_SDE_21_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18494), .Z1_t (new_AGEMA_signal_18495), .Z1_f (new_AGEMA_signal_18496) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_21_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_21_MUX_inst_Y), .A0_f (new_AGEMA_signal_18494), .A1_t (new_AGEMA_signal_18495), .A1_f (new_AGEMA_signal_18496), .B0_t (RoundOutput[21]), .B0_f (new_AGEMA_signal_17369), .B1_t (new_AGEMA_signal_17370), .B1_f (new_AGEMA_signal_17371), .Z0_t (RoundInput[21]), .Z0_f (new_AGEMA_signal_5429), .Z1_t (new_AGEMA_signal_5430), .Z1_f (new_AGEMA_signal_5431) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_22_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[22]), .A0_f (new_AGEMA_signal_17372), .A1_t (new_AGEMA_signal_17373), .A1_f (new_AGEMA_signal_17374), .B0_t (plaintext_s0_t[22]), .B0_f (plaintext_s0_f[22]), .B1_t (plaintext_s1_t[22]), .B1_f (plaintext_s1_f[22]), .Z0_t (RoundReg_Inst_ff_SDE_22_MUX_inst_X), .Z0_f (new_AGEMA_signal_17984), .Z1_t (new_AGEMA_signal_17985), .Z1_f (new_AGEMA_signal_17986) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_22_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_22_MUX_inst_X), .B0_f (new_AGEMA_signal_17984), .B1_t (new_AGEMA_signal_17985), .B1_f (new_AGEMA_signal_17986), .Z0_t (RoundReg_Inst_ff_SDE_22_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18497), .Z1_t (new_AGEMA_signal_18498), .Z1_f (new_AGEMA_signal_18499) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_22_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_22_MUX_inst_Y), .A0_f (new_AGEMA_signal_18497), .A1_t (new_AGEMA_signal_18498), .A1_f (new_AGEMA_signal_18499), .B0_t (RoundOutput[22]), .B0_f (new_AGEMA_signal_17372), .B1_t (new_AGEMA_signal_17373), .B1_f (new_AGEMA_signal_17374), .Z0_t (RoundInput[22]), .Z0_f (new_AGEMA_signal_5438), .Z1_t (new_AGEMA_signal_5439), .Z1_f (new_AGEMA_signal_5440) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_23_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[23]), .A0_f (new_AGEMA_signal_17375), .A1_t (new_AGEMA_signal_17376), .A1_f (new_AGEMA_signal_17377), .B0_t (plaintext_s0_t[23]), .B0_f (plaintext_s0_f[23]), .B1_t (plaintext_s1_t[23]), .B1_f (plaintext_s1_f[23]), .Z0_t (RoundReg_Inst_ff_SDE_23_MUX_inst_X), .Z0_f (new_AGEMA_signal_17990), .Z1_t (new_AGEMA_signal_17991), .Z1_f (new_AGEMA_signal_17992) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_23_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_23_MUX_inst_X), .B0_f (new_AGEMA_signal_17990), .B1_t (new_AGEMA_signal_17991), .B1_f (new_AGEMA_signal_17992), .Z0_t (RoundReg_Inst_ff_SDE_23_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18500), .Z1_t (new_AGEMA_signal_18501), .Z1_f (new_AGEMA_signal_18502) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_23_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_23_MUX_inst_Y), .A0_f (new_AGEMA_signal_18500), .A1_t (new_AGEMA_signal_18501), .A1_f (new_AGEMA_signal_18502), .B0_t (RoundOutput[23]), .B0_f (new_AGEMA_signal_17375), .B1_t (new_AGEMA_signal_17376), .B1_f (new_AGEMA_signal_17377), .Z0_t (RoundInput[23]), .Z0_f (new_AGEMA_signal_5447), .Z1_t (new_AGEMA_signal_5448), .Z1_f (new_AGEMA_signal_5449) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_24_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[24]), .A0_f (new_AGEMA_signal_17378), .A1_t (new_AGEMA_signal_17379), .A1_f (new_AGEMA_signal_17380), .B0_t (plaintext_s0_t[24]), .B0_f (plaintext_s0_f[24]), .B1_t (plaintext_s1_t[24]), .B1_f (plaintext_s1_f[24]), .Z0_t (RoundReg_Inst_ff_SDE_24_MUX_inst_X), .Z0_f (new_AGEMA_signal_17996), .Z1_t (new_AGEMA_signal_17997), .Z1_f (new_AGEMA_signal_17998) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_24_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_24_MUX_inst_X), .B0_f (new_AGEMA_signal_17996), .B1_t (new_AGEMA_signal_17997), .B1_f (new_AGEMA_signal_17998), .Z0_t (RoundReg_Inst_ff_SDE_24_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18503), .Z1_t (new_AGEMA_signal_18504), .Z1_f (new_AGEMA_signal_18505) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_24_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_24_MUX_inst_Y), .A0_f (new_AGEMA_signal_18503), .A1_t (new_AGEMA_signal_18504), .A1_f (new_AGEMA_signal_18505), .B0_t (RoundOutput[24]), .B0_f (new_AGEMA_signal_17378), .B1_t (new_AGEMA_signal_17379), .B1_f (new_AGEMA_signal_17380), .Z0_t (RoundInput[24]), .Z0_f (new_AGEMA_signal_5456), .Z1_t (new_AGEMA_signal_5457), .Z1_f (new_AGEMA_signal_5458) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_25_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[25]), .A0_f (new_AGEMA_signal_17807), .A1_t (new_AGEMA_signal_17808), .A1_f (new_AGEMA_signal_17809), .B0_t (plaintext_s0_t[25]), .B0_f (plaintext_s0_f[25]), .B1_t (plaintext_s1_t[25]), .B1_f (plaintext_s1_f[25]), .Z0_t (RoundReg_Inst_ff_SDE_25_MUX_inst_X), .Z0_f (new_AGEMA_signal_18509), .Z1_t (new_AGEMA_signal_18510), .Z1_f (new_AGEMA_signal_18511) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_25_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_25_MUX_inst_X), .B0_f (new_AGEMA_signal_18509), .B1_t (new_AGEMA_signal_18510), .B1_f (new_AGEMA_signal_18511), .Z0_t (RoundReg_Inst_ff_SDE_25_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18959), .Z1_t (new_AGEMA_signal_18960), .Z1_f (new_AGEMA_signal_18961) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_25_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_25_MUX_inst_Y), .A0_f (new_AGEMA_signal_18959), .A1_t (new_AGEMA_signal_18960), .A1_f (new_AGEMA_signal_18961), .B0_t (RoundOutput[25]), .B0_f (new_AGEMA_signal_17807), .B1_t (new_AGEMA_signal_17808), .B1_f (new_AGEMA_signal_17809), .Z0_t (RoundInput[25]), .Z0_f (new_AGEMA_signal_5465), .Z1_t (new_AGEMA_signal_5466), .Z1_f (new_AGEMA_signal_5467) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_26_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[26]), .A0_f (new_AGEMA_signal_17384), .A1_t (new_AGEMA_signal_17385), .A1_f (new_AGEMA_signal_17386), .B0_t (plaintext_s0_t[26]), .B0_f (plaintext_s0_f[26]), .B1_t (plaintext_s1_t[26]), .B1_f (plaintext_s1_f[26]), .Z0_t (RoundReg_Inst_ff_SDE_26_MUX_inst_X), .Z0_f (new_AGEMA_signal_18002), .Z1_t (new_AGEMA_signal_18003), .Z1_f (new_AGEMA_signal_18004) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_26_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_26_MUX_inst_X), .B0_f (new_AGEMA_signal_18002), .B1_t (new_AGEMA_signal_18003), .B1_f (new_AGEMA_signal_18004), .Z0_t (RoundReg_Inst_ff_SDE_26_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18512), .Z1_t (new_AGEMA_signal_18513), .Z1_f (new_AGEMA_signal_18514) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_26_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_26_MUX_inst_Y), .A0_f (new_AGEMA_signal_18512), .A1_t (new_AGEMA_signal_18513), .A1_f (new_AGEMA_signal_18514), .B0_t (RoundOutput[26]), .B0_f (new_AGEMA_signal_17384), .B1_t (new_AGEMA_signal_17385), .B1_f (new_AGEMA_signal_17386), .Z0_t (RoundInput[26]), .Z0_f (new_AGEMA_signal_5474), .Z1_t (new_AGEMA_signal_5475), .Z1_f (new_AGEMA_signal_5476) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_27_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[27]), .A0_f (new_AGEMA_signal_17810), .A1_t (new_AGEMA_signal_17811), .A1_f (new_AGEMA_signal_17812), .B0_t (plaintext_s0_t[27]), .B0_f (plaintext_s0_f[27]), .B1_t (plaintext_s1_t[27]), .B1_f (plaintext_s1_f[27]), .Z0_t (RoundReg_Inst_ff_SDE_27_MUX_inst_X), .Z0_f (new_AGEMA_signal_18518), .Z1_t (new_AGEMA_signal_18519), .Z1_f (new_AGEMA_signal_18520) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_27_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_27_MUX_inst_X), .B0_f (new_AGEMA_signal_18518), .B1_t (new_AGEMA_signal_18519), .B1_f (new_AGEMA_signal_18520), .Z0_t (RoundReg_Inst_ff_SDE_27_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18962), .Z1_t (new_AGEMA_signal_18963), .Z1_f (new_AGEMA_signal_18964) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_27_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_27_MUX_inst_Y), .A0_f (new_AGEMA_signal_18962), .A1_t (new_AGEMA_signal_18963), .A1_f (new_AGEMA_signal_18964), .B0_t (RoundOutput[27]), .B0_f (new_AGEMA_signal_17810), .B1_t (new_AGEMA_signal_17811), .B1_f (new_AGEMA_signal_17812), .Z0_t (RoundInput[27]), .Z0_f (new_AGEMA_signal_5483), .Z1_t (new_AGEMA_signal_5484), .Z1_f (new_AGEMA_signal_5485) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_28_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[28]), .A0_f (new_AGEMA_signal_17813), .A1_t (new_AGEMA_signal_17814), .A1_f (new_AGEMA_signal_17815), .B0_t (plaintext_s0_t[28]), .B0_f (plaintext_s0_f[28]), .B1_t (plaintext_s1_t[28]), .B1_f (plaintext_s1_f[28]), .Z0_t (RoundReg_Inst_ff_SDE_28_MUX_inst_X), .Z0_f (new_AGEMA_signal_18524), .Z1_t (new_AGEMA_signal_18525), .Z1_f (new_AGEMA_signal_18526) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_28_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_28_MUX_inst_X), .B0_f (new_AGEMA_signal_18524), .B1_t (new_AGEMA_signal_18525), .B1_f (new_AGEMA_signal_18526), .Z0_t (RoundReg_Inst_ff_SDE_28_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18965), .Z1_t (new_AGEMA_signal_18966), .Z1_f (new_AGEMA_signal_18967) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_28_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_28_MUX_inst_Y), .A0_f (new_AGEMA_signal_18965), .A1_t (new_AGEMA_signal_18966), .A1_f (new_AGEMA_signal_18967), .B0_t (RoundOutput[28]), .B0_f (new_AGEMA_signal_17813), .B1_t (new_AGEMA_signal_17814), .B1_f (new_AGEMA_signal_17815), .Z0_t (RoundInput[28]), .Z0_f (new_AGEMA_signal_5492), .Z1_t (new_AGEMA_signal_5493), .Z1_f (new_AGEMA_signal_5494) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_29_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[29]), .A0_f (new_AGEMA_signal_17393), .A1_t (new_AGEMA_signal_17394), .A1_f (new_AGEMA_signal_17395), .B0_t (plaintext_s0_t[29]), .B0_f (plaintext_s0_f[29]), .B1_t (plaintext_s1_t[29]), .B1_f (plaintext_s1_f[29]), .Z0_t (RoundReg_Inst_ff_SDE_29_MUX_inst_X), .Z0_f (new_AGEMA_signal_18008), .Z1_t (new_AGEMA_signal_18009), .Z1_f (new_AGEMA_signal_18010) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_29_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_29_MUX_inst_X), .B0_f (new_AGEMA_signal_18008), .B1_t (new_AGEMA_signal_18009), .B1_f (new_AGEMA_signal_18010), .Z0_t (RoundReg_Inst_ff_SDE_29_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18527), .Z1_t (new_AGEMA_signal_18528), .Z1_f (new_AGEMA_signal_18529) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_29_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_29_MUX_inst_Y), .A0_f (new_AGEMA_signal_18527), .A1_t (new_AGEMA_signal_18528), .A1_f (new_AGEMA_signal_18529), .B0_t (RoundOutput[29]), .B0_f (new_AGEMA_signal_17393), .B1_t (new_AGEMA_signal_17394), .B1_f (new_AGEMA_signal_17395), .Z0_t (RoundInput[29]), .Z0_f (new_AGEMA_signal_5501), .Z1_t (new_AGEMA_signal_5502), .Z1_f (new_AGEMA_signal_5503) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_30_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[30]), .A0_f (new_AGEMA_signal_17399), .A1_t (new_AGEMA_signal_17400), .A1_f (new_AGEMA_signal_17401), .B0_t (plaintext_s0_t[30]), .B0_f (plaintext_s0_f[30]), .B1_t (plaintext_s1_t[30]), .B1_f (plaintext_s1_f[30]), .Z0_t (RoundReg_Inst_ff_SDE_30_MUX_inst_X), .Z0_f (new_AGEMA_signal_18014), .Z1_t (new_AGEMA_signal_18015), .Z1_f (new_AGEMA_signal_18016) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_30_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_30_MUX_inst_X), .B0_f (new_AGEMA_signal_18014), .B1_t (new_AGEMA_signal_18015), .B1_f (new_AGEMA_signal_18016), .Z0_t (RoundReg_Inst_ff_SDE_30_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18530), .Z1_t (new_AGEMA_signal_18531), .Z1_f (new_AGEMA_signal_18532) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_30_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_30_MUX_inst_Y), .A0_f (new_AGEMA_signal_18530), .A1_t (new_AGEMA_signal_18531), .A1_f (new_AGEMA_signal_18532), .B0_t (RoundOutput[30]), .B0_f (new_AGEMA_signal_17399), .B1_t (new_AGEMA_signal_17400), .B1_f (new_AGEMA_signal_17401), .Z0_t (RoundInput[30]), .Z0_f (new_AGEMA_signal_5519), .Z1_t (new_AGEMA_signal_5520), .Z1_f (new_AGEMA_signal_5521) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_31_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[31]), .A0_f (new_AGEMA_signal_17402), .A1_t (new_AGEMA_signal_17403), .A1_f (new_AGEMA_signal_17404), .B0_t (plaintext_s0_t[31]), .B0_f (plaintext_s0_f[31]), .B1_t (plaintext_s1_t[31]), .B1_f (plaintext_s1_f[31]), .Z0_t (RoundReg_Inst_ff_SDE_31_MUX_inst_X), .Z0_f (new_AGEMA_signal_18020), .Z1_t (new_AGEMA_signal_18021), .Z1_f (new_AGEMA_signal_18022) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_31_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_31_MUX_inst_X), .B0_f (new_AGEMA_signal_18020), .B1_t (new_AGEMA_signal_18021), .B1_f (new_AGEMA_signal_18022), .Z0_t (RoundReg_Inst_ff_SDE_31_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18533), .Z1_t (new_AGEMA_signal_18534), .Z1_f (new_AGEMA_signal_18535) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_31_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_31_MUX_inst_Y), .A0_f (new_AGEMA_signal_18533), .A1_t (new_AGEMA_signal_18534), .A1_f (new_AGEMA_signal_18535), .B0_t (RoundOutput[31]), .B0_f (new_AGEMA_signal_17402), .B1_t (new_AGEMA_signal_17403), .B1_f (new_AGEMA_signal_17404), .Z0_t (RoundInput[31]), .Z0_f (new_AGEMA_signal_5528), .Z1_t (new_AGEMA_signal_5529), .Z1_f (new_AGEMA_signal_5530) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_32_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[32]), .A0_f (new_AGEMA_signal_17405), .A1_t (new_AGEMA_signal_17406), .A1_f (new_AGEMA_signal_17407), .B0_t (plaintext_s0_t[32]), .B0_f (plaintext_s0_f[32]), .B1_t (plaintext_s1_t[32]), .B1_f (plaintext_s1_f[32]), .Z0_t (RoundReg_Inst_ff_SDE_32_MUX_inst_X), .Z0_f (new_AGEMA_signal_18026), .Z1_t (new_AGEMA_signal_18027), .Z1_f (new_AGEMA_signal_18028) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_32_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_32_MUX_inst_X), .B0_f (new_AGEMA_signal_18026), .B1_t (new_AGEMA_signal_18027), .B1_f (new_AGEMA_signal_18028), .Z0_t (RoundReg_Inst_ff_SDE_32_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18536), .Z1_t (new_AGEMA_signal_18537), .Z1_f (new_AGEMA_signal_18538) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_32_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_32_MUX_inst_Y), .A0_f (new_AGEMA_signal_18536), .A1_t (new_AGEMA_signal_18537), .A1_f (new_AGEMA_signal_18538), .B0_t (RoundOutput[32]), .B0_f (new_AGEMA_signal_17405), .B1_t (new_AGEMA_signal_17406), .B1_f (new_AGEMA_signal_17407), .Z0_t (RoundInput[32]), .Z0_f (new_AGEMA_signal_5537), .Z1_t (new_AGEMA_signal_5538), .Z1_f (new_AGEMA_signal_5539) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_33_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[33]), .A0_f (new_AGEMA_signal_17816), .A1_t (new_AGEMA_signal_17817), .A1_f (new_AGEMA_signal_17818), .B0_t (plaintext_s0_t[33]), .B0_f (plaintext_s0_f[33]), .B1_t (plaintext_s1_t[33]), .B1_f (plaintext_s1_f[33]), .Z0_t (RoundReg_Inst_ff_SDE_33_MUX_inst_X), .Z0_f (new_AGEMA_signal_18542), .Z1_t (new_AGEMA_signal_18543), .Z1_f (new_AGEMA_signal_18544) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_33_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_33_MUX_inst_X), .B0_f (new_AGEMA_signal_18542), .B1_t (new_AGEMA_signal_18543), .B1_f (new_AGEMA_signal_18544), .Z0_t (RoundReg_Inst_ff_SDE_33_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18968), .Z1_t (new_AGEMA_signal_18969), .Z1_f (new_AGEMA_signal_18970) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_33_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_33_MUX_inst_Y), .A0_f (new_AGEMA_signal_18968), .A1_t (new_AGEMA_signal_18969), .A1_f (new_AGEMA_signal_18970), .B0_t (RoundOutput[33]), .B0_f (new_AGEMA_signal_17816), .B1_t (new_AGEMA_signal_17817), .B1_f (new_AGEMA_signal_17818), .Z0_t (RoundInput[33]), .Z0_f (new_AGEMA_signal_5546), .Z1_t (new_AGEMA_signal_5547), .Z1_f (new_AGEMA_signal_5548) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_34_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[34]), .A0_f (new_AGEMA_signal_17411), .A1_t (new_AGEMA_signal_17412), .A1_f (new_AGEMA_signal_17413), .B0_t (plaintext_s0_t[34]), .B0_f (plaintext_s0_f[34]), .B1_t (plaintext_s1_t[34]), .B1_f (plaintext_s1_f[34]), .Z0_t (RoundReg_Inst_ff_SDE_34_MUX_inst_X), .Z0_f (new_AGEMA_signal_18032), .Z1_t (new_AGEMA_signal_18033), .Z1_f (new_AGEMA_signal_18034) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_34_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_34_MUX_inst_X), .B0_f (new_AGEMA_signal_18032), .B1_t (new_AGEMA_signal_18033), .B1_f (new_AGEMA_signal_18034), .Z0_t (RoundReg_Inst_ff_SDE_34_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18545), .Z1_t (new_AGEMA_signal_18546), .Z1_f (new_AGEMA_signal_18547) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_34_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_34_MUX_inst_Y), .A0_f (new_AGEMA_signal_18545), .A1_t (new_AGEMA_signal_18546), .A1_f (new_AGEMA_signal_18547), .B0_t (RoundOutput[34]), .B0_f (new_AGEMA_signal_17411), .B1_t (new_AGEMA_signal_17412), .B1_f (new_AGEMA_signal_17413), .Z0_t (RoundInput[34]), .Z0_f (new_AGEMA_signal_5555), .Z1_t (new_AGEMA_signal_5556), .Z1_f (new_AGEMA_signal_5557) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_35_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[35]), .A0_f (new_AGEMA_signal_17819), .A1_t (new_AGEMA_signal_17820), .A1_f (new_AGEMA_signal_17821), .B0_t (plaintext_s0_t[35]), .B0_f (plaintext_s0_f[35]), .B1_t (plaintext_s1_t[35]), .B1_f (plaintext_s1_f[35]), .Z0_t (RoundReg_Inst_ff_SDE_35_MUX_inst_X), .Z0_f (new_AGEMA_signal_18551), .Z1_t (new_AGEMA_signal_18552), .Z1_f (new_AGEMA_signal_18553) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_35_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_35_MUX_inst_X), .B0_f (new_AGEMA_signal_18551), .B1_t (new_AGEMA_signal_18552), .B1_f (new_AGEMA_signal_18553), .Z0_t (RoundReg_Inst_ff_SDE_35_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18971), .Z1_t (new_AGEMA_signal_18972), .Z1_f (new_AGEMA_signal_18973) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_35_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_35_MUX_inst_Y), .A0_f (new_AGEMA_signal_18971), .A1_t (new_AGEMA_signal_18972), .A1_f (new_AGEMA_signal_18973), .B0_t (RoundOutput[35]), .B0_f (new_AGEMA_signal_17819), .B1_t (new_AGEMA_signal_17820), .B1_f (new_AGEMA_signal_17821), .Z0_t (RoundInput[35]), .Z0_f (new_AGEMA_signal_5564), .Z1_t (new_AGEMA_signal_5565), .Z1_f (new_AGEMA_signal_5566) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_36_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[36]), .A0_f (new_AGEMA_signal_17822), .A1_t (new_AGEMA_signal_17823), .A1_f (new_AGEMA_signal_17824), .B0_t (plaintext_s0_t[36]), .B0_f (plaintext_s0_f[36]), .B1_t (plaintext_s1_t[36]), .B1_f (plaintext_s1_f[36]), .Z0_t (RoundReg_Inst_ff_SDE_36_MUX_inst_X), .Z0_f (new_AGEMA_signal_18557), .Z1_t (new_AGEMA_signal_18558), .Z1_f (new_AGEMA_signal_18559) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_36_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_36_MUX_inst_X), .B0_f (new_AGEMA_signal_18557), .B1_t (new_AGEMA_signal_18558), .B1_f (new_AGEMA_signal_18559), .Z0_t (RoundReg_Inst_ff_SDE_36_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18974), .Z1_t (new_AGEMA_signal_18975), .Z1_f (new_AGEMA_signal_18976) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_36_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_36_MUX_inst_Y), .A0_f (new_AGEMA_signal_18974), .A1_t (new_AGEMA_signal_18975), .A1_f (new_AGEMA_signal_18976), .B0_t (RoundOutput[36]), .B0_f (new_AGEMA_signal_17822), .B1_t (new_AGEMA_signal_17823), .B1_f (new_AGEMA_signal_17824), .Z0_t (RoundInput[36]), .Z0_f (new_AGEMA_signal_5573), .Z1_t (new_AGEMA_signal_5574), .Z1_f (new_AGEMA_signal_5575) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_37_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[37]), .A0_f (new_AGEMA_signal_17420), .A1_t (new_AGEMA_signal_17421), .A1_f (new_AGEMA_signal_17422), .B0_t (plaintext_s0_t[37]), .B0_f (plaintext_s0_f[37]), .B1_t (plaintext_s1_t[37]), .B1_f (plaintext_s1_f[37]), .Z0_t (RoundReg_Inst_ff_SDE_37_MUX_inst_X), .Z0_f (new_AGEMA_signal_18038), .Z1_t (new_AGEMA_signal_18039), .Z1_f (new_AGEMA_signal_18040) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_37_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_37_MUX_inst_X), .B0_f (new_AGEMA_signal_18038), .B1_t (new_AGEMA_signal_18039), .B1_f (new_AGEMA_signal_18040), .Z0_t (RoundReg_Inst_ff_SDE_37_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18560), .Z1_t (new_AGEMA_signal_18561), .Z1_f (new_AGEMA_signal_18562) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_37_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_37_MUX_inst_Y), .A0_f (new_AGEMA_signal_18560), .A1_t (new_AGEMA_signal_18561), .A1_f (new_AGEMA_signal_18562), .B0_t (RoundOutput[37]), .B0_f (new_AGEMA_signal_17420), .B1_t (new_AGEMA_signal_17421), .B1_f (new_AGEMA_signal_17422), .Z0_t (RoundInput[37]), .Z0_f (new_AGEMA_signal_5582), .Z1_t (new_AGEMA_signal_5583), .Z1_f (new_AGEMA_signal_5584) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_38_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[38]), .A0_f (new_AGEMA_signal_17423), .A1_t (new_AGEMA_signal_17424), .A1_f (new_AGEMA_signal_17425), .B0_t (plaintext_s0_t[38]), .B0_f (plaintext_s0_f[38]), .B1_t (plaintext_s1_t[38]), .B1_f (plaintext_s1_f[38]), .Z0_t (RoundReg_Inst_ff_SDE_38_MUX_inst_X), .Z0_f (new_AGEMA_signal_18044), .Z1_t (new_AGEMA_signal_18045), .Z1_f (new_AGEMA_signal_18046) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_38_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_38_MUX_inst_X), .B0_f (new_AGEMA_signal_18044), .B1_t (new_AGEMA_signal_18045), .B1_f (new_AGEMA_signal_18046), .Z0_t (RoundReg_Inst_ff_SDE_38_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18563), .Z1_t (new_AGEMA_signal_18564), .Z1_f (new_AGEMA_signal_18565) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_38_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_38_MUX_inst_Y), .A0_f (new_AGEMA_signal_18563), .A1_t (new_AGEMA_signal_18564), .A1_f (new_AGEMA_signal_18565), .B0_t (RoundOutput[38]), .B0_f (new_AGEMA_signal_17423), .B1_t (new_AGEMA_signal_17424), .B1_f (new_AGEMA_signal_17425), .Z0_t (RoundInput[38]), .Z0_f (new_AGEMA_signal_5591), .Z1_t (new_AGEMA_signal_5592), .Z1_f (new_AGEMA_signal_5593) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_39_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[39]), .A0_f (new_AGEMA_signal_17426), .A1_t (new_AGEMA_signal_17427), .A1_f (new_AGEMA_signal_17428), .B0_t (plaintext_s0_t[39]), .B0_f (plaintext_s0_f[39]), .B1_t (plaintext_s1_t[39]), .B1_f (plaintext_s1_f[39]), .Z0_t (RoundReg_Inst_ff_SDE_39_MUX_inst_X), .Z0_f (new_AGEMA_signal_18050), .Z1_t (new_AGEMA_signal_18051), .Z1_f (new_AGEMA_signal_18052) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_39_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_39_MUX_inst_X), .B0_f (new_AGEMA_signal_18050), .B1_t (new_AGEMA_signal_18051), .B1_f (new_AGEMA_signal_18052), .Z0_t (RoundReg_Inst_ff_SDE_39_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18566), .Z1_t (new_AGEMA_signal_18567), .Z1_f (new_AGEMA_signal_18568) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_39_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_39_MUX_inst_Y), .A0_f (new_AGEMA_signal_18566), .A1_t (new_AGEMA_signal_18567), .A1_f (new_AGEMA_signal_18568), .B0_t (RoundOutput[39]), .B0_f (new_AGEMA_signal_17426), .B1_t (new_AGEMA_signal_17427), .B1_f (new_AGEMA_signal_17428), .Z0_t (RoundInput[39]), .Z0_f (new_AGEMA_signal_5600), .Z1_t (new_AGEMA_signal_5601), .Z1_f (new_AGEMA_signal_5602) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_40_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[40]), .A0_f (new_AGEMA_signal_17432), .A1_t (new_AGEMA_signal_17433), .A1_f (new_AGEMA_signal_17434), .B0_t (plaintext_s0_t[40]), .B0_f (plaintext_s0_f[40]), .B1_t (plaintext_s1_t[40]), .B1_f (plaintext_s1_f[40]), .Z0_t (RoundReg_Inst_ff_SDE_40_MUX_inst_X), .Z0_f (new_AGEMA_signal_18056), .Z1_t (new_AGEMA_signal_18057), .Z1_f (new_AGEMA_signal_18058) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_40_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_40_MUX_inst_X), .B0_f (new_AGEMA_signal_18056), .B1_t (new_AGEMA_signal_18057), .B1_f (new_AGEMA_signal_18058), .Z0_t (RoundReg_Inst_ff_SDE_40_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18569), .Z1_t (new_AGEMA_signal_18570), .Z1_f (new_AGEMA_signal_18571) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_40_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_40_MUX_inst_Y), .A0_f (new_AGEMA_signal_18569), .A1_t (new_AGEMA_signal_18570), .A1_f (new_AGEMA_signal_18571), .B0_t (RoundOutput[40]), .B0_f (new_AGEMA_signal_17432), .B1_t (new_AGEMA_signal_17433), .B1_f (new_AGEMA_signal_17434), .Z0_t (RoundInput[40]), .Z0_f (new_AGEMA_signal_5618), .Z1_t (new_AGEMA_signal_5619), .Z1_f (new_AGEMA_signal_5620) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_41_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[41]), .A0_f (new_AGEMA_signal_17828), .A1_t (new_AGEMA_signal_17829), .A1_f (new_AGEMA_signal_17830), .B0_t (plaintext_s0_t[41]), .B0_f (plaintext_s0_f[41]), .B1_t (plaintext_s1_t[41]), .B1_f (plaintext_s1_f[41]), .Z0_t (RoundReg_Inst_ff_SDE_41_MUX_inst_X), .Z0_f (new_AGEMA_signal_18575), .Z1_t (new_AGEMA_signal_18576), .Z1_f (new_AGEMA_signal_18577) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_41_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_41_MUX_inst_X), .B0_f (new_AGEMA_signal_18575), .B1_t (new_AGEMA_signal_18576), .B1_f (new_AGEMA_signal_18577), .Z0_t (RoundReg_Inst_ff_SDE_41_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18977), .Z1_t (new_AGEMA_signal_18978), .Z1_f (new_AGEMA_signal_18979) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_41_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_41_MUX_inst_Y), .A0_f (new_AGEMA_signal_18977), .A1_t (new_AGEMA_signal_18978), .A1_f (new_AGEMA_signal_18979), .B0_t (RoundOutput[41]), .B0_f (new_AGEMA_signal_17828), .B1_t (new_AGEMA_signal_17829), .B1_f (new_AGEMA_signal_17830), .Z0_t (RoundInput[41]), .Z0_f (new_AGEMA_signal_5627), .Z1_t (new_AGEMA_signal_5628), .Z1_f (new_AGEMA_signal_5629) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_42_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[42]), .A0_f (new_AGEMA_signal_17438), .A1_t (new_AGEMA_signal_17439), .A1_f (new_AGEMA_signal_17440), .B0_t (plaintext_s0_t[42]), .B0_f (plaintext_s0_f[42]), .B1_t (plaintext_s1_t[42]), .B1_f (plaintext_s1_f[42]), .Z0_t (RoundReg_Inst_ff_SDE_42_MUX_inst_X), .Z0_f (new_AGEMA_signal_18062), .Z1_t (new_AGEMA_signal_18063), .Z1_f (new_AGEMA_signal_18064) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_42_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_42_MUX_inst_X), .B0_f (new_AGEMA_signal_18062), .B1_t (new_AGEMA_signal_18063), .B1_f (new_AGEMA_signal_18064), .Z0_t (RoundReg_Inst_ff_SDE_42_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18578), .Z1_t (new_AGEMA_signal_18579), .Z1_f (new_AGEMA_signal_18580) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_42_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_42_MUX_inst_Y), .A0_f (new_AGEMA_signal_18578), .A1_t (new_AGEMA_signal_18579), .A1_f (new_AGEMA_signal_18580), .B0_t (RoundOutput[42]), .B0_f (new_AGEMA_signal_17438), .B1_t (new_AGEMA_signal_17439), .B1_f (new_AGEMA_signal_17440), .Z0_t (RoundInput[42]), .Z0_f (new_AGEMA_signal_5636), .Z1_t (new_AGEMA_signal_5637), .Z1_f (new_AGEMA_signal_5638) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_43_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[43]), .A0_f (new_AGEMA_signal_17831), .A1_t (new_AGEMA_signal_17832), .A1_f (new_AGEMA_signal_17833), .B0_t (plaintext_s0_t[43]), .B0_f (plaintext_s0_f[43]), .B1_t (plaintext_s1_t[43]), .B1_f (plaintext_s1_f[43]), .Z0_t (RoundReg_Inst_ff_SDE_43_MUX_inst_X), .Z0_f (new_AGEMA_signal_18584), .Z1_t (new_AGEMA_signal_18585), .Z1_f (new_AGEMA_signal_18586) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_43_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_43_MUX_inst_X), .B0_f (new_AGEMA_signal_18584), .B1_t (new_AGEMA_signal_18585), .B1_f (new_AGEMA_signal_18586), .Z0_t (RoundReg_Inst_ff_SDE_43_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18980), .Z1_t (new_AGEMA_signal_18981), .Z1_f (new_AGEMA_signal_18982) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_43_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_43_MUX_inst_Y), .A0_f (new_AGEMA_signal_18980), .A1_t (new_AGEMA_signal_18981), .A1_f (new_AGEMA_signal_18982), .B0_t (RoundOutput[43]), .B0_f (new_AGEMA_signal_17831), .B1_t (new_AGEMA_signal_17832), .B1_f (new_AGEMA_signal_17833), .Z0_t (RoundInput[43]), .Z0_f (new_AGEMA_signal_5645), .Z1_t (new_AGEMA_signal_5646), .Z1_f (new_AGEMA_signal_5647) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_44_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[44]), .A0_f (new_AGEMA_signal_17834), .A1_t (new_AGEMA_signal_17835), .A1_f (new_AGEMA_signal_17836), .B0_t (plaintext_s0_t[44]), .B0_f (plaintext_s0_f[44]), .B1_t (plaintext_s1_t[44]), .B1_f (plaintext_s1_f[44]), .Z0_t (RoundReg_Inst_ff_SDE_44_MUX_inst_X), .Z0_f (new_AGEMA_signal_18590), .Z1_t (new_AGEMA_signal_18591), .Z1_f (new_AGEMA_signal_18592) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_44_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_44_MUX_inst_X), .B0_f (new_AGEMA_signal_18590), .B1_t (new_AGEMA_signal_18591), .B1_f (new_AGEMA_signal_18592), .Z0_t (RoundReg_Inst_ff_SDE_44_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18983), .Z1_t (new_AGEMA_signal_18984), .Z1_f (new_AGEMA_signal_18985) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_44_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_44_MUX_inst_Y), .A0_f (new_AGEMA_signal_18983), .A1_t (new_AGEMA_signal_18984), .A1_f (new_AGEMA_signal_18985), .B0_t (RoundOutput[44]), .B0_f (new_AGEMA_signal_17834), .B1_t (new_AGEMA_signal_17835), .B1_f (new_AGEMA_signal_17836), .Z0_t (RoundInput[44]), .Z0_f (new_AGEMA_signal_5654), .Z1_t (new_AGEMA_signal_5655), .Z1_f (new_AGEMA_signal_5656) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_45_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[45]), .A0_f (new_AGEMA_signal_17447), .A1_t (new_AGEMA_signal_17448), .A1_f (new_AGEMA_signal_17449), .B0_t (plaintext_s0_t[45]), .B0_f (plaintext_s0_f[45]), .B1_t (plaintext_s1_t[45]), .B1_f (plaintext_s1_f[45]), .Z0_t (RoundReg_Inst_ff_SDE_45_MUX_inst_X), .Z0_f (new_AGEMA_signal_18068), .Z1_t (new_AGEMA_signal_18069), .Z1_f (new_AGEMA_signal_18070) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_45_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_45_MUX_inst_X), .B0_f (new_AGEMA_signal_18068), .B1_t (new_AGEMA_signal_18069), .B1_f (new_AGEMA_signal_18070), .Z0_t (RoundReg_Inst_ff_SDE_45_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18593), .Z1_t (new_AGEMA_signal_18594), .Z1_f (new_AGEMA_signal_18595) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_45_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_45_MUX_inst_Y), .A0_f (new_AGEMA_signal_18593), .A1_t (new_AGEMA_signal_18594), .A1_f (new_AGEMA_signal_18595), .B0_t (RoundOutput[45]), .B0_f (new_AGEMA_signal_17447), .B1_t (new_AGEMA_signal_17448), .B1_f (new_AGEMA_signal_17449), .Z0_t (RoundInput[45]), .Z0_f (new_AGEMA_signal_5663), .Z1_t (new_AGEMA_signal_5664), .Z1_f (new_AGEMA_signal_5665) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_46_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[46]), .A0_f (new_AGEMA_signal_17450), .A1_t (new_AGEMA_signal_17451), .A1_f (new_AGEMA_signal_17452), .B0_t (plaintext_s0_t[46]), .B0_f (plaintext_s0_f[46]), .B1_t (plaintext_s1_t[46]), .B1_f (plaintext_s1_f[46]), .Z0_t (RoundReg_Inst_ff_SDE_46_MUX_inst_X), .Z0_f (new_AGEMA_signal_18074), .Z1_t (new_AGEMA_signal_18075), .Z1_f (new_AGEMA_signal_18076) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_46_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_46_MUX_inst_X), .B0_f (new_AGEMA_signal_18074), .B1_t (new_AGEMA_signal_18075), .B1_f (new_AGEMA_signal_18076), .Z0_t (RoundReg_Inst_ff_SDE_46_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18596), .Z1_t (new_AGEMA_signal_18597), .Z1_f (new_AGEMA_signal_18598) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_46_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_46_MUX_inst_Y), .A0_f (new_AGEMA_signal_18596), .A1_t (new_AGEMA_signal_18597), .A1_f (new_AGEMA_signal_18598), .B0_t (RoundOutput[46]), .B0_f (new_AGEMA_signal_17450), .B1_t (new_AGEMA_signal_17451), .B1_f (new_AGEMA_signal_17452), .Z0_t (RoundInput[46]), .Z0_f (new_AGEMA_signal_5672), .Z1_t (new_AGEMA_signal_5673), .Z1_f (new_AGEMA_signal_5674) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_47_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[47]), .A0_f (new_AGEMA_signal_17453), .A1_t (new_AGEMA_signal_17454), .A1_f (new_AGEMA_signal_17455), .B0_t (plaintext_s0_t[47]), .B0_f (plaintext_s0_f[47]), .B1_t (plaintext_s1_t[47]), .B1_f (plaintext_s1_f[47]), .Z0_t (RoundReg_Inst_ff_SDE_47_MUX_inst_X), .Z0_f (new_AGEMA_signal_18080), .Z1_t (new_AGEMA_signal_18081), .Z1_f (new_AGEMA_signal_18082) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_47_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_47_MUX_inst_X), .B0_f (new_AGEMA_signal_18080), .B1_t (new_AGEMA_signal_18081), .B1_f (new_AGEMA_signal_18082), .Z0_t (RoundReg_Inst_ff_SDE_47_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18599), .Z1_t (new_AGEMA_signal_18600), .Z1_f (new_AGEMA_signal_18601) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_47_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_47_MUX_inst_Y), .A0_f (new_AGEMA_signal_18599), .A1_t (new_AGEMA_signal_18600), .A1_f (new_AGEMA_signal_18601), .B0_t (RoundOutput[47]), .B0_f (new_AGEMA_signal_17453), .B1_t (new_AGEMA_signal_17454), .B1_f (new_AGEMA_signal_17455), .Z0_t (RoundInput[47]), .Z0_f (new_AGEMA_signal_5681), .Z1_t (new_AGEMA_signal_5682), .Z1_f (new_AGEMA_signal_5683) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_48_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[48]), .A0_f (new_AGEMA_signal_17456), .A1_t (new_AGEMA_signal_17457), .A1_f (new_AGEMA_signal_17458), .B0_t (plaintext_s0_t[48]), .B0_f (plaintext_s0_f[48]), .B1_t (plaintext_s1_t[48]), .B1_f (plaintext_s1_f[48]), .Z0_t (RoundReg_Inst_ff_SDE_48_MUX_inst_X), .Z0_f (new_AGEMA_signal_18086), .Z1_t (new_AGEMA_signal_18087), .Z1_f (new_AGEMA_signal_18088) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_48_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_48_MUX_inst_X), .B0_f (new_AGEMA_signal_18086), .B1_t (new_AGEMA_signal_18087), .B1_f (new_AGEMA_signal_18088), .Z0_t (RoundReg_Inst_ff_SDE_48_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18602), .Z1_t (new_AGEMA_signal_18603), .Z1_f (new_AGEMA_signal_18604) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_48_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_48_MUX_inst_Y), .A0_f (new_AGEMA_signal_18602), .A1_t (new_AGEMA_signal_18603), .A1_f (new_AGEMA_signal_18604), .B0_t (RoundOutput[48]), .B0_f (new_AGEMA_signal_17456), .B1_t (new_AGEMA_signal_17457), .B1_f (new_AGEMA_signal_17458), .Z0_t (RoundInput[48]), .Z0_f (new_AGEMA_signal_5690), .Z1_t (new_AGEMA_signal_5691), .Z1_f (new_AGEMA_signal_5692) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_49_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[49]), .A0_f (new_AGEMA_signal_17837), .A1_t (new_AGEMA_signal_17838), .A1_f (new_AGEMA_signal_17839), .B0_t (plaintext_s0_t[49]), .B0_f (plaintext_s0_f[49]), .B1_t (plaintext_s1_t[49]), .B1_f (plaintext_s1_f[49]), .Z0_t (RoundReg_Inst_ff_SDE_49_MUX_inst_X), .Z0_f (new_AGEMA_signal_18608), .Z1_t (new_AGEMA_signal_18609), .Z1_f (new_AGEMA_signal_18610) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_49_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_49_MUX_inst_X), .B0_f (new_AGEMA_signal_18608), .B1_t (new_AGEMA_signal_18609), .B1_f (new_AGEMA_signal_18610), .Z0_t (RoundReg_Inst_ff_SDE_49_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18986), .Z1_t (new_AGEMA_signal_18987), .Z1_f (new_AGEMA_signal_18988) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_49_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_49_MUX_inst_Y), .A0_f (new_AGEMA_signal_18986), .A1_t (new_AGEMA_signal_18987), .A1_f (new_AGEMA_signal_18988), .B0_t (RoundOutput[49]), .B0_f (new_AGEMA_signal_17837), .B1_t (new_AGEMA_signal_17838), .B1_f (new_AGEMA_signal_17839), .Z0_t (RoundInput[49]), .Z0_f (new_AGEMA_signal_5699), .Z1_t (new_AGEMA_signal_5700), .Z1_f (new_AGEMA_signal_5701) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_50_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[50]), .A0_f (new_AGEMA_signal_17465), .A1_t (new_AGEMA_signal_17466), .A1_f (new_AGEMA_signal_17467), .B0_t (plaintext_s0_t[50]), .B0_f (plaintext_s0_f[50]), .B1_t (plaintext_s1_t[50]), .B1_f (plaintext_s1_f[50]), .Z0_t (RoundReg_Inst_ff_SDE_50_MUX_inst_X), .Z0_f (new_AGEMA_signal_18092), .Z1_t (new_AGEMA_signal_18093), .Z1_f (new_AGEMA_signal_18094) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_50_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_50_MUX_inst_X), .B0_f (new_AGEMA_signal_18092), .B1_t (new_AGEMA_signal_18093), .B1_f (new_AGEMA_signal_18094), .Z0_t (RoundReg_Inst_ff_SDE_50_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18611), .Z1_t (new_AGEMA_signal_18612), .Z1_f (new_AGEMA_signal_18613) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_50_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_50_MUX_inst_Y), .A0_f (new_AGEMA_signal_18611), .A1_t (new_AGEMA_signal_18612), .A1_f (new_AGEMA_signal_18613), .B0_t (RoundOutput[50]), .B0_f (new_AGEMA_signal_17465), .B1_t (new_AGEMA_signal_17466), .B1_f (new_AGEMA_signal_17467), .Z0_t (RoundInput[50]), .Z0_f (new_AGEMA_signal_5717), .Z1_t (new_AGEMA_signal_5718), .Z1_f (new_AGEMA_signal_5719) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_51_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[51]), .A0_f (new_AGEMA_signal_17843), .A1_t (new_AGEMA_signal_17844), .A1_f (new_AGEMA_signal_17845), .B0_t (plaintext_s0_t[51]), .B0_f (plaintext_s0_f[51]), .B1_t (plaintext_s1_t[51]), .B1_f (plaintext_s1_f[51]), .Z0_t (RoundReg_Inst_ff_SDE_51_MUX_inst_X), .Z0_f (new_AGEMA_signal_18617), .Z1_t (new_AGEMA_signal_18618), .Z1_f (new_AGEMA_signal_18619) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_51_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_51_MUX_inst_X), .B0_f (new_AGEMA_signal_18617), .B1_t (new_AGEMA_signal_18618), .B1_f (new_AGEMA_signal_18619), .Z0_t (RoundReg_Inst_ff_SDE_51_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18989), .Z1_t (new_AGEMA_signal_18990), .Z1_f (new_AGEMA_signal_18991) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_51_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_51_MUX_inst_Y), .A0_f (new_AGEMA_signal_18989), .A1_t (new_AGEMA_signal_18990), .A1_f (new_AGEMA_signal_18991), .B0_t (RoundOutput[51]), .B0_f (new_AGEMA_signal_17843), .B1_t (new_AGEMA_signal_17844), .B1_f (new_AGEMA_signal_17845), .Z0_t (RoundInput[51]), .Z0_f (new_AGEMA_signal_5726), .Z1_t (new_AGEMA_signal_5727), .Z1_f (new_AGEMA_signal_5728) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_52_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[52]), .A0_f (new_AGEMA_signal_17846), .A1_t (new_AGEMA_signal_17847), .A1_f (new_AGEMA_signal_17848), .B0_t (plaintext_s0_t[52]), .B0_f (plaintext_s0_f[52]), .B1_t (plaintext_s1_t[52]), .B1_f (plaintext_s1_f[52]), .Z0_t (RoundReg_Inst_ff_SDE_52_MUX_inst_X), .Z0_f (new_AGEMA_signal_18623), .Z1_t (new_AGEMA_signal_18624), .Z1_f (new_AGEMA_signal_18625) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_52_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_52_MUX_inst_X), .B0_f (new_AGEMA_signal_18623), .B1_t (new_AGEMA_signal_18624), .B1_f (new_AGEMA_signal_18625), .Z0_t (RoundReg_Inst_ff_SDE_52_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18992), .Z1_t (new_AGEMA_signal_18993), .Z1_f (new_AGEMA_signal_18994) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_52_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_52_MUX_inst_Y), .A0_f (new_AGEMA_signal_18992), .A1_t (new_AGEMA_signal_18993), .A1_f (new_AGEMA_signal_18994), .B0_t (RoundOutput[52]), .B0_f (new_AGEMA_signal_17846), .B1_t (new_AGEMA_signal_17847), .B1_f (new_AGEMA_signal_17848), .Z0_t (RoundInput[52]), .Z0_f (new_AGEMA_signal_5735), .Z1_t (new_AGEMA_signal_5736), .Z1_f (new_AGEMA_signal_5737) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_53_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[53]), .A0_f (new_AGEMA_signal_17474), .A1_t (new_AGEMA_signal_17475), .A1_f (new_AGEMA_signal_17476), .B0_t (plaintext_s0_t[53]), .B0_f (plaintext_s0_f[53]), .B1_t (plaintext_s1_t[53]), .B1_f (plaintext_s1_f[53]), .Z0_t (RoundReg_Inst_ff_SDE_53_MUX_inst_X), .Z0_f (new_AGEMA_signal_18098), .Z1_t (new_AGEMA_signal_18099), .Z1_f (new_AGEMA_signal_18100) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_53_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_53_MUX_inst_X), .B0_f (new_AGEMA_signal_18098), .B1_t (new_AGEMA_signal_18099), .B1_f (new_AGEMA_signal_18100), .Z0_t (RoundReg_Inst_ff_SDE_53_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18626), .Z1_t (new_AGEMA_signal_18627), .Z1_f (new_AGEMA_signal_18628) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_53_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_53_MUX_inst_Y), .A0_f (new_AGEMA_signal_18626), .A1_t (new_AGEMA_signal_18627), .A1_f (new_AGEMA_signal_18628), .B0_t (RoundOutput[53]), .B0_f (new_AGEMA_signal_17474), .B1_t (new_AGEMA_signal_17475), .B1_f (new_AGEMA_signal_17476), .Z0_t (RoundInput[53]), .Z0_f (new_AGEMA_signal_5744), .Z1_t (new_AGEMA_signal_5745), .Z1_f (new_AGEMA_signal_5746) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_54_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[54]), .A0_f (new_AGEMA_signal_17477), .A1_t (new_AGEMA_signal_17478), .A1_f (new_AGEMA_signal_17479), .B0_t (plaintext_s0_t[54]), .B0_f (plaintext_s0_f[54]), .B1_t (plaintext_s1_t[54]), .B1_f (plaintext_s1_f[54]), .Z0_t (RoundReg_Inst_ff_SDE_54_MUX_inst_X), .Z0_f (new_AGEMA_signal_18104), .Z1_t (new_AGEMA_signal_18105), .Z1_f (new_AGEMA_signal_18106) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_54_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_54_MUX_inst_X), .B0_f (new_AGEMA_signal_18104), .B1_t (new_AGEMA_signal_18105), .B1_f (new_AGEMA_signal_18106), .Z0_t (RoundReg_Inst_ff_SDE_54_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18629), .Z1_t (new_AGEMA_signal_18630), .Z1_f (new_AGEMA_signal_18631) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_54_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_54_MUX_inst_Y), .A0_f (new_AGEMA_signal_18629), .A1_t (new_AGEMA_signal_18630), .A1_f (new_AGEMA_signal_18631), .B0_t (RoundOutput[54]), .B0_f (new_AGEMA_signal_17477), .B1_t (new_AGEMA_signal_17478), .B1_f (new_AGEMA_signal_17479), .Z0_t (RoundInput[54]), .Z0_f (new_AGEMA_signal_5753), .Z1_t (new_AGEMA_signal_5754), .Z1_f (new_AGEMA_signal_5755) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_55_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[55]), .A0_f (new_AGEMA_signal_17480), .A1_t (new_AGEMA_signal_17481), .A1_f (new_AGEMA_signal_17482), .B0_t (plaintext_s0_t[55]), .B0_f (plaintext_s0_f[55]), .B1_t (plaintext_s1_t[55]), .B1_f (plaintext_s1_f[55]), .Z0_t (RoundReg_Inst_ff_SDE_55_MUX_inst_X), .Z0_f (new_AGEMA_signal_18110), .Z1_t (new_AGEMA_signal_18111), .Z1_f (new_AGEMA_signal_18112) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_55_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_55_MUX_inst_X), .B0_f (new_AGEMA_signal_18110), .B1_t (new_AGEMA_signal_18111), .B1_f (new_AGEMA_signal_18112), .Z0_t (RoundReg_Inst_ff_SDE_55_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18632), .Z1_t (new_AGEMA_signal_18633), .Z1_f (new_AGEMA_signal_18634) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_55_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_55_MUX_inst_Y), .A0_f (new_AGEMA_signal_18632), .A1_t (new_AGEMA_signal_18633), .A1_f (new_AGEMA_signal_18634), .B0_t (RoundOutput[55]), .B0_f (new_AGEMA_signal_17480), .B1_t (new_AGEMA_signal_17481), .B1_f (new_AGEMA_signal_17482), .Z0_t (RoundInput[55]), .Z0_f (new_AGEMA_signal_5762), .Z1_t (new_AGEMA_signal_5763), .Z1_f (new_AGEMA_signal_5764) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_56_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[56]), .A0_f (new_AGEMA_signal_17483), .A1_t (new_AGEMA_signal_17484), .A1_f (new_AGEMA_signal_17485), .B0_t (plaintext_s0_t[56]), .B0_f (plaintext_s0_f[56]), .B1_t (plaintext_s1_t[56]), .B1_f (plaintext_s1_f[56]), .Z0_t (RoundReg_Inst_ff_SDE_56_MUX_inst_X), .Z0_f (new_AGEMA_signal_18116), .Z1_t (new_AGEMA_signal_18117), .Z1_f (new_AGEMA_signal_18118) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_56_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_56_MUX_inst_X), .B0_f (new_AGEMA_signal_18116), .B1_t (new_AGEMA_signal_18117), .B1_f (new_AGEMA_signal_18118), .Z0_t (RoundReg_Inst_ff_SDE_56_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18635), .Z1_t (new_AGEMA_signal_18636), .Z1_f (new_AGEMA_signal_18637) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_56_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_56_MUX_inst_Y), .A0_f (new_AGEMA_signal_18635), .A1_t (new_AGEMA_signal_18636), .A1_f (new_AGEMA_signal_18637), .B0_t (RoundOutput[56]), .B0_f (new_AGEMA_signal_17483), .B1_t (new_AGEMA_signal_17484), .B1_f (new_AGEMA_signal_17485), .Z0_t (RoundInput[56]), .Z0_f (new_AGEMA_signal_5771), .Z1_t (new_AGEMA_signal_5772), .Z1_f (new_AGEMA_signal_5773) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_57_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[57]), .A0_f (new_AGEMA_signal_17849), .A1_t (new_AGEMA_signal_17850), .A1_f (new_AGEMA_signal_17851), .B0_t (plaintext_s0_t[57]), .B0_f (plaintext_s0_f[57]), .B1_t (plaintext_s1_t[57]), .B1_f (plaintext_s1_f[57]), .Z0_t (RoundReg_Inst_ff_SDE_57_MUX_inst_X), .Z0_f (new_AGEMA_signal_18641), .Z1_t (new_AGEMA_signal_18642), .Z1_f (new_AGEMA_signal_18643) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_57_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_57_MUX_inst_X), .B0_f (new_AGEMA_signal_18641), .B1_t (new_AGEMA_signal_18642), .B1_f (new_AGEMA_signal_18643), .Z0_t (RoundReg_Inst_ff_SDE_57_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18995), .Z1_t (new_AGEMA_signal_18996), .Z1_f (new_AGEMA_signal_18997) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_57_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_57_MUX_inst_Y), .A0_f (new_AGEMA_signal_18995), .A1_t (new_AGEMA_signal_18996), .A1_f (new_AGEMA_signal_18997), .B0_t (RoundOutput[57]), .B0_f (new_AGEMA_signal_17849), .B1_t (new_AGEMA_signal_17850), .B1_f (new_AGEMA_signal_17851), .Z0_t (RoundInput[57]), .Z0_f (new_AGEMA_signal_5780), .Z1_t (new_AGEMA_signal_5781), .Z1_f (new_AGEMA_signal_5782) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_58_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[58]), .A0_f (new_AGEMA_signal_17489), .A1_t (new_AGEMA_signal_17490), .A1_f (new_AGEMA_signal_17491), .B0_t (plaintext_s0_t[58]), .B0_f (plaintext_s0_f[58]), .B1_t (plaintext_s1_t[58]), .B1_f (plaintext_s1_f[58]), .Z0_t (RoundReg_Inst_ff_SDE_58_MUX_inst_X), .Z0_f (new_AGEMA_signal_18122), .Z1_t (new_AGEMA_signal_18123), .Z1_f (new_AGEMA_signal_18124) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_58_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_58_MUX_inst_X), .B0_f (new_AGEMA_signal_18122), .B1_t (new_AGEMA_signal_18123), .B1_f (new_AGEMA_signal_18124), .Z0_t (RoundReg_Inst_ff_SDE_58_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18644), .Z1_t (new_AGEMA_signal_18645), .Z1_f (new_AGEMA_signal_18646) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_58_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_58_MUX_inst_Y), .A0_f (new_AGEMA_signal_18644), .A1_t (new_AGEMA_signal_18645), .A1_f (new_AGEMA_signal_18646), .B0_t (RoundOutput[58]), .B0_f (new_AGEMA_signal_17489), .B1_t (new_AGEMA_signal_17490), .B1_f (new_AGEMA_signal_17491), .Z0_t (RoundInput[58]), .Z0_f (new_AGEMA_signal_5789), .Z1_t (new_AGEMA_signal_5790), .Z1_f (new_AGEMA_signal_5791) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_59_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[59]), .A0_f (new_AGEMA_signal_17852), .A1_t (new_AGEMA_signal_17853), .A1_f (new_AGEMA_signal_17854), .B0_t (plaintext_s0_t[59]), .B0_f (plaintext_s0_f[59]), .B1_t (plaintext_s1_t[59]), .B1_f (plaintext_s1_f[59]), .Z0_t (RoundReg_Inst_ff_SDE_59_MUX_inst_X), .Z0_f (new_AGEMA_signal_18650), .Z1_t (new_AGEMA_signal_18651), .Z1_f (new_AGEMA_signal_18652) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_59_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_59_MUX_inst_X), .B0_f (new_AGEMA_signal_18650), .B1_t (new_AGEMA_signal_18651), .B1_f (new_AGEMA_signal_18652), .Z0_t (RoundReg_Inst_ff_SDE_59_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18998), .Z1_t (new_AGEMA_signal_18999), .Z1_f (new_AGEMA_signal_19000) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_59_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_59_MUX_inst_Y), .A0_f (new_AGEMA_signal_18998), .A1_t (new_AGEMA_signal_18999), .A1_f (new_AGEMA_signal_19000), .B0_t (RoundOutput[59]), .B0_f (new_AGEMA_signal_17852), .B1_t (new_AGEMA_signal_17853), .B1_f (new_AGEMA_signal_17854), .Z0_t (RoundInput[59]), .Z0_f (new_AGEMA_signal_5798), .Z1_t (new_AGEMA_signal_5799), .Z1_f (new_AGEMA_signal_5800) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_60_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[60]), .A0_f (new_AGEMA_signal_17855), .A1_t (new_AGEMA_signal_17856), .A1_f (new_AGEMA_signal_17857), .B0_t (plaintext_s0_t[60]), .B0_f (plaintext_s0_f[60]), .B1_t (plaintext_s1_t[60]), .B1_f (plaintext_s1_f[60]), .Z0_t (RoundReg_Inst_ff_SDE_60_MUX_inst_X), .Z0_f (new_AGEMA_signal_18656), .Z1_t (new_AGEMA_signal_18657), .Z1_f (new_AGEMA_signal_18658) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_60_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_60_MUX_inst_X), .B0_f (new_AGEMA_signal_18656), .B1_t (new_AGEMA_signal_18657), .B1_f (new_AGEMA_signal_18658), .Z0_t (RoundReg_Inst_ff_SDE_60_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19001), .Z1_t (new_AGEMA_signal_19002), .Z1_f (new_AGEMA_signal_19003) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_60_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_60_MUX_inst_Y), .A0_f (new_AGEMA_signal_19001), .A1_t (new_AGEMA_signal_19002), .A1_f (new_AGEMA_signal_19003), .B0_t (RoundOutput[60]), .B0_f (new_AGEMA_signal_17855), .B1_t (new_AGEMA_signal_17856), .B1_f (new_AGEMA_signal_17857), .Z0_t (RoundInput[60]), .Z0_f (new_AGEMA_signal_5816), .Z1_t (new_AGEMA_signal_5817), .Z1_f (new_AGEMA_signal_5818) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_61_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[61]), .A0_f (new_AGEMA_signal_17501), .A1_t (new_AGEMA_signal_17502), .A1_f (new_AGEMA_signal_17503), .B0_t (plaintext_s0_t[61]), .B0_f (plaintext_s0_f[61]), .B1_t (plaintext_s1_t[61]), .B1_f (plaintext_s1_f[61]), .Z0_t (RoundReg_Inst_ff_SDE_61_MUX_inst_X), .Z0_f (new_AGEMA_signal_18128), .Z1_t (new_AGEMA_signal_18129), .Z1_f (new_AGEMA_signal_18130) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_61_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_61_MUX_inst_X), .B0_f (new_AGEMA_signal_18128), .B1_t (new_AGEMA_signal_18129), .B1_f (new_AGEMA_signal_18130), .Z0_t (RoundReg_Inst_ff_SDE_61_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18659), .Z1_t (new_AGEMA_signal_18660), .Z1_f (new_AGEMA_signal_18661) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_61_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_61_MUX_inst_Y), .A0_f (new_AGEMA_signal_18659), .A1_t (new_AGEMA_signal_18660), .A1_f (new_AGEMA_signal_18661), .B0_t (RoundOutput[61]), .B0_f (new_AGEMA_signal_17501), .B1_t (new_AGEMA_signal_17502), .B1_f (new_AGEMA_signal_17503), .Z0_t (RoundInput[61]), .Z0_f (new_AGEMA_signal_5825), .Z1_t (new_AGEMA_signal_5826), .Z1_f (new_AGEMA_signal_5827) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_62_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[62]), .A0_f (new_AGEMA_signal_17504), .A1_t (new_AGEMA_signal_17505), .A1_f (new_AGEMA_signal_17506), .B0_t (plaintext_s0_t[62]), .B0_f (plaintext_s0_f[62]), .B1_t (plaintext_s1_t[62]), .B1_f (plaintext_s1_f[62]), .Z0_t (RoundReg_Inst_ff_SDE_62_MUX_inst_X), .Z0_f (new_AGEMA_signal_18134), .Z1_t (new_AGEMA_signal_18135), .Z1_f (new_AGEMA_signal_18136) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_62_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_62_MUX_inst_X), .B0_f (new_AGEMA_signal_18134), .B1_t (new_AGEMA_signal_18135), .B1_f (new_AGEMA_signal_18136), .Z0_t (RoundReg_Inst_ff_SDE_62_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18662), .Z1_t (new_AGEMA_signal_18663), .Z1_f (new_AGEMA_signal_18664) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_62_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_62_MUX_inst_Y), .A0_f (new_AGEMA_signal_18662), .A1_t (new_AGEMA_signal_18663), .A1_f (new_AGEMA_signal_18664), .B0_t (RoundOutput[62]), .B0_f (new_AGEMA_signal_17504), .B1_t (new_AGEMA_signal_17505), .B1_f (new_AGEMA_signal_17506), .Z0_t (RoundInput[62]), .Z0_f (new_AGEMA_signal_5834), .Z1_t (new_AGEMA_signal_5835), .Z1_f (new_AGEMA_signal_5836) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_63_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[63]), .A0_f (new_AGEMA_signal_17507), .A1_t (new_AGEMA_signal_17508), .A1_f (new_AGEMA_signal_17509), .B0_t (plaintext_s0_t[63]), .B0_f (plaintext_s0_f[63]), .B1_t (plaintext_s1_t[63]), .B1_f (plaintext_s1_f[63]), .Z0_t (RoundReg_Inst_ff_SDE_63_MUX_inst_X), .Z0_f (new_AGEMA_signal_18140), .Z1_t (new_AGEMA_signal_18141), .Z1_f (new_AGEMA_signal_18142) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_63_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_63_MUX_inst_X), .B0_f (new_AGEMA_signal_18140), .B1_t (new_AGEMA_signal_18141), .B1_f (new_AGEMA_signal_18142), .Z0_t (RoundReg_Inst_ff_SDE_63_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18665), .Z1_t (new_AGEMA_signal_18666), .Z1_f (new_AGEMA_signal_18667) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_63_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_63_MUX_inst_Y), .A0_f (new_AGEMA_signal_18665), .A1_t (new_AGEMA_signal_18666), .A1_f (new_AGEMA_signal_18667), .B0_t (RoundOutput[63]), .B0_f (new_AGEMA_signal_17507), .B1_t (new_AGEMA_signal_17508), .B1_f (new_AGEMA_signal_17509), .Z0_t (RoundInput[63]), .Z0_f (new_AGEMA_signal_5843), .Z1_t (new_AGEMA_signal_5844), .Z1_f (new_AGEMA_signal_5845) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_64_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[64]), .A0_f (new_AGEMA_signal_17510), .A1_t (new_AGEMA_signal_17511), .A1_f (new_AGEMA_signal_17512), .B0_t (plaintext_s0_t[64]), .B0_f (plaintext_s0_f[64]), .B1_t (plaintext_s1_t[64]), .B1_f (plaintext_s1_f[64]), .Z0_t (RoundReg_Inst_ff_SDE_64_MUX_inst_X), .Z0_f (new_AGEMA_signal_18146), .Z1_t (new_AGEMA_signal_18147), .Z1_f (new_AGEMA_signal_18148) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_64_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_64_MUX_inst_X), .B0_f (new_AGEMA_signal_18146), .B1_t (new_AGEMA_signal_18147), .B1_f (new_AGEMA_signal_18148), .Z0_t (RoundReg_Inst_ff_SDE_64_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18668), .Z1_t (new_AGEMA_signal_18669), .Z1_f (new_AGEMA_signal_18670) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_64_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_64_MUX_inst_Y), .A0_f (new_AGEMA_signal_18668), .A1_t (new_AGEMA_signal_18669), .A1_f (new_AGEMA_signal_18670), .B0_t (RoundOutput[64]), .B0_f (new_AGEMA_signal_17510), .B1_t (new_AGEMA_signal_17511), .B1_f (new_AGEMA_signal_17512), .Z0_t (RoundInput[64]), .Z0_f (new_AGEMA_signal_5852), .Z1_t (new_AGEMA_signal_5853), .Z1_f (new_AGEMA_signal_5854) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_65_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[65]), .A0_f (new_AGEMA_signal_17858), .A1_t (new_AGEMA_signal_17859), .A1_f (new_AGEMA_signal_17860), .B0_t (plaintext_s0_t[65]), .B0_f (plaintext_s0_f[65]), .B1_t (plaintext_s1_t[65]), .B1_f (plaintext_s1_f[65]), .Z0_t (RoundReg_Inst_ff_SDE_65_MUX_inst_X), .Z0_f (new_AGEMA_signal_18674), .Z1_t (new_AGEMA_signal_18675), .Z1_f (new_AGEMA_signal_18676) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_65_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_65_MUX_inst_X), .B0_f (new_AGEMA_signal_18674), .B1_t (new_AGEMA_signal_18675), .B1_f (new_AGEMA_signal_18676), .Z0_t (RoundReg_Inst_ff_SDE_65_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19004), .Z1_t (new_AGEMA_signal_19005), .Z1_f (new_AGEMA_signal_19006) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_65_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_65_MUX_inst_Y), .A0_f (new_AGEMA_signal_19004), .A1_t (new_AGEMA_signal_19005), .A1_f (new_AGEMA_signal_19006), .B0_t (RoundOutput[65]), .B0_f (new_AGEMA_signal_17858), .B1_t (new_AGEMA_signal_17859), .B1_f (new_AGEMA_signal_17860), .Z0_t (RoundInput[65]), .Z0_f (new_AGEMA_signal_5861), .Z1_t (new_AGEMA_signal_5862), .Z1_f (new_AGEMA_signal_5863) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_66_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[66]), .A0_f (new_AGEMA_signal_17516), .A1_t (new_AGEMA_signal_17517), .A1_f (new_AGEMA_signal_17518), .B0_t (plaintext_s0_t[66]), .B0_f (plaintext_s0_f[66]), .B1_t (plaintext_s1_t[66]), .B1_f (plaintext_s1_f[66]), .Z0_t (RoundReg_Inst_ff_SDE_66_MUX_inst_X), .Z0_f (new_AGEMA_signal_18152), .Z1_t (new_AGEMA_signal_18153), .Z1_f (new_AGEMA_signal_18154) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_66_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_66_MUX_inst_X), .B0_f (new_AGEMA_signal_18152), .B1_t (new_AGEMA_signal_18153), .B1_f (new_AGEMA_signal_18154), .Z0_t (RoundReg_Inst_ff_SDE_66_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18677), .Z1_t (new_AGEMA_signal_18678), .Z1_f (new_AGEMA_signal_18679) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_66_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_66_MUX_inst_Y), .A0_f (new_AGEMA_signal_18677), .A1_t (new_AGEMA_signal_18678), .A1_f (new_AGEMA_signal_18679), .B0_t (RoundOutput[66]), .B0_f (new_AGEMA_signal_17516), .B1_t (new_AGEMA_signal_17517), .B1_f (new_AGEMA_signal_17518), .Z0_t (RoundInput[66]), .Z0_f (new_AGEMA_signal_5870), .Z1_t (new_AGEMA_signal_5871), .Z1_f (new_AGEMA_signal_5872) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_67_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[67]), .A0_f (new_AGEMA_signal_17861), .A1_t (new_AGEMA_signal_17862), .A1_f (new_AGEMA_signal_17863), .B0_t (plaintext_s0_t[67]), .B0_f (plaintext_s0_f[67]), .B1_t (plaintext_s1_t[67]), .B1_f (plaintext_s1_f[67]), .Z0_t (RoundReg_Inst_ff_SDE_67_MUX_inst_X), .Z0_f (new_AGEMA_signal_18683), .Z1_t (new_AGEMA_signal_18684), .Z1_f (new_AGEMA_signal_18685) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_67_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_67_MUX_inst_X), .B0_f (new_AGEMA_signal_18683), .B1_t (new_AGEMA_signal_18684), .B1_f (new_AGEMA_signal_18685), .Z0_t (RoundReg_Inst_ff_SDE_67_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19007), .Z1_t (new_AGEMA_signal_19008), .Z1_f (new_AGEMA_signal_19009) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_67_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_67_MUX_inst_Y), .A0_f (new_AGEMA_signal_19007), .A1_t (new_AGEMA_signal_19008), .A1_f (new_AGEMA_signal_19009), .B0_t (RoundOutput[67]), .B0_f (new_AGEMA_signal_17861), .B1_t (new_AGEMA_signal_17862), .B1_f (new_AGEMA_signal_17863), .Z0_t (RoundInput[67]), .Z0_f (new_AGEMA_signal_5879), .Z1_t (new_AGEMA_signal_5880), .Z1_f (new_AGEMA_signal_5881) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_68_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[68]), .A0_f (new_AGEMA_signal_17864), .A1_t (new_AGEMA_signal_17865), .A1_f (new_AGEMA_signal_17866), .B0_t (plaintext_s0_t[68]), .B0_f (plaintext_s0_f[68]), .B1_t (plaintext_s1_t[68]), .B1_f (plaintext_s1_f[68]), .Z0_t (RoundReg_Inst_ff_SDE_68_MUX_inst_X), .Z0_f (new_AGEMA_signal_18689), .Z1_t (new_AGEMA_signal_18690), .Z1_f (new_AGEMA_signal_18691) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_68_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_68_MUX_inst_X), .B0_f (new_AGEMA_signal_18689), .B1_t (new_AGEMA_signal_18690), .B1_f (new_AGEMA_signal_18691), .Z0_t (RoundReg_Inst_ff_SDE_68_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19010), .Z1_t (new_AGEMA_signal_19011), .Z1_f (new_AGEMA_signal_19012) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_68_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_68_MUX_inst_Y), .A0_f (new_AGEMA_signal_19010), .A1_t (new_AGEMA_signal_19011), .A1_f (new_AGEMA_signal_19012), .B0_t (RoundOutput[68]), .B0_f (new_AGEMA_signal_17864), .B1_t (new_AGEMA_signal_17865), .B1_f (new_AGEMA_signal_17866), .Z0_t (RoundInput[68]), .Z0_f (new_AGEMA_signal_5888), .Z1_t (new_AGEMA_signal_5889), .Z1_f (new_AGEMA_signal_5890) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_69_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[69]), .A0_f (new_AGEMA_signal_17525), .A1_t (new_AGEMA_signal_17526), .A1_f (new_AGEMA_signal_17527), .B0_t (plaintext_s0_t[69]), .B0_f (plaintext_s0_f[69]), .B1_t (plaintext_s1_t[69]), .B1_f (plaintext_s1_f[69]), .Z0_t (RoundReg_Inst_ff_SDE_69_MUX_inst_X), .Z0_f (new_AGEMA_signal_18158), .Z1_t (new_AGEMA_signal_18159), .Z1_f (new_AGEMA_signal_18160) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_69_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_69_MUX_inst_X), .B0_f (new_AGEMA_signal_18158), .B1_t (new_AGEMA_signal_18159), .B1_f (new_AGEMA_signal_18160), .Z0_t (RoundReg_Inst_ff_SDE_69_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18692), .Z1_t (new_AGEMA_signal_18693), .Z1_f (new_AGEMA_signal_18694) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_69_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_69_MUX_inst_Y), .A0_f (new_AGEMA_signal_18692), .A1_t (new_AGEMA_signal_18693), .A1_f (new_AGEMA_signal_18694), .B0_t (RoundOutput[69]), .B0_f (new_AGEMA_signal_17525), .B1_t (new_AGEMA_signal_17526), .B1_f (new_AGEMA_signal_17527), .Z0_t (RoundInput[69]), .Z0_f (new_AGEMA_signal_5897), .Z1_t (new_AGEMA_signal_5898), .Z1_f (new_AGEMA_signal_5899) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_70_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[70]), .A0_f (new_AGEMA_signal_17531), .A1_t (new_AGEMA_signal_17532), .A1_f (new_AGEMA_signal_17533), .B0_t (plaintext_s0_t[70]), .B0_f (plaintext_s0_f[70]), .B1_t (plaintext_s1_t[70]), .B1_f (plaintext_s1_f[70]), .Z0_t (RoundReg_Inst_ff_SDE_70_MUX_inst_X), .Z0_f (new_AGEMA_signal_18164), .Z1_t (new_AGEMA_signal_18165), .Z1_f (new_AGEMA_signal_18166) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_70_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_70_MUX_inst_X), .B0_f (new_AGEMA_signal_18164), .B1_t (new_AGEMA_signal_18165), .B1_f (new_AGEMA_signal_18166), .Z0_t (RoundReg_Inst_ff_SDE_70_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18695), .Z1_t (new_AGEMA_signal_18696), .Z1_f (new_AGEMA_signal_18697) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_70_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_70_MUX_inst_Y), .A0_f (new_AGEMA_signal_18695), .A1_t (new_AGEMA_signal_18696), .A1_f (new_AGEMA_signal_18697), .B0_t (RoundOutput[70]), .B0_f (new_AGEMA_signal_17531), .B1_t (new_AGEMA_signal_17532), .B1_f (new_AGEMA_signal_17533), .Z0_t (RoundInput[70]), .Z0_f (new_AGEMA_signal_5915), .Z1_t (new_AGEMA_signal_5916), .Z1_f (new_AGEMA_signal_5917) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_71_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[71]), .A0_f (new_AGEMA_signal_17534), .A1_t (new_AGEMA_signal_17535), .A1_f (new_AGEMA_signal_17536), .B0_t (plaintext_s0_t[71]), .B0_f (plaintext_s0_f[71]), .B1_t (plaintext_s1_t[71]), .B1_f (plaintext_s1_f[71]), .Z0_t (RoundReg_Inst_ff_SDE_71_MUX_inst_X), .Z0_f (new_AGEMA_signal_18170), .Z1_t (new_AGEMA_signal_18171), .Z1_f (new_AGEMA_signal_18172) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_71_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_71_MUX_inst_X), .B0_f (new_AGEMA_signal_18170), .B1_t (new_AGEMA_signal_18171), .B1_f (new_AGEMA_signal_18172), .Z0_t (RoundReg_Inst_ff_SDE_71_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18698), .Z1_t (new_AGEMA_signal_18699), .Z1_f (new_AGEMA_signal_18700) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_71_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_71_MUX_inst_Y), .A0_f (new_AGEMA_signal_18698), .A1_t (new_AGEMA_signal_18699), .A1_f (new_AGEMA_signal_18700), .B0_t (RoundOutput[71]), .B0_f (new_AGEMA_signal_17534), .B1_t (new_AGEMA_signal_17535), .B1_f (new_AGEMA_signal_17536), .Z0_t (RoundInput[71]), .Z0_f (new_AGEMA_signal_5924), .Z1_t (new_AGEMA_signal_5925), .Z1_f (new_AGEMA_signal_5926) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_72_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[72]), .A0_f (new_AGEMA_signal_17537), .A1_t (new_AGEMA_signal_17538), .A1_f (new_AGEMA_signal_17539), .B0_t (plaintext_s0_t[72]), .B0_f (plaintext_s0_f[72]), .B1_t (plaintext_s1_t[72]), .B1_f (plaintext_s1_f[72]), .Z0_t (RoundReg_Inst_ff_SDE_72_MUX_inst_X), .Z0_f (new_AGEMA_signal_18176), .Z1_t (new_AGEMA_signal_18177), .Z1_f (new_AGEMA_signal_18178) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_72_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_72_MUX_inst_X), .B0_f (new_AGEMA_signal_18176), .B1_t (new_AGEMA_signal_18177), .B1_f (new_AGEMA_signal_18178), .Z0_t (RoundReg_Inst_ff_SDE_72_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18701), .Z1_t (new_AGEMA_signal_18702), .Z1_f (new_AGEMA_signal_18703) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_72_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_72_MUX_inst_Y), .A0_f (new_AGEMA_signal_18701), .A1_t (new_AGEMA_signal_18702), .A1_f (new_AGEMA_signal_18703), .B0_t (RoundOutput[72]), .B0_f (new_AGEMA_signal_17537), .B1_t (new_AGEMA_signal_17538), .B1_f (new_AGEMA_signal_17539), .Z0_t (RoundInput[72]), .Z0_f (new_AGEMA_signal_5933), .Z1_t (new_AGEMA_signal_5934), .Z1_f (new_AGEMA_signal_5935) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_73_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[73]), .A0_f (new_AGEMA_signal_17867), .A1_t (new_AGEMA_signal_17868), .A1_f (new_AGEMA_signal_17869), .B0_t (plaintext_s0_t[73]), .B0_f (plaintext_s0_f[73]), .B1_t (plaintext_s1_t[73]), .B1_f (plaintext_s1_f[73]), .Z0_t (RoundReg_Inst_ff_SDE_73_MUX_inst_X), .Z0_f (new_AGEMA_signal_18707), .Z1_t (new_AGEMA_signal_18708), .Z1_f (new_AGEMA_signal_18709) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_73_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_73_MUX_inst_X), .B0_f (new_AGEMA_signal_18707), .B1_t (new_AGEMA_signal_18708), .B1_f (new_AGEMA_signal_18709), .Z0_t (RoundReg_Inst_ff_SDE_73_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19013), .Z1_t (new_AGEMA_signal_19014), .Z1_f (new_AGEMA_signal_19015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_73_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_73_MUX_inst_Y), .A0_f (new_AGEMA_signal_19013), .A1_t (new_AGEMA_signal_19014), .A1_f (new_AGEMA_signal_19015), .B0_t (RoundOutput[73]), .B0_f (new_AGEMA_signal_17867), .B1_t (new_AGEMA_signal_17868), .B1_f (new_AGEMA_signal_17869), .Z0_t (RoundInput[73]), .Z0_f (new_AGEMA_signal_5942), .Z1_t (new_AGEMA_signal_5943), .Z1_f (new_AGEMA_signal_5944) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_74_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[74]), .A0_f (new_AGEMA_signal_17543), .A1_t (new_AGEMA_signal_17544), .A1_f (new_AGEMA_signal_17545), .B0_t (plaintext_s0_t[74]), .B0_f (plaintext_s0_f[74]), .B1_t (plaintext_s1_t[74]), .B1_f (plaintext_s1_f[74]), .Z0_t (RoundReg_Inst_ff_SDE_74_MUX_inst_X), .Z0_f (new_AGEMA_signal_18182), .Z1_t (new_AGEMA_signal_18183), .Z1_f (new_AGEMA_signal_18184) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_74_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_74_MUX_inst_X), .B0_f (new_AGEMA_signal_18182), .B1_t (new_AGEMA_signal_18183), .B1_f (new_AGEMA_signal_18184), .Z0_t (RoundReg_Inst_ff_SDE_74_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18710), .Z1_t (new_AGEMA_signal_18711), .Z1_f (new_AGEMA_signal_18712) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_74_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_74_MUX_inst_Y), .A0_f (new_AGEMA_signal_18710), .A1_t (new_AGEMA_signal_18711), .A1_f (new_AGEMA_signal_18712), .B0_t (RoundOutput[74]), .B0_f (new_AGEMA_signal_17543), .B1_t (new_AGEMA_signal_17544), .B1_f (new_AGEMA_signal_17545), .Z0_t (RoundInput[74]), .Z0_f (new_AGEMA_signal_5951), .Z1_t (new_AGEMA_signal_5952), .Z1_f (new_AGEMA_signal_5953) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_75_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[75]), .A0_f (new_AGEMA_signal_17870), .A1_t (new_AGEMA_signal_17871), .A1_f (new_AGEMA_signal_17872), .B0_t (plaintext_s0_t[75]), .B0_f (plaintext_s0_f[75]), .B1_t (plaintext_s1_t[75]), .B1_f (plaintext_s1_f[75]), .Z0_t (RoundReg_Inst_ff_SDE_75_MUX_inst_X), .Z0_f (new_AGEMA_signal_18716), .Z1_t (new_AGEMA_signal_18717), .Z1_f (new_AGEMA_signal_18718) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_75_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_75_MUX_inst_X), .B0_f (new_AGEMA_signal_18716), .B1_t (new_AGEMA_signal_18717), .B1_f (new_AGEMA_signal_18718), .Z0_t (RoundReg_Inst_ff_SDE_75_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19016), .Z1_t (new_AGEMA_signal_19017), .Z1_f (new_AGEMA_signal_19018) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_75_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_75_MUX_inst_Y), .A0_f (new_AGEMA_signal_19016), .A1_t (new_AGEMA_signal_19017), .A1_f (new_AGEMA_signal_19018), .B0_t (RoundOutput[75]), .B0_f (new_AGEMA_signal_17870), .B1_t (new_AGEMA_signal_17871), .B1_f (new_AGEMA_signal_17872), .Z0_t (RoundInput[75]), .Z0_f (new_AGEMA_signal_5960), .Z1_t (new_AGEMA_signal_5961), .Z1_f (new_AGEMA_signal_5962) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_76_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[76]), .A0_f (new_AGEMA_signal_17873), .A1_t (new_AGEMA_signal_17874), .A1_f (new_AGEMA_signal_17875), .B0_t (plaintext_s0_t[76]), .B0_f (plaintext_s0_f[76]), .B1_t (plaintext_s1_t[76]), .B1_f (plaintext_s1_f[76]), .Z0_t (RoundReg_Inst_ff_SDE_76_MUX_inst_X), .Z0_f (new_AGEMA_signal_18722), .Z1_t (new_AGEMA_signal_18723), .Z1_f (new_AGEMA_signal_18724) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_76_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_76_MUX_inst_X), .B0_f (new_AGEMA_signal_18722), .B1_t (new_AGEMA_signal_18723), .B1_f (new_AGEMA_signal_18724), .Z0_t (RoundReg_Inst_ff_SDE_76_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19019), .Z1_t (new_AGEMA_signal_19020), .Z1_f (new_AGEMA_signal_19021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_76_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_76_MUX_inst_Y), .A0_f (new_AGEMA_signal_19019), .A1_t (new_AGEMA_signal_19020), .A1_f (new_AGEMA_signal_19021), .B0_t (RoundOutput[76]), .B0_f (new_AGEMA_signal_17873), .B1_t (new_AGEMA_signal_17874), .B1_f (new_AGEMA_signal_17875), .Z0_t (RoundInput[76]), .Z0_f (new_AGEMA_signal_5969), .Z1_t (new_AGEMA_signal_5970), .Z1_f (new_AGEMA_signal_5971) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_77_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[77]), .A0_f (new_AGEMA_signal_17552), .A1_t (new_AGEMA_signal_17553), .A1_f (new_AGEMA_signal_17554), .B0_t (plaintext_s0_t[77]), .B0_f (plaintext_s0_f[77]), .B1_t (plaintext_s1_t[77]), .B1_f (plaintext_s1_f[77]), .Z0_t (RoundReg_Inst_ff_SDE_77_MUX_inst_X), .Z0_f (new_AGEMA_signal_18188), .Z1_t (new_AGEMA_signal_18189), .Z1_f (new_AGEMA_signal_18190) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_77_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_77_MUX_inst_X), .B0_f (new_AGEMA_signal_18188), .B1_t (new_AGEMA_signal_18189), .B1_f (new_AGEMA_signal_18190), .Z0_t (RoundReg_Inst_ff_SDE_77_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18725), .Z1_t (new_AGEMA_signal_18726), .Z1_f (new_AGEMA_signal_18727) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_77_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_77_MUX_inst_Y), .A0_f (new_AGEMA_signal_18725), .A1_t (new_AGEMA_signal_18726), .A1_f (new_AGEMA_signal_18727), .B0_t (RoundOutput[77]), .B0_f (new_AGEMA_signal_17552), .B1_t (new_AGEMA_signal_17553), .B1_f (new_AGEMA_signal_17554), .Z0_t (RoundInput[77]), .Z0_f (new_AGEMA_signal_5978), .Z1_t (new_AGEMA_signal_5979), .Z1_f (new_AGEMA_signal_5980) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_78_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[78]), .A0_f (new_AGEMA_signal_17555), .A1_t (new_AGEMA_signal_17556), .A1_f (new_AGEMA_signal_17557), .B0_t (plaintext_s0_t[78]), .B0_f (plaintext_s0_f[78]), .B1_t (plaintext_s1_t[78]), .B1_f (plaintext_s1_f[78]), .Z0_t (RoundReg_Inst_ff_SDE_78_MUX_inst_X), .Z0_f (new_AGEMA_signal_18194), .Z1_t (new_AGEMA_signal_18195), .Z1_f (new_AGEMA_signal_18196) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_78_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_78_MUX_inst_X), .B0_f (new_AGEMA_signal_18194), .B1_t (new_AGEMA_signal_18195), .B1_f (new_AGEMA_signal_18196), .Z0_t (RoundReg_Inst_ff_SDE_78_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18728), .Z1_t (new_AGEMA_signal_18729), .Z1_f (new_AGEMA_signal_18730) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_78_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_78_MUX_inst_Y), .A0_f (new_AGEMA_signal_18728), .A1_t (new_AGEMA_signal_18729), .A1_f (new_AGEMA_signal_18730), .B0_t (RoundOutput[78]), .B0_f (new_AGEMA_signal_17555), .B1_t (new_AGEMA_signal_17556), .B1_f (new_AGEMA_signal_17557), .Z0_t (RoundInput[78]), .Z0_f (new_AGEMA_signal_5987), .Z1_t (new_AGEMA_signal_5988), .Z1_f (new_AGEMA_signal_5989) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_79_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[79]), .A0_f (new_AGEMA_signal_17558), .A1_t (new_AGEMA_signal_17559), .A1_f (new_AGEMA_signal_17560), .B0_t (plaintext_s0_t[79]), .B0_f (plaintext_s0_f[79]), .B1_t (plaintext_s1_t[79]), .B1_f (plaintext_s1_f[79]), .Z0_t (RoundReg_Inst_ff_SDE_79_MUX_inst_X), .Z0_f (new_AGEMA_signal_18200), .Z1_t (new_AGEMA_signal_18201), .Z1_f (new_AGEMA_signal_18202) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_79_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_79_MUX_inst_X), .B0_f (new_AGEMA_signal_18200), .B1_t (new_AGEMA_signal_18201), .B1_f (new_AGEMA_signal_18202), .Z0_t (RoundReg_Inst_ff_SDE_79_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18731), .Z1_t (new_AGEMA_signal_18732), .Z1_f (new_AGEMA_signal_18733) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_79_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_79_MUX_inst_Y), .A0_f (new_AGEMA_signal_18731), .A1_t (new_AGEMA_signal_18732), .A1_f (new_AGEMA_signal_18733), .B0_t (RoundOutput[79]), .B0_f (new_AGEMA_signal_17558), .B1_t (new_AGEMA_signal_17559), .B1_f (new_AGEMA_signal_17560), .Z0_t (RoundInput[79]), .Z0_f (new_AGEMA_signal_5996), .Z1_t (new_AGEMA_signal_5997), .Z1_f (new_AGEMA_signal_5998) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_80_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[80]), .A0_f (new_AGEMA_signal_17564), .A1_t (new_AGEMA_signal_17565), .A1_f (new_AGEMA_signal_17566), .B0_t (plaintext_s0_t[80]), .B0_f (plaintext_s0_f[80]), .B1_t (plaintext_s1_t[80]), .B1_f (plaintext_s1_f[80]), .Z0_t (RoundReg_Inst_ff_SDE_80_MUX_inst_X), .Z0_f (new_AGEMA_signal_18206), .Z1_t (new_AGEMA_signal_18207), .Z1_f (new_AGEMA_signal_18208) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_80_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_80_MUX_inst_X), .B0_f (new_AGEMA_signal_18206), .B1_t (new_AGEMA_signal_18207), .B1_f (new_AGEMA_signal_18208), .Z0_t (RoundReg_Inst_ff_SDE_80_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18734), .Z1_t (new_AGEMA_signal_18735), .Z1_f (new_AGEMA_signal_18736) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_80_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_80_MUX_inst_Y), .A0_f (new_AGEMA_signal_18734), .A1_t (new_AGEMA_signal_18735), .A1_f (new_AGEMA_signal_18736), .B0_t (RoundOutput[80]), .B0_f (new_AGEMA_signal_17564), .B1_t (new_AGEMA_signal_17565), .B1_f (new_AGEMA_signal_17566), .Z0_t (RoundInput[80]), .Z0_f (new_AGEMA_signal_6014), .Z1_t (new_AGEMA_signal_6015), .Z1_f (new_AGEMA_signal_6016) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_81_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[81]), .A0_f (new_AGEMA_signal_17876), .A1_t (new_AGEMA_signal_17877), .A1_f (new_AGEMA_signal_17878), .B0_t (plaintext_s0_t[81]), .B0_f (plaintext_s0_f[81]), .B1_t (plaintext_s1_t[81]), .B1_f (plaintext_s1_f[81]), .Z0_t (RoundReg_Inst_ff_SDE_81_MUX_inst_X), .Z0_f (new_AGEMA_signal_18740), .Z1_t (new_AGEMA_signal_18741), .Z1_f (new_AGEMA_signal_18742) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_81_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_81_MUX_inst_X), .B0_f (new_AGEMA_signal_18740), .B1_t (new_AGEMA_signal_18741), .B1_f (new_AGEMA_signal_18742), .Z0_t (RoundReg_Inst_ff_SDE_81_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19022), .Z1_t (new_AGEMA_signal_19023), .Z1_f (new_AGEMA_signal_19024) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_81_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_81_MUX_inst_Y), .A0_f (new_AGEMA_signal_19022), .A1_t (new_AGEMA_signal_19023), .A1_f (new_AGEMA_signal_19024), .B0_t (RoundOutput[81]), .B0_f (new_AGEMA_signal_17876), .B1_t (new_AGEMA_signal_17877), .B1_f (new_AGEMA_signal_17878), .Z0_t (RoundInput[81]), .Z0_f (new_AGEMA_signal_6023), .Z1_t (new_AGEMA_signal_6024), .Z1_f (new_AGEMA_signal_6025) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_82_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[82]), .A0_f (new_AGEMA_signal_17570), .A1_t (new_AGEMA_signal_17571), .A1_f (new_AGEMA_signal_17572), .B0_t (plaintext_s0_t[82]), .B0_f (plaintext_s0_f[82]), .B1_t (plaintext_s1_t[82]), .B1_f (plaintext_s1_f[82]), .Z0_t (RoundReg_Inst_ff_SDE_82_MUX_inst_X), .Z0_f (new_AGEMA_signal_18212), .Z1_t (new_AGEMA_signal_18213), .Z1_f (new_AGEMA_signal_18214) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_82_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_82_MUX_inst_X), .B0_f (new_AGEMA_signal_18212), .B1_t (new_AGEMA_signal_18213), .B1_f (new_AGEMA_signal_18214), .Z0_t (RoundReg_Inst_ff_SDE_82_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18743), .Z1_t (new_AGEMA_signal_18744), .Z1_f (new_AGEMA_signal_18745) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_82_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_82_MUX_inst_Y), .A0_f (new_AGEMA_signal_18743), .A1_t (new_AGEMA_signal_18744), .A1_f (new_AGEMA_signal_18745), .B0_t (RoundOutput[82]), .B0_f (new_AGEMA_signal_17570), .B1_t (new_AGEMA_signal_17571), .B1_f (new_AGEMA_signal_17572), .Z0_t (RoundInput[82]), .Z0_f (new_AGEMA_signal_6032), .Z1_t (new_AGEMA_signal_6033), .Z1_f (new_AGEMA_signal_6034) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_83_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[83]), .A0_f (new_AGEMA_signal_17879), .A1_t (new_AGEMA_signal_17880), .A1_f (new_AGEMA_signal_17881), .B0_t (plaintext_s0_t[83]), .B0_f (plaintext_s0_f[83]), .B1_t (plaintext_s1_t[83]), .B1_f (plaintext_s1_f[83]), .Z0_t (RoundReg_Inst_ff_SDE_83_MUX_inst_X), .Z0_f (new_AGEMA_signal_18749), .Z1_t (new_AGEMA_signal_18750), .Z1_f (new_AGEMA_signal_18751) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_83_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_83_MUX_inst_X), .B0_f (new_AGEMA_signal_18749), .B1_t (new_AGEMA_signal_18750), .B1_f (new_AGEMA_signal_18751), .Z0_t (RoundReg_Inst_ff_SDE_83_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19025), .Z1_t (new_AGEMA_signal_19026), .Z1_f (new_AGEMA_signal_19027) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_83_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_83_MUX_inst_Y), .A0_f (new_AGEMA_signal_19025), .A1_t (new_AGEMA_signal_19026), .A1_f (new_AGEMA_signal_19027), .B0_t (RoundOutput[83]), .B0_f (new_AGEMA_signal_17879), .B1_t (new_AGEMA_signal_17880), .B1_f (new_AGEMA_signal_17881), .Z0_t (RoundInput[83]), .Z0_f (new_AGEMA_signal_6041), .Z1_t (new_AGEMA_signal_6042), .Z1_f (new_AGEMA_signal_6043) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_84_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[84]), .A0_f (new_AGEMA_signal_17882), .A1_t (new_AGEMA_signal_17883), .A1_f (new_AGEMA_signal_17884), .B0_t (plaintext_s0_t[84]), .B0_f (plaintext_s0_f[84]), .B1_t (plaintext_s1_t[84]), .B1_f (plaintext_s1_f[84]), .Z0_t (RoundReg_Inst_ff_SDE_84_MUX_inst_X), .Z0_f (new_AGEMA_signal_18755), .Z1_t (new_AGEMA_signal_18756), .Z1_f (new_AGEMA_signal_18757) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_84_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_84_MUX_inst_X), .B0_f (new_AGEMA_signal_18755), .B1_t (new_AGEMA_signal_18756), .B1_f (new_AGEMA_signal_18757), .Z0_t (RoundReg_Inst_ff_SDE_84_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19028), .Z1_t (new_AGEMA_signal_19029), .Z1_f (new_AGEMA_signal_19030) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_84_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_84_MUX_inst_Y), .A0_f (new_AGEMA_signal_19028), .A1_t (new_AGEMA_signal_19029), .A1_f (new_AGEMA_signal_19030), .B0_t (RoundOutput[84]), .B0_f (new_AGEMA_signal_17882), .B1_t (new_AGEMA_signal_17883), .B1_f (new_AGEMA_signal_17884), .Z0_t (RoundInput[84]), .Z0_f (new_AGEMA_signal_6050), .Z1_t (new_AGEMA_signal_6051), .Z1_f (new_AGEMA_signal_6052) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_85_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[85]), .A0_f (new_AGEMA_signal_17579), .A1_t (new_AGEMA_signal_17580), .A1_f (new_AGEMA_signal_17581), .B0_t (plaintext_s0_t[85]), .B0_f (plaintext_s0_f[85]), .B1_t (plaintext_s1_t[85]), .B1_f (plaintext_s1_f[85]), .Z0_t (RoundReg_Inst_ff_SDE_85_MUX_inst_X), .Z0_f (new_AGEMA_signal_18218), .Z1_t (new_AGEMA_signal_18219), .Z1_f (new_AGEMA_signal_18220) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_85_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_85_MUX_inst_X), .B0_f (new_AGEMA_signal_18218), .B1_t (new_AGEMA_signal_18219), .B1_f (new_AGEMA_signal_18220), .Z0_t (RoundReg_Inst_ff_SDE_85_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18758), .Z1_t (new_AGEMA_signal_18759), .Z1_f (new_AGEMA_signal_18760) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_85_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_85_MUX_inst_Y), .A0_f (new_AGEMA_signal_18758), .A1_t (new_AGEMA_signal_18759), .A1_f (new_AGEMA_signal_18760), .B0_t (RoundOutput[85]), .B0_f (new_AGEMA_signal_17579), .B1_t (new_AGEMA_signal_17580), .B1_f (new_AGEMA_signal_17581), .Z0_t (RoundInput[85]), .Z0_f (new_AGEMA_signal_6059), .Z1_t (new_AGEMA_signal_6060), .Z1_f (new_AGEMA_signal_6061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_86_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[86]), .A0_f (new_AGEMA_signal_17582), .A1_t (new_AGEMA_signal_17583), .A1_f (new_AGEMA_signal_17584), .B0_t (plaintext_s0_t[86]), .B0_f (plaintext_s0_f[86]), .B1_t (plaintext_s1_t[86]), .B1_f (plaintext_s1_f[86]), .Z0_t (RoundReg_Inst_ff_SDE_86_MUX_inst_X), .Z0_f (new_AGEMA_signal_18224), .Z1_t (new_AGEMA_signal_18225), .Z1_f (new_AGEMA_signal_18226) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_86_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_86_MUX_inst_X), .B0_f (new_AGEMA_signal_18224), .B1_t (new_AGEMA_signal_18225), .B1_f (new_AGEMA_signal_18226), .Z0_t (RoundReg_Inst_ff_SDE_86_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18761), .Z1_t (new_AGEMA_signal_18762), .Z1_f (new_AGEMA_signal_18763) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_86_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_86_MUX_inst_Y), .A0_f (new_AGEMA_signal_18761), .A1_t (new_AGEMA_signal_18762), .A1_f (new_AGEMA_signal_18763), .B0_t (RoundOutput[86]), .B0_f (new_AGEMA_signal_17582), .B1_t (new_AGEMA_signal_17583), .B1_f (new_AGEMA_signal_17584), .Z0_t (RoundInput[86]), .Z0_f (new_AGEMA_signal_6068), .Z1_t (new_AGEMA_signal_6069), .Z1_f (new_AGEMA_signal_6070) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_87_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[87]), .A0_f (new_AGEMA_signal_17585), .A1_t (new_AGEMA_signal_17586), .A1_f (new_AGEMA_signal_17587), .B0_t (plaintext_s0_t[87]), .B0_f (plaintext_s0_f[87]), .B1_t (plaintext_s1_t[87]), .B1_f (plaintext_s1_f[87]), .Z0_t (RoundReg_Inst_ff_SDE_87_MUX_inst_X), .Z0_f (new_AGEMA_signal_18230), .Z1_t (new_AGEMA_signal_18231), .Z1_f (new_AGEMA_signal_18232) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_87_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_87_MUX_inst_X), .B0_f (new_AGEMA_signal_18230), .B1_t (new_AGEMA_signal_18231), .B1_f (new_AGEMA_signal_18232), .Z0_t (RoundReg_Inst_ff_SDE_87_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18764), .Z1_t (new_AGEMA_signal_18765), .Z1_f (new_AGEMA_signal_18766) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_87_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_87_MUX_inst_Y), .A0_f (new_AGEMA_signal_18764), .A1_t (new_AGEMA_signal_18765), .A1_f (new_AGEMA_signal_18766), .B0_t (RoundOutput[87]), .B0_f (new_AGEMA_signal_17585), .B1_t (new_AGEMA_signal_17586), .B1_f (new_AGEMA_signal_17587), .Z0_t (RoundInput[87]), .Z0_f (new_AGEMA_signal_6077), .Z1_t (new_AGEMA_signal_6078), .Z1_f (new_AGEMA_signal_6079) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_88_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[88]), .A0_f (new_AGEMA_signal_17588), .A1_t (new_AGEMA_signal_17589), .A1_f (new_AGEMA_signal_17590), .B0_t (plaintext_s0_t[88]), .B0_f (plaintext_s0_f[88]), .B1_t (plaintext_s1_t[88]), .B1_f (plaintext_s1_f[88]), .Z0_t (RoundReg_Inst_ff_SDE_88_MUX_inst_X), .Z0_f (new_AGEMA_signal_18236), .Z1_t (new_AGEMA_signal_18237), .Z1_f (new_AGEMA_signal_18238) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_88_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_88_MUX_inst_X), .B0_f (new_AGEMA_signal_18236), .B1_t (new_AGEMA_signal_18237), .B1_f (new_AGEMA_signal_18238), .Z0_t (RoundReg_Inst_ff_SDE_88_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18767), .Z1_t (new_AGEMA_signal_18768), .Z1_f (new_AGEMA_signal_18769) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_88_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_88_MUX_inst_Y), .A0_f (new_AGEMA_signal_18767), .A1_t (new_AGEMA_signal_18768), .A1_f (new_AGEMA_signal_18769), .B0_t (RoundOutput[88]), .B0_f (new_AGEMA_signal_17588), .B1_t (new_AGEMA_signal_17589), .B1_f (new_AGEMA_signal_17590), .Z0_t (RoundInput[88]), .Z0_f (new_AGEMA_signal_6086), .Z1_t (new_AGEMA_signal_6087), .Z1_f (new_AGEMA_signal_6088) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_89_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[89]), .A0_f (new_AGEMA_signal_17885), .A1_t (new_AGEMA_signal_17886), .A1_f (new_AGEMA_signal_17887), .B0_t (plaintext_s0_t[89]), .B0_f (plaintext_s0_f[89]), .B1_t (plaintext_s1_t[89]), .B1_f (plaintext_s1_f[89]), .Z0_t (RoundReg_Inst_ff_SDE_89_MUX_inst_X), .Z0_f (new_AGEMA_signal_18773), .Z1_t (new_AGEMA_signal_18774), .Z1_f (new_AGEMA_signal_18775) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_89_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_89_MUX_inst_X), .B0_f (new_AGEMA_signal_18773), .B1_t (new_AGEMA_signal_18774), .B1_f (new_AGEMA_signal_18775), .Z0_t (RoundReg_Inst_ff_SDE_89_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19031), .Z1_t (new_AGEMA_signal_19032), .Z1_f (new_AGEMA_signal_19033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_89_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_89_MUX_inst_Y), .A0_f (new_AGEMA_signal_19031), .A1_t (new_AGEMA_signal_19032), .A1_f (new_AGEMA_signal_19033), .B0_t (RoundOutput[89]), .B0_f (new_AGEMA_signal_17885), .B1_t (new_AGEMA_signal_17886), .B1_f (new_AGEMA_signal_17887), .Z0_t (RoundInput[89]), .Z0_f (new_AGEMA_signal_6095), .Z1_t (new_AGEMA_signal_6096), .Z1_f (new_AGEMA_signal_6097) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_90_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[90]), .A0_f (new_AGEMA_signal_17597), .A1_t (new_AGEMA_signal_17598), .A1_f (new_AGEMA_signal_17599), .B0_t (plaintext_s0_t[90]), .B0_f (plaintext_s0_f[90]), .B1_t (plaintext_s1_t[90]), .B1_f (plaintext_s1_f[90]), .Z0_t (RoundReg_Inst_ff_SDE_90_MUX_inst_X), .Z0_f (new_AGEMA_signal_18242), .Z1_t (new_AGEMA_signal_18243), .Z1_f (new_AGEMA_signal_18244) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_90_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_90_MUX_inst_X), .B0_f (new_AGEMA_signal_18242), .B1_t (new_AGEMA_signal_18243), .B1_f (new_AGEMA_signal_18244), .Z0_t (RoundReg_Inst_ff_SDE_90_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18776), .Z1_t (new_AGEMA_signal_18777), .Z1_f (new_AGEMA_signal_18778) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_90_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_90_MUX_inst_Y), .A0_f (new_AGEMA_signal_18776), .A1_t (new_AGEMA_signal_18777), .A1_f (new_AGEMA_signal_18778), .B0_t (RoundOutput[90]), .B0_f (new_AGEMA_signal_17597), .B1_t (new_AGEMA_signal_17598), .B1_f (new_AGEMA_signal_17599), .Z0_t (RoundInput[90]), .Z0_f (new_AGEMA_signal_6113), .Z1_t (new_AGEMA_signal_6114), .Z1_f (new_AGEMA_signal_6115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_91_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[91]), .A0_f (new_AGEMA_signal_17888), .A1_t (new_AGEMA_signal_17889), .A1_f (new_AGEMA_signal_17890), .B0_t (plaintext_s0_t[91]), .B0_f (plaintext_s0_f[91]), .B1_t (plaintext_s1_t[91]), .B1_f (plaintext_s1_f[91]), .Z0_t (RoundReg_Inst_ff_SDE_91_MUX_inst_X), .Z0_f (new_AGEMA_signal_18782), .Z1_t (new_AGEMA_signal_18783), .Z1_f (new_AGEMA_signal_18784) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_91_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_91_MUX_inst_X), .B0_f (new_AGEMA_signal_18782), .B1_t (new_AGEMA_signal_18783), .B1_f (new_AGEMA_signal_18784), .Z0_t (RoundReg_Inst_ff_SDE_91_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19034), .Z1_t (new_AGEMA_signal_19035), .Z1_f (new_AGEMA_signal_19036) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_91_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_91_MUX_inst_Y), .A0_f (new_AGEMA_signal_19034), .A1_t (new_AGEMA_signal_19035), .A1_f (new_AGEMA_signal_19036), .B0_t (RoundOutput[91]), .B0_f (new_AGEMA_signal_17888), .B1_t (new_AGEMA_signal_17889), .B1_f (new_AGEMA_signal_17890), .Z0_t (RoundInput[91]), .Z0_f (new_AGEMA_signal_6122), .Z1_t (new_AGEMA_signal_6123), .Z1_f (new_AGEMA_signal_6124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_92_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[92]), .A0_f (new_AGEMA_signal_17891), .A1_t (new_AGEMA_signal_17892), .A1_f (new_AGEMA_signal_17893), .B0_t (plaintext_s0_t[92]), .B0_f (plaintext_s0_f[92]), .B1_t (plaintext_s1_t[92]), .B1_f (plaintext_s1_f[92]), .Z0_t (RoundReg_Inst_ff_SDE_92_MUX_inst_X), .Z0_f (new_AGEMA_signal_18788), .Z1_t (new_AGEMA_signal_18789), .Z1_f (new_AGEMA_signal_18790) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_92_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_92_MUX_inst_X), .B0_f (new_AGEMA_signal_18788), .B1_t (new_AGEMA_signal_18789), .B1_f (new_AGEMA_signal_18790), .Z0_t (RoundReg_Inst_ff_SDE_92_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19037), .Z1_t (new_AGEMA_signal_19038), .Z1_f (new_AGEMA_signal_19039) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_92_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_92_MUX_inst_Y), .A0_f (new_AGEMA_signal_19037), .A1_t (new_AGEMA_signal_19038), .A1_f (new_AGEMA_signal_19039), .B0_t (RoundOutput[92]), .B0_f (new_AGEMA_signal_17891), .B1_t (new_AGEMA_signal_17892), .B1_f (new_AGEMA_signal_17893), .Z0_t (RoundInput[92]), .Z0_f (new_AGEMA_signal_6131), .Z1_t (new_AGEMA_signal_6132), .Z1_f (new_AGEMA_signal_6133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_93_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[93]), .A0_f (new_AGEMA_signal_17606), .A1_t (new_AGEMA_signal_17607), .A1_f (new_AGEMA_signal_17608), .B0_t (plaintext_s0_t[93]), .B0_f (plaintext_s0_f[93]), .B1_t (plaintext_s1_t[93]), .B1_f (plaintext_s1_f[93]), .Z0_t (RoundReg_Inst_ff_SDE_93_MUX_inst_X), .Z0_f (new_AGEMA_signal_18248), .Z1_t (new_AGEMA_signal_18249), .Z1_f (new_AGEMA_signal_18250) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_93_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_93_MUX_inst_X), .B0_f (new_AGEMA_signal_18248), .B1_t (new_AGEMA_signal_18249), .B1_f (new_AGEMA_signal_18250), .Z0_t (RoundReg_Inst_ff_SDE_93_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18791), .Z1_t (new_AGEMA_signal_18792), .Z1_f (new_AGEMA_signal_18793) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_93_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_93_MUX_inst_Y), .A0_f (new_AGEMA_signal_18791), .A1_t (new_AGEMA_signal_18792), .A1_f (new_AGEMA_signal_18793), .B0_t (RoundOutput[93]), .B0_f (new_AGEMA_signal_17606), .B1_t (new_AGEMA_signal_17607), .B1_f (new_AGEMA_signal_17608), .Z0_t (RoundInput[93]), .Z0_f (new_AGEMA_signal_6140), .Z1_t (new_AGEMA_signal_6141), .Z1_f (new_AGEMA_signal_6142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_94_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[94]), .A0_f (new_AGEMA_signal_17609), .A1_t (new_AGEMA_signal_17610), .A1_f (new_AGEMA_signal_17611), .B0_t (plaintext_s0_t[94]), .B0_f (plaintext_s0_f[94]), .B1_t (plaintext_s1_t[94]), .B1_f (plaintext_s1_f[94]), .Z0_t (RoundReg_Inst_ff_SDE_94_MUX_inst_X), .Z0_f (new_AGEMA_signal_18254), .Z1_t (new_AGEMA_signal_18255), .Z1_f (new_AGEMA_signal_18256) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_94_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_94_MUX_inst_X), .B0_f (new_AGEMA_signal_18254), .B1_t (new_AGEMA_signal_18255), .B1_f (new_AGEMA_signal_18256), .Z0_t (RoundReg_Inst_ff_SDE_94_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18794), .Z1_t (new_AGEMA_signal_18795), .Z1_f (new_AGEMA_signal_18796) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_94_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_94_MUX_inst_Y), .A0_f (new_AGEMA_signal_18794), .A1_t (new_AGEMA_signal_18795), .A1_f (new_AGEMA_signal_18796), .B0_t (RoundOutput[94]), .B0_f (new_AGEMA_signal_17609), .B1_t (new_AGEMA_signal_17610), .B1_f (new_AGEMA_signal_17611), .Z0_t (RoundInput[94]), .Z0_f (new_AGEMA_signal_6149), .Z1_t (new_AGEMA_signal_6150), .Z1_f (new_AGEMA_signal_6151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_95_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[95]), .A0_f (new_AGEMA_signal_17612), .A1_t (new_AGEMA_signal_17613), .A1_f (new_AGEMA_signal_17614), .B0_t (plaintext_s0_t[95]), .B0_f (plaintext_s0_f[95]), .B1_t (plaintext_s1_t[95]), .B1_f (plaintext_s1_f[95]), .Z0_t (RoundReg_Inst_ff_SDE_95_MUX_inst_X), .Z0_f (new_AGEMA_signal_18260), .Z1_t (new_AGEMA_signal_18261), .Z1_f (new_AGEMA_signal_18262) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_95_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_95_MUX_inst_X), .B0_f (new_AGEMA_signal_18260), .B1_t (new_AGEMA_signal_18261), .B1_f (new_AGEMA_signal_18262), .Z0_t (RoundReg_Inst_ff_SDE_95_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18797), .Z1_t (new_AGEMA_signal_18798), .Z1_f (new_AGEMA_signal_18799) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_95_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_95_MUX_inst_Y), .A0_f (new_AGEMA_signal_18797), .A1_t (new_AGEMA_signal_18798), .A1_f (new_AGEMA_signal_18799), .B0_t (RoundOutput[95]), .B0_f (new_AGEMA_signal_17612), .B1_t (new_AGEMA_signal_17613), .B1_f (new_AGEMA_signal_17614), .Z0_t (RoundInput[95]), .Z0_f (new_AGEMA_signal_6158), .Z1_t (new_AGEMA_signal_6159), .Z1_f (new_AGEMA_signal_6160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_96_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[96]), .A0_f (new_AGEMA_signal_17615), .A1_t (new_AGEMA_signal_17616), .A1_f (new_AGEMA_signal_17617), .B0_t (plaintext_s0_t[96]), .B0_f (plaintext_s0_f[96]), .B1_t (plaintext_s1_t[96]), .B1_f (plaintext_s1_f[96]), .Z0_t (RoundReg_Inst_ff_SDE_96_MUX_inst_X), .Z0_f (new_AGEMA_signal_18266), .Z1_t (new_AGEMA_signal_18267), .Z1_f (new_AGEMA_signal_18268) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_96_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_96_MUX_inst_X), .B0_f (new_AGEMA_signal_18266), .B1_t (new_AGEMA_signal_18267), .B1_f (new_AGEMA_signal_18268), .Z0_t (RoundReg_Inst_ff_SDE_96_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18800), .Z1_t (new_AGEMA_signal_18801), .Z1_f (new_AGEMA_signal_18802) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_96_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_96_MUX_inst_Y), .A0_f (new_AGEMA_signal_18800), .A1_t (new_AGEMA_signal_18801), .A1_f (new_AGEMA_signal_18802), .B0_t (RoundOutput[96]), .B0_f (new_AGEMA_signal_17615), .B1_t (new_AGEMA_signal_17616), .B1_f (new_AGEMA_signal_17617), .Z0_t (RoundInput[96]), .Z0_f (new_AGEMA_signal_6167), .Z1_t (new_AGEMA_signal_6168), .Z1_f (new_AGEMA_signal_6169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_97_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[97]), .A0_f (new_AGEMA_signal_17894), .A1_t (new_AGEMA_signal_17895), .A1_f (new_AGEMA_signal_17896), .B0_t (plaintext_s0_t[97]), .B0_f (plaintext_s0_f[97]), .B1_t (plaintext_s1_t[97]), .B1_f (plaintext_s1_f[97]), .Z0_t (RoundReg_Inst_ff_SDE_97_MUX_inst_X), .Z0_f (new_AGEMA_signal_18806), .Z1_t (new_AGEMA_signal_18807), .Z1_f (new_AGEMA_signal_18808) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_97_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_97_MUX_inst_X), .B0_f (new_AGEMA_signal_18806), .B1_t (new_AGEMA_signal_18807), .B1_f (new_AGEMA_signal_18808), .Z0_t (RoundReg_Inst_ff_SDE_97_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19040), .Z1_t (new_AGEMA_signal_19041), .Z1_f (new_AGEMA_signal_19042) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_97_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_97_MUX_inst_Y), .A0_f (new_AGEMA_signal_19040), .A1_t (new_AGEMA_signal_19041), .A1_f (new_AGEMA_signal_19042), .B0_t (RoundOutput[97]), .B0_f (new_AGEMA_signal_17894), .B1_t (new_AGEMA_signal_17895), .B1_f (new_AGEMA_signal_17896), .Z0_t (RoundInput[97]), .Z0_f (new_AGEMA_signal_6176), .Z1_t (new_AGEMA_signal_6177), .Z1_f (new_AGEMA_signal_6178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_98_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[98]), .A0_f (new_AGEMA_signal_17621), .A1_t (new_AGEMA_signal_17622), .A1_f (new_AGEMA_signal_17623), .B0_t (plaintext_s0_t[98]), .B0_f (plaintext_s0_f[98]), .B1_t (plaintext_s1_t[98]), .B1_f (plaintext_s1_f[98]), .Z0_t (RoundReg_Inst_ff_SDE_98_MUX_inst_X), .Z0_f (new_AGEMA_signal_18272), .Z1_t (new_AGEMA_signal_18273), .Z1_f (new_AGEMA_signal_18274) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_98_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_98_MUX_inst_X), .B0_f (new_AGEMA_signal_18272), .B1_t (new_AGEMA_signal_18273), .B1_f (new_AGEMA_signal_18274), .Z0_t (RoundReg_Inst_ff_SDE_98_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18809), .Z1_t (new_AGEMA_signal_18810), .Z1_f (new_AGEMA_signal_18811) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_98_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_98_MUX_inst_Y), .A0_f (new_AGEMA_signal_18809), .A1_t (new_AGEMA_signal_18810), .A1_f (new_AGEMA_signal_18811), .B0_t (RoundOutput[98]), .B0_f (new_AGEMA_signal_17621), .B1_t (new_AGEMA_signal_17622), .B1_f (new_AGEMA_signal_17623), .Z0_t (RoundInput[98]), .Z0_f (new_AGEMA_signal_6185), .Z1_t (new_AGEMA_signal_6186), .Z1_f (new_AGEMA_signal_6187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_99_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[99]), .A0_f (new_AGEMA_signal_17897), .A1_t (new_AGEMA_signal_17898), .A1_f (new_AGEMA_signal_17899), .B0_t (plaintext_s0_t[99]), .B0_f (plaintext_s0_f[99]), .B1_t (plaintext_s1_t[99]), .B1_f (plaintext_s1_f[99]), .Z0_t (RoundReg_Inst_ff_SDE_99_MUX_inst_X), .Z0_f (new_AGEMA_signal_18815), .Z1_t (new_AGEMA_signal_18816), .Z1_f (new_AGEMA_signal_18817) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_99_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_99_MUX_inst_X), .B0_f (new_AGEMA_signal_18815), .B1_t (new_AGEMA_signal_18816), .B1_f (new_AGEMA_signal_18817), .Z0_t (RoundReg_Inst_ff_SDE_99_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19043), .Z1_t (new_AGEMA_signal_19044), .Z1_f (new_AGEMA_signal_19045) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_99_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_99_MUX_inst_Y), .A0_f (new_AGEMA_signal_19043), .A1_t (new_AGEMA_signal_19044), .A1_f (new_AGEMA_signal_19045), .B0_t (RoundOutput[99]), .B0_f (new_AGEMA_signal_17897), .B1_t (new_AGEMA_signal_17898), .B1_f (new_AGEMA_signal_17899), .Z0_t (RoundInput[99]), .Z0_f (new_AGEMA_signal_6194), .Z1_t (new_AGEMA_signal_6195), .Z1_f (new_AGEMA_signal_6196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_100_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[100]), .A0_f (new_AGEMA_signal_17759), .A1_t (new_AGEMA_signal_17760), .A1_f (new_AGEMA_signal_17761), .B0_t (plaintext_s0_t[100]), .B0_f (plaintext_s0_f[100]), .B1_t (plaintext_s1_t[100]), .B1_f (plaintext_s1_f[100]), .Z0_t (RoundReg_Inst_ff_SDE_100_MUX_inst_X), .Z0_f (new_AGEMA_signal_18821), .Z1_t (new_AGEMA_signal_18822), .Z1_f (new_AGEMA_signal_18823) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_100_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_100_MUX_inst_X), .B0_f (new_AGEMA_signal_18821), .B1_t (new_AGEMA_signal_18822), .B1_f (new_AGEMA_signal_18823), .Z0_t (RoundReg_Inst_ff_SDE_100_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19046), .Z1_t (new_AGEMA_signal_19047), .Z1_f (new_AGEMA_signal_19048) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_100_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_100_MUX_inst_Y), .A0_f (new_AGEMA_signal_19046), .A1_t (new_AGEMA_signal_19047), .A1_f (new_AGEMA_signal_19048), .B0_t (RoundOutput[100]), .B0_f (new_AGEMA_signal_17759), .B1_t (new_AGEMA_signal_17760), .B1_f (new_AGEMA_signal_17761), .Z0_t (RoundInput[100]), .Z0_f (new_AGEMA_signal_5069), .Z1_t (new_AGEMA_signal_5070), .Z1_f (new_AGEMA_signal_5071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_101_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[101]), .A0_f (new_AGEMA_signal_17252), .A1_t (new_AGEMA_signal_17253), .A1_f (new_AGEMA_signal_17254), .B0_t (plaintext_s0_t[101]), .B0_f (plaintext_s0_f[101]), .B1_t (plaintext_s1_t[101]), .B1_f (plaintext_s1_f[101]), .Z0_t (RoundReg_Inst_ff_SDE_101_MUX_inst_X), .Z0_f (new_AGEMA_signal_18278), .Z1_t (new_AGEMA_signal_18279), .Z1_f (new_AGEMA_signal_18280) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_101_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_101_MUX_inst_X), .B0_f (new_AGEMA_signal_18278), .B1_t (new_AGEMA_signal_18279), .B1_f (new_AGEMA_signal_18280), .Z0_t (RoundReg_Inst_ff_SDE_101_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18824), .Z1_t (new_AGEMA_signal_18825), .Z1_f (new_AGEMA_signal_18826) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_101_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_101_MUX_inst_Y), .A0_f (new_AGEMA_signal_18824), .A1_t (new_AGEMA_signal_18825), .A1_f (new_AGEMA_signal_18826), .B0_t (RoundOutput[101]), .B0_f (new_AGEMA_signal_17252), .B1_t (new_AGEMA_signal_17253), .B1_f (new_AGEMA_signal_17254), .Z0_t (RoundInput[101]), .Z0_f (new_AGEMA_signal_5078), .Z1_t (new_AGEMA_signal_5079), .Z1_f (new_AGEMA_signal_5080) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_102_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[102]), .A0_f (new_AGEMA_signal_17255), .A1_t (new_AGEMA_signal_17256), .A1_f (new_AGEMA_signal_17257), .B0_t (plaintext_s0_t[102]), .B0_f (plaintext_s0_f[102]), .B1_t (plaintext_s1_t[102]), .B1_f (plaintext_s1_f[102]), .Z0_t (RoundReg_Inst_ff_SDE_102_MUX_inst_X), .Z0_f (new_AGEMA_signal_18284), .Z1_t (new_AGEMA_signal_18285), .Z1_f (new_AGEMA_signal_18286) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_102_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_102_MUX_inst_X), .B0_f (new_AGEMA_signal_18284), .B1_t (new_AGEMA_signal_18285), .B1_f (new_AGEMA_signal_18286), .Z0_t (RoundReg_Inst_ff_SDE_102_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18827), .Z1_t (new_AGEMA_signal_18828), .Z1_f (new_AGEMA_signal_18829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_102_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_102_MUX_inst_Y), .A0_f (new_AGEMA_signal_18827), .A1_t (new_AGEMA_signal_18828), .A1_f (new_AGEMA_signal_18829), .B0_t (RoundOutput[102]), .B0_f (new_AGEMA_signal_17255), .B1_t (new_AGEMA_signal_17256), .B1_f (new_AGEMA_signal_17257), .Z0_t (RoundInput[102]), .Z0_f (new_AGEMA_signal_5087), .Z1_t (new_AGEMA_signal_5088), .Z1_f (new_AGEMA_signal_5089) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_103_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[103]), .A0_f (new_AGEMA_signal_17258), .A1_t (new_AGEMA_signal_17259), .A1_f (new_AGEMA_signal_17260), .B0_t (plaintext_s0_t[103]), .B0_f (plaintext_s0_f[103]), .B1_t (plaintext_s1_t[103]), .B1_f (plaintext_s1_f[103]), .Z0_t (RoundReg_Inst_ff_SDE_103_MUX_inst_X), .Z0_f (new_AGEMA_signal_18290), .Z1_t (new_AGEMA_signal_18291), .Z1_f (new_AGEMA_signal_18292) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_103_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_103_MUX_inst_X), .B0_f (new_AGEMA_signal_18290), .B1_t (new_AGEMA_signal_18291), .B1_f (new_AGEMA_signal_18292), .Z0_t (RoundReg_Inst_ff_SDE_103_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18830), .Z1_t (new_AGEMA_signal_18831), .Z1_f (new_AGEMA_signal_18832) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_103_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_103_MUX_inst_Y), .A0_f (new_AGEMA_signal_18830), .A1_t (new_AGEMA_signal_18831), .A1_f (new_AGEMA_signal_18832), .B0_t (RoundOutput[103]), .B0_f (new_AGEMA_signal_17258), .B1_t (new_AGEMA_signal_17259), .B1_f (new_AGEMA_signal_17260), .Z0_t (RoundInput[103]), .Z0_f (new_AGEMA_signal_5096), .Z1_t (new_AGEMA_signal_5097), .Z1_f (new_AGEMA_signal_5098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_104_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[104]), .A0_f (new_AGEMA_signal_17261), .A1_t (new_AGEMA_signal_17262), .A1_f (new_AGEMA_signal_17263), .B0_t (plaintext_s0_t[104]), .B0_f (plaintext_s0_f[104]), .B1_t (plaintext_s1_t[104]), .B1_f (plaintext_s1_f[104]), .Z0_t (RoundReg_Inst_ff_SDE_104_MUX_inst_X), .Z0_f (new_AGEMA_signal_18296), .Z1_t (new_AGEMA_signal_18297), .Z1_f (new_AGEMA_signal_18298) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_104_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_104_MUX_inst_X), .B0_f (new_AGEMA_signal_18296), .B1_t (new_AGEMA_signal_18297), .B1_f (new_AGEMA_signal_18298), .Z0_t (RoundReg_Inst_ff_SDE_104_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18833), .Z1_t (new_AGEMA_signal_18834), .Z1_f (new_AGEMA_signal_18835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_104_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_104_MUX_inst_Y), .A0_f (new_AGEMA_signal_18833), .A1_t (new_AGEMA_signal_18834), .A1_f (new_AGEMA_signal_18835), .B0_t (RoundOutput[104]), .B0_f (new_AGEMA_signal_17261), .B1_t (new_AGEMA_signal_17262), .B1_f (new_AGEMA_signal_17263), .Z0_t (RoundInput[104]), .Z0_f (new_AGEMA_signal_5105), .Z1_t (new_AGEMA_signal_5106), .Z1_f (new_AGEMA_signal_5107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_105_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[105]), .A0_f (new_AGEMA_signal_17762), .A1_t (new_AGEMA_signal_17763), .A1_f (new_AGEMA_signal_17764), .B0_t (plaintext_s0_t[105]), .B0_f (plaintext_s0_f[105]), .B1_t (plaintext_s1_t[105]), .B1_f (plaintext_s1_f[105]), .Z0_t (RoundReg_Inst_ff_SDE_105_MUX_inst_X), .Z0_f (new_AGEMA_signal_18839), .Z1_t (new_AGEMA_signal_18840), .Z1_f (new_AGEMA_signal_18841) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_105_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_105_MUX_inst_X), .B0_f (new_AGEMA_signal_18839), .B1_t (new_AGEMA_signal_18840), .B1_f (new_AGEMA_signal_18841), .Z0_t (RoundReg_Inst_ff_SDE_105_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19049), .Z1_t (new_AGEMA_signal_19050), .Z1_f (new_AGEMA_signal_19051) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_105_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_105_MUX_inst_Y), .A0_f (new_AGEMA_signal_19049), .A1_t (new_AGEMA_signal_19050), .A1_f (new_AGEMA_signal_19051), .B0_t (RoundOutput[105]), .B0_f (new_AGEMA_signal_17762), .B1_t (new_AGEMA_signal_17763), .B1_f (new_AGEMA_signal_17764), .Z0_t (RoundInput[105]), .Z0_f (new_AGEMA_signal_5114), .Z1_t (new_AGEMA_signal_5115), .Z1_f (new_AGEMA_signal_5116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_106_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[106]), .A0_f (new_AGEMA_signal_17267), .A1_t (new_AGEMA_signal_17268), .A1_f (new_AGEMA_signal_17269), .B0_t (plaintext_s0_t[106]), .B0_f (plaintext_s0_f[106]), .B1_t (plaintext_s1_t[106]), .B1_f (plaintext_s1_f[106]), .Z0_t (RoundReg_Inst_ff_SDE_106_MUX_inst_X), .Z0_f (new_AGEMA_signal_18302), .Z1_t (new_AGEMA_signal_18303), .Z1_f (new_AGEMA_signal_18304) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_106_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_106_MUX_inst_X), .B0_f (new_AGEMA_signal_18302), .B1_t (new_AGEMA_signal_18303), .B1_f (new_AGEMA_signal_18304), .Z0_t (RoundReg_Inst_ff_SDE_106_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18842), .Z1_t (new_AGEMA_signal_18843), .Z1_f (new_AGEMA_signal_18844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_106_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_106_MUX_inst_Y), .A0_f (new_AGEMA_signal_18842), .A1_t (new_AGEMA_signal_18843), .A1_f (new_AGEMA_signal_18844), .B0_t (RoundOutput[106]), .B0_f (new_AGEMA_signal_17267), .B1_t (new_AGEMA_signal_17268), .B1_f (new_AGEMA_signal_17269), .Z0_t (RoundInput[106]), .Z0_f (new_AGEMA_signal_5123), .Z1_t (new_AGEMA_signal_5124), .Z1_f (new_AGEMA_signal_5125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_107_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[107]), .A0_f (new_AGEMA_signal_17765), .A1_t (new_AGEMA_signal_17766), .A1_f (new_AGEMA_signal_17767), .B0_t (plaintext_s0_t[107]), .B0_f (plaintext_s0_f[107]), .B1_t (plaintext_s1_t[107]), .B1_f (plaintext_s1_f[107]), .Z0_t (RoundReg_Inst_ff_SDE_107_MUX_inst_X), .Z0_f (new_AGEMA_signal_18848), .Z1_t (new_AGEMA_signal_18849), .Z1_f (new_AGEMA_signal_18850) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_107_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_107_MUX_inst_X), .B0_f (new_AGEMA_signal_18848), .B1_t (new_AGEMA_signal_18849), .B1_f (new_AGEMA_signal_18850), .Z0_t (RoundReg_Inst_ff_SDE_107_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19052), .Z1_t (new_AGEMA_signal_19053), .Z1_f (new_AGEMA_signal_19054) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_107_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_107_MUX_inst_Y), .A0_f (new_AGEMA_signal_19052), .A1_t (new_AGEMA_signal_19053), .A1_f (new_AGEMA_signal_19054), .B0_t (RoundOutput[107]), .B0_f (new_AGEMA_signal_17765), .B1_t (new_AGEMA_signal_17766), .B1_f (new_AGEMA_signal_17767), .Z0_t (RoundInput[107]), .Z0_f (new_AGEMA_signal_5132), .Z1_t (new_AGEMA_signal_5133), .Z1_f (new_AGEMA_signal_5134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_108_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[108]), .A0_f (new_AGEMA_signal_17768), .A1_t (new_AGEMA_signal_17769), .A1_f (new_AGEMA_signal_17770), .B0_t (plaintext_s0_t[108]), .B0_f (plaintext_s0_f[108]), .B1_t (plaintext_s1_t[108]), .B1_f (plaintext_s1_f[108]), .Z0_t (RoundReg_Inst_ff_SDE_108_MUX_inst_X), .Z0_f (new_AGEMA_signal_18854), .Z1_t (new_AGEMA_signal_18855), .Z1_f (new_AGEMA_signal_18856) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_108_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_108_MUX_inst_X), .B0_f (new_AGEMA_signal_18854), .B1_t (new_AGEMA_signal_18855), .B1_f (new_AGEMA_signal_18856), .Z0_t (RoundReg_Inst_ff_SDE_108_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19055), .Z1_t (new_AGEMA_signal_19056), .Z1_f (new_AGEMA_signal_19057) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_108_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_108_MUX_inst_Y), .A0_f (new_AGEMA_signal_19055), .A1_t (new_AGEMA_signal_19056), .A1_f (new_AGEMA_signal_19057), .B0_t (RoundOutput[108]), .B0_f (new_AGEMA_signal_17768), .B1_t (new_AGEMA_signal_17769), .B1_f (new_AGEMA_signal_17770), .Z0_t (RoundInput[108]), .Z0_f (new_AGEMA_signal_5141), .Z1_t (new_AGEMA_signal_5142), .Z1_f (new_AGEMA_signal_5143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_109_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[109]), .A0_f (new_AGEMA_signal_17276), .A1_t (new_AGEMA_signal_17277), .A1_f (new_AGEMA_signal_17278), .B0_t (plaintext_s0_t[109]), .B0_f (plaintext_s0_f[109]), .B1_t (plaintext_s1_t[109]), .B1_f (plaintext_s1_f[109]), .Z0_t (RoundReg_Inst_ff_SDE_109_MUX_inst_X), .Z0_f (new_AGEMA_signal_18308), .Z1_t (new_AGEMA_signal_18309), .Z1_f (new_AGEMA_signal_18310) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_109_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_109_MUX_inst_X), .B0_f (new_AGEMA_signal_18308), .B1_t (new_AGEMA_signal_18309), .B1_f (new_AGEMA_signal_18310), .Z0_t (RoundReg_Inst_ff_SDE_109_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18857), .Z1_t (new_AGEMA_signal_18858), .Z1_f (new_AGEMA_signal_18859) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_109_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_109_MUX_inst_Y), .A0_f (new_AGEMA_signal_18857), .A1_t (new_AGEMA_signal_18858), .A1_f (new_AGEMA_signal_18859), .B0_t (RoundOutput[109]), .B0_f (new_AGEMA_signal_17276), .B1_t (new_AGEMA_signal_17277), .B1_f (new_AGEMA_signal_17278), .Z0_t (RoundInput[109]), .Z0_f (new_AGEMA_signal_5150), .Z1_t (new_AGEMA_signal_5151), .Z1_f (new_AGEMA_signal_5152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_110_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[110]), .A0_f (new_AGEMA_signal_17282), .A1_t (new_AGEMA_signal_17283), .A1_f (new_AGEMA_signal_17284), .B0_t (plaintext_s0_t[110]), .B0_f (plaintext_s0_f[110]), .B1_t (plaintext_s1_t[110]), .B1_f (plaintext_s1_f[110]), .Z0_t (RoundReg_Inst_ff_SDE_110_MUX_inst_X), .Z0_f (new_AGEMA_signal_18314), .Z1_t (new_AGEMA_signal_18315), .Z1_f (new_AGEMA_signal_18316) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_110_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_110_MUX_inst_X), .B0_f (new_AGEMA_signal_18314), .B1_t (new_AGEMA_signal_18315), .B1_f (new_AGEMA_signal_18316), .Z0_t (RoundReg_Inst_ff_SDE_110_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18860), .Z1_t (new_AGEMA_signal_18861), .Z1_f (new_AGEMA_signal_18862) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_110_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_110_MUX_inst_Y), .A0_f (new_AGEMA_signal_18860), .A1_t (new_AGEMA_signal_18861), .A1_f (new_AGEMA_signal_18862), .B0_t (RoundOutput[110]), .B0_f (new_AGEMA_signal_17282), .B1_t (new_AGEMA_signal_17283), .B1_f (new_AGEMA_signal_17284), .Z0_t (RoundInput[110]), .Z0_f (new_AGEMA_signal_5168), .Z1_t (new_AGEMA_signal_5169), .Z1_f (new_AGEMA_signal_5170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_111_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[111]), .A0_f (new_AGEMA_signal_17285), .A1_t (new_AGEMA_signal_17286), .A1_f (new_AGEMA_signal_17287), .B0_t (plaintext_s0_t[111]), .B0_f (plaintext_s0_f[111]), .B1_t (plaintext_s1_t[111]), .B1_f (plaintext_s1_f[111]), .Z0_t (RoundReg_Inst_ff_SDE_111_MUX_inst_X), .Z0_f (new_AGEMA_signal_18320), .Z1_t (new_AGEMA_signal_18321), .Z1_f (new_AGEMA_signal_18322) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_111_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_111_MUX_inst_X), .B0_f (new_AGEMA_signal_18320), .B1_t (new_AGEMA_signal_18321), .B1_f (new_AGEMA_signal_18322), .Z0_t (RoundReg_Inst_ff_SDE_111_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18863), .Z1_t (new_AGEMA_signal_18864), .Z1_f (new_AGEMA_signal_18865) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_111_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_111_MUX_inst_Y), .A0_f (new_AGEMA_signal_18863), .A1_t (new_AGEMA_signal_18864), .A1_f (new_AGEMA_signal_18865), .B0_t (RoundOutput[111]), .B0_f (new_AGEMA_signal_17285), .B1_t (new_AGEMA_signal_17286), .B1_f (new_AGEMA_signal_17287), .Z0_t (RoundInput[111]), .Z0_f (new_AGEMA_signal_5177), .Z1_t (new_AGEMA_signal_5178), .Z1_f (new_AGEMA_signal_5179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_112_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[112]), .A0_f (new_AGEMA_signal_17288), .A1_t (new_AGEMA_signal_17289), .A1_f (new_AGEMA_signal_17290), .B0_t (plaintext_s0_t[112]), .B0_f (plaintext_s0_f[112]), .B1_t (plaintext_s1_t[112]), .B1_f (plaintext_s1_f[112]), .Z0_t (RoundReg_Inst_ff_SDE_112_MUX_inst_X), .Z0_f (new_AGEMA_signal_18326), .Z1_t (new_AGEMA_signal_18327), .Z1_f (new_AGEMA_signal_18328) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_112_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_112_MUX_inst_X), .B0_f (new_AGEMA_signal_18326), .B1_t (new_AGEMA_signal_18327), .B1_f (new_AGEMA_signal_18328), .Z0_t (RoundReg_Inst_ff_SDE_112_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18866), .Z1_t (new_AGEMA_signal_18867), .Z1_f (new_AGEMA_signal_18868) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_112_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_112_MUX_inst_Y), .A0_f (new_AGEMA_signal_18866), .A1_t (new_AGEMA_signal_18867), .A1_f (new_AGEMA_signal_18868), .B0_t (RoundOutput[112]), .B0_f (new_AGEMA_signal_17288), .B1_t (new_AGEMA_signal_17289), .B1_f (new_AGEMA_signal_17290), .Z0_t (RoundInput[112]), .Z0_f (new_AGEMA_signal_5186), .Z1_t (new_AGEMA_signal_5187), .Z1_f (new_AGEMA_signal_5188) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_113_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[113]), .A0_f (new_AGEMA_signal_17771), .A1_t (new_AGEMA_signal_17772), .A1_f (new_AGEMA_signal_17773), .B0_t (plaintext_s0_t[113]), .B0_f (plaintext_s0_f[113]), .B1_t (plaintext_s1_t[113]), .B1_f (plaintext_s1_f[113]), .Z0_t (RoundReg_Inst_ff_SDE_113_MUX_inst_X), .Z0_f (new_AGEMA_signal_18872), .Z1_t (new_AGEMA_signal_18873), .Z1_f (new_AGEMA_signal_18874) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_113_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_113_MUX_inst_X), .B0_f (new_AGEMA_signal_18872), .B1_t (new_AGEMA_signal_18873), .B1_f (new_AGEMA_signal_18874), .Z0_t (RoundReg_Inst_ff_SDE_113_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19058), .Z1_t (new_AGEMA_signal_19059), .Z1_f (new_AGEMA_signal_19060) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_113_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_113_MUX_inst_Y), .A0_f (new_AGEMA_signal_19058), .A1_t (new_AGEMA_signal_19059), .A1_f (new_AGEMA_signal_19060), .B0_t (RoundOutput[113]), .B0_f (new_AGEMA_signal_17771), .B1_t (new_AGEMA_signal_17772), .B1_f (new_AGEMA_signal_17773), .Z0_t (RoundInput[113]), .Z0_f (new_AGEMA_signal_5195), .Z1_t (new_AGEMA_signal_5196), .Z1_f (new_AGEMA_signal_5197) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_114_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[114]), .A0_f (new_AGEMA_signal_17294), .A1_t (new_AGEMA_signal_17295), .A1_f (new_AGEMA_signal_17296), .B0_t (plaintext_s0_t[114]), .B0_f (plaintext_s0_f[114]), .B1_t (plaintext_s1_t[114]), .B1_f (plaintext_s1_f[114]), .Z0_t (RoundReg_Inst_ff_SDE_114_MUX_inst_X), .Z0_f (new_AGEMA_signal_18332), .Z1_t (new_AGEMA_signal_18333), .Z1_f (new_AGEMA_signal_18334) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_114_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_114_MUX_inst_X), .B0_f (new_AGEMA_signal_18332), .B1_t (new_AGEMA_signal_18333), .B1_f (new_AGEMA_signal_18334), .Z0_t (RoundReg_Inst_ff_SDE_114_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18875), .Z1_t (new_AGEMA_signal_18876), .Z1_f (new_AGEMA_signal_18877) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_114_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_114_MUX_inst_Y), .A0_f (new_AGEMA_signal_18875), .A1_t (new_AGEMA_signal_18876), .A1_f (new_AGEMA_signal_18877), .B0_t (RoundOutput[114]), .B0_f (new_AGEMA_signal_17294), .B1_t (new_AGEMA_signal_17295), .B1_f (new_AGEMA_signal_17296), .Z0_t (RoundInput[114]), .Z0_f (new_AGEMA_signal_5204), .Z1_t (new_AGEMA_signal_5205), .Z1_f (new_AGEMA_signal_5206) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_115_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[115]), .A0_f (new_AGEMA_signal_17774), .A1_t (new_AGEMA_signal_17775), .A1_f (new_AGEMA_signal_17776), .B0_t (plaintext_s0_t[115]), .B0_f (plaintext_s0_f[115]), .B1_t (plaintext_s1_t[115]), .B1_f (plaintext_s1_f[115]), .Z0_t (RoundReg_Inst_ff_SDE_115_MUX_inst_X), .Z0_f (new_AGEMA_signal_18881), .Z1_t (new_AGEMA_signal_18882), .Z1_f (new_AGEMA_signal_18883) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_115_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_115_MUX_inst_X), .B0_f (new_AGEMA_signal_18881), .B1_t (new_AGEMA_signal_18882), .B1_f (new_AGEMA_signal_18883), .Z0_t (RoundReg_Inst_ff_SDE_115_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19061), .Z1_t (new_AGEMA_signal_19062), .Z1_f (new_AGEMA_signal_19063) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_115_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_115_MUX_inst_Y), .A0_f (new_AGEMA_signal_19061), .A1_t (new_AGEMA_signal_19062), .A1_f (new_AGEMA_signal_19063), .B0_t (RoundOutput[115]), .B0_f (new_AGEMA_signal_17774), .B1_t (new_AGEMA_signal_17775), .B1_f (new_AGEMA_signal_17776), .Z0_t (RoundInput[115]), .Z0_f (new_AGEMA_signal_5213), .Z1_t (new_AGEMA_signal_5214), .Z1_f (new_AGEMA_signal_5215) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_116_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[116]), .A0_f (new_AGEMA_signal_17777), .A1_t (new_AGEMA_signal_17778), .A1_f (new_AGEMA_signal_17779), .B0_t (plaintext_s0_t[116]), .B0_f (plaintext_s0_f[116]), .B1_t (plaintext_s1_t[116]), .B1_f (plaintext_s1_f[116]), .Z0_t (RoundReg_Inst_ff_SDE_116_MUX_inst_X), .Z0_f (new_AGEMA_signal_18887), .Z1_t (new_AGEMA_signal_18888), .Z1_f (new_AGEMA_signal_18889) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_116_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_116_MUX_inst_X), .B0_f (new_AGEMA_signal_18887), .B1_t (new_AGEMA_signal_18888), .B1_f (new_AGEMA_signal_18889), .Z0_t (RoundReg_Inst_ff_SDE_116_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19064), .Z1_t (new_AGEMA_signal_19065), .Z1_f (new_AGEMA_signal_19066) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_116_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_116_MUX_inst_Y), .A0_f (new_AGEMA_signal_19064), .A1_t (new_AGEMA_signal_19065), .A1_f (new_AGEMA_signal_19066), .B0_t (RoundOutput[116]), .B0_f (new_AGEMA_signal_17777), .B1_t (new_AGEMA_signal_17778), .B1_f (new_AGEMA_signal_17779), .Z0_t (RoundInput[116]), .Z0_f (new_AGEMA_signal_5222), .Z1_t (new_AGEMA_signal_5223), .Z1_f (new_AGEMA_signal_5224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_117_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[117]), .A0_f (new_AGEMA_signal_17303), .A1_t (new_AGEMA_signal_17304), .A1_f (new_AGEMA_signal_17305), .B0_t (plaintext_s0_t[117]), .B0_f (plaintext_s0_f[117]), .B1_t (plaintext_s1_t[117]), .B1_f (plaintext_s1_f[117]), .Z0_t (RoundReg_Inst_ff_SDE_117_MUX_inst_X), .Z0_f (new_AGEMA_signal_18338), .Z1_t (new_AGEMA_signal_18339), .Z1_f (new_AGEMA_signal_18340) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_117_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_117_MUX_inst_X), .B0_f (new_AGEMA_signal_18338), .B1_t (new_AGEMA_signal_18339), .B1_f (new_AGEMA_signal_18340), .Z0_t (RoundReg_Inst_ff_SDE_117_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18890), .Z1_t (new_AGEMA_signal_18891), .Z1_f (new_AGEMA_signal_18892) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_117_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_117_MUX_inst_Y), .A0_f (new_AGEMA_signal_18890), .A1_t (new_AGEMA_signal_18891), .A1_f (new_AGEMA_signal_18892), .B0_t (RoundOutput[117]), .B0_f (new_AGEMA_signal_17303), .B1_t (new_AGEMA_signal_17304), .B1_f (new_AGEMA_signal_17305), .Z0_t (RoundInput[117]), .Z0_f (new_AGEMA_signal_5231), .Z1_t (new_AGEMA_signal_5232), .Z1_f (new_AGEMA_signal_5233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_118_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[118]), .A0_f (new_AGEMA_signal_17306), .A1_t (new_AGEMA_signal_17307), .A1_f (new_AGEMA_signal_17308), .B0_t (plaintext_s0_t[118]), .B0_f (plaintext_s0_f[118]), .B1_t (plaintext_s1_t[118]), .B1_f (plaintext_s1_f[118]), .Z0_t (RoundReg_Inst_ff_SDE_118_MUX_inst_X), .Z0_f (new_AGEMA_signal_18344), .Z1_t (new_AGEMA_signal_18345), .Z1_f (new_AGEMA_signal_18346) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_118_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_118_MUX_inst_X), .B0_f (new_AGEMA_signal_18344), .B1_t (new_AGEMA_signal_18345), .B1_f (new_AGEMA_signal_18346), .Z0_t (RoundReg_Inst_ff_SDE_118_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18893), .Z1_t (new_AGEMA_signal_18894), .Z1_f (new_AGEMA_signal_18895) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_118_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_118_MUX_inst_Y), .A0_f (new_AGEMA_signal_18893), .A1_t (new_AGEMA_signal_18894), .A1_f (new_AGEMA_signal_18895), .B0_t (RoundOutput[118]), .B0_f (new_AGEMA_signal_17306), .B1_t (new_AGEMA_signal_17307), .B1_f (new_AGEMA_signal_17308), .Z0_t (RoundInput[118]), .Z0_f (new_AGEMA_signal_5240), .Z1_t (new_AGEMA_signal_5241), .Z1_f (new_AGEMA_signal_5242) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_119_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[119]), .A0_f (new_AGEMA_signal_17309), .A1_t (new_AGEMA_signal_17310), .A1_f (new_AGEMA_signal_17311), .B0_t (plaintext_s0_t[119]), .B0_f (plaintext_s0_f[119]), .B1_t (plaintext_s1_t[119]), .B1_f (plaintext_s1_f[119]), .Z0_t (RoundReg_Inst_ff_SDE_119_MUX_inst_X), .Z0_f (new_AGEMA_signal_18350), .Z1_t (new_AGEMA_signal_18351), .Z1_f (new_AGEMA_signal_18352) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_119_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_119_MUX_inst_X), .B0_f (new_AGEMA_signal_18350), .B1_t (new_AGEMA_signal_18351), .B1_f (new_AGEMA_signal_18352), .Z0_t (RoundReg_Inst_ff_SDE_119_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18896), .Z1_t (new_AGEMA_signal_18897), .Z1_f (new_AGEMA_signal_18898) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_119_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_119_MUX_inst_Y), .A0_f (new_AGEMA_signal_18896), .A1_t (new_AGEMA_signal_18897), .A1_f (new_AGEMA_signal_18898), .B0_t (RoundOutput[119]), .B0_f (new_AGEMA_signal_17309), .B1_t (new_AGEMA_signal_17310), .B1_f (new_AGEMA_signal_17311), .Z0_t (RoundInput[119]), .Z0_f (new_AGEMA_signal_5249), .Z1_t (new_AGEMA_signal_5250), .Z1_f (new_AGEMA_signal_5251) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_120_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[120]), .A0_f (new_AGEMA_signal_17315), .A1_t (new_AGEMA_signal_17316), .A1_f (new_AGEMA_signal_17317), .B0_t (plaintext_s0_t[120]), .B0_f (plaintext_s0_f[120]), .B1_t (plaintext_s1_t[120]), .B1_f (plaintext_s1_f[120]), .Z0_t (RoundReg_Inst_ff_SDE_120_MUX_inst_X), .Z0_f (new_AGEMA_signal_18356), .Z1_t (new_AGEMA_signal_18357), .Z1_f (new_AGEMA_signal_18358) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_120_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_120_MUX_inst_X), .B0_f (new_AGEMA_signal_18356), .B1_t (new_AGEMA_signal_18357), .B1_f (new_AGEMA_signal_18358), .Z0_t (RoundReg_Inst_ff_SDE_120_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18899), .Z1_t (new_AGEMA_signal_18900), .Z1_f (new_AGEMA_signal_18901) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_120_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_120_MUX_inst_Y), .A0_f (new_AGEMA_signal_18899), .A1_t (new_AGEMA_signal_18900), .A1_f (new_AGEMA_signal_18901), .B0_t (RoundOutput[120]), .B0_f (new_AGEMA_signal_17315), .B1_t (new_AGEMA_signal_17316), .B1_f (new_AGEMA_signal_17317), .Z0_t (RoundInput[120]), .Z0_f (new_AGEMA_signal_5267), .Z1_t (new_AGEMA_signal_5268), .Z1_f (new_AGEMA_signal_5269) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_121_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[121]), .A0_f (new_AGEMA_signal_17783), .A1_t (new_AGEMA_signal_17784), .A1_f (new_AGEMA_signal_17785), .B0_t (plaintext_s0_t[121]), .B0_f (plaintext_s0_f[121]), .B1_t (plaintext_s1_t[121]), .B1_f (plaintext_s1_f[121]), .Z0_t (RoundReg_Inst_ff_SDE_121_MUX_inst_X), .Z0_f (new_AGEMA_signal_18905), .Z1_t (new_AGEMA_signal_18906), .Z1_f (new_AGEMA_signal_18907) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_121_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_121_MUX_inst_X), .B0_f (new_AGEMA_signal_18905), .B1_t (new_AGEMA_signal_18906), .B1_f (new_AGEMA_signal_18907), .Z0_t (RoundReg_Inst_ff_SDE_121_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19067), .Z1_t (new_AGEMA_signal_19068), .Z1_f (new_AGEMA_signal_19069) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_121_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_121_MUX_inst_Y), .A0_f (new_AGEMA_signal_19067), .A1_t (new_AGEMA_signal_19068), .A1_f (new_AGEMA_signal_19069), .B0_t (RoundOutput[121]), .B0_f (new_AGEMA_signal_17783), .B1_t (new_AGEMA_signal_17784), .B1_f (new_AGEMA_signal_17785), .Z0_t (RoundInput[121]), .Z0_f (new_AGEMA_signal_5276), .Z1_t (new_AGEMA_signal_5277), .Z1_f (new_AGEMA_signal_5278) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_122_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[122]), .A0_f (new_AGEMA_signal_17321), .A1_t (new_AGEMA_signal_17322), .A1_f (new_AGEMA_signal_17323), .B0_t (plaintext_s0_t[122]), .B0_f (plaintext_s0_f[122]), .B1_t (plaintext_s1_t[122]), .B1_f (plaintext_s1_f[122]), .Z0_t (RoundReg_Inst_ff_SDE_122_MUX_inst_X), .Z0_f (new_AGEMA_signal_18362), .Z1_t (new_AGEMA_signal_18363), .Z1_f (new_AGEMA_signal_18364) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_122_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_122_MUX_inst_X), .B0_f (new_AGEMA_signal_18362), .B1_t (new_AGEMA_signal_18363), .B1_f (new_AGEMA_signal_18364), .Z0_t (RoundReg_Inst_ff_SDE_122_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18908), .Z1_t (new_AGEMA_signal_18909), .Z1_f (new_AGEMA_signal_18910) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_122_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_122_MUX_inst_Y), .A0_f (new_AGEMA_signal_18908), .A1_t (new_AGEMA_signal_18909), .A1_f (new_AGEMA_signal_18910), .B0_t (RoundOutput[122]), .B0_f (new_AGEMA_signal_17321), .B1_t (new_AGEMA_signal_17322), .B1_f (new_AGEMA_signal_17323), .Z0_t (RoundInput[122]), .Z0_f (new_AGEMA_signal_5285), .Z1_t (new_AGEMA_signal_5286), .Z1_f (new_AGEMA_signal_5287) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_123_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[123]), .A0_f (new_AGEMA_signal_17786), .A1_t (new_AGEMA_signal_17787), .A1_f (new_AGEMA_signal_17788), .B0_t (plaintext_s0_t[123]), .B0_f (plaintext_s0_f[123]), .B1_t (plaintext_s1_t[123]), .B1_f (plaintext_s1_f[123]), .Z0_t (RoundReg_Inst_ff_SDE_123_MUX_inst_X), .Z0_f (new_AGEMA_signal_18914), .Z1_t (new_AGEMA_signal_18915), .Z1_f (new_AGEMA_signal_18916) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_123_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_123_MUX_inst_X), .B0_f (new_AGEMA_signal_18914), .B1_t (new_AGEMA_signal_18915), .B1_f (new_AGEMA_signal_18916), .Z0_t (RoundReg_Inst_ff_SDE_123_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19070), .Z1_t (new_AGEMA_signal_19071), .Z1_f (new_AGEMA_signal_19072) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_123_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_123_MUX_inst_Y), .A0_f (new_AGEMA_signal_19070), .A1_t (new_AGEMA_signal_19071), .A1_f (new_AGEMA_signal_19072), .B0_t (RoundOutput[123]), .B0_f (new_AGEMA_signal_17786), .B1_t (new_AGEMA_signal_17787), .B1_f (new_AGEMA_signal_17788), .Z0_t (RoundInput[123]), .Z0_f (new_AGEMA_signal_5294), .Z1_t (new_AGEMA_signal_5295), .Z1_f (new_AGEMA_signal_5296) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_124_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[124]), .A0_f (new_AGEMA_signal_17789), .A1_t (new_AGEMA_signal_17790), .A1_f (new_AGEMA_signal_17791), .B0_t (plaintext_s0_t[124]), .B0_f (plaintext_s0_f[124]), .B1_t (plaintext_s1_t[124]), .B1_f (plaintext_s1_f[124]), .Z0_t (RoundReg_Inst_ff_SDE_124_MUX_inst_X), .Z0_f (new_AGEMA_signal_18920), .Z1_t (new_AGEMA_signal_18921), .Z1_f (new_AGEMA_signal_18922) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_124_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_124_MUX_inst_X), .B0_f (new_AGEMA_signal_18920), .B1_t (new_AGEMA_signal_18921), .B1_f (new_AGEMA_signal_18922), .Z0_t (RoundReg_Inst_ff_SDE_124_MUX_inst_Y), .Z0_f (new_AGEMA_signal_19073), .Z1_t (new_AGEMA_signal_19074), .Z1_f (new_AGEMA_signal_19075) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_124_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_124_MUX_inst_Y), .A0_f (new_AGEMA_signal_19073), .A1_t (new_AGEMA_signal_19074), .A1_f (new_AGEMA_signal_19075), .B0_t (RoundOutput[124]), .B0_f (new_AGEMA_signal_17789), .B1_t (new_AGEMA_signal_17790), .B1_f (new_AGEMA_signal_17791), .Z0_t (RoundInput[124]), .Z0_f (new_AGEMA_signal_5303), .Z1_t (new_AGEMA_signal_5304), .Z1_f (new_AGEMA_signal_5305) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_125_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[125]), .A0_f (new_AGEMA_signal_17330), .A1_t (new_AGEMA_signal_17331), .A1_f (new_AGEMA_signal_17332), .B0_t (plaintext_s0_t[125]), .B0_f (plaintext_s0_f[125]), .B1_t (plaintext_s1_t[125]), .B1_f (plaintext_s1_f[125]), .Z0_t (RoundReg_Inst_ff_SDE_125_MUX_inst_X), .Z0_f (new_AGEMA_signal_18368), .Z1_t (new_AGEMA_signal_18369), .Z1_f (new_AGEMA_signal_18370) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_125_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_125_MUX_inst_X), .B0_f (new_AGEMA_signal_18368), .B1_t (new_AGEMA_signal_18369), .B1_f (new_AGEMA_signal_18370), .Z0_t (RoundReg_Inst_ff_SDE_125_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18923), .Z1_t (new_AGEMA_signal_18924), .Z1_f (new_AGEMA_signal_18925) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_125_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_125_MUX_inst_Y), .A0_f (new_AGEMA_signal_18923), .A1_t (new_AGEMA_signal_18924), .A1_f (new_AGEMA_signal_18925), .B0_t (RoundOutput[125]), .B0_f (new_AGEMA_signal_17330), .B1_t (new_AGEMA_signal_17331), .B1_f (new_AGEMA_signal_17332), .Z0_t (RoundInput[125]), .Z0_f (new_AGEMA_signal_5312), .Z1_t (new_AGEMA_signal_5313), .Z1_f (new_AGEMA_signal_5314) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_126_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[126]), .A0_f (new_AGEMA_signal_17333), .A1_t (new_AGEMA_signal_17334), .A1_f (new_AGEMA_signal_17335), .B0_t (plaintext_s0_t[126]), .B0_f (plaintext_s0_f[126]), .B1_t (plaintext_s1_t[126]), .B1_f (plaintext_s1_f[126]), .Z0_t (RoundReg_Inst_ff_SDE_126_MUX_inst_X), .Z0_f (new_AGEMA_signal_18374), .Z1_t (new_AGEMA_signal_18375), .Z1_f (new_AGEMA_signal_18376) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_126_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_126_MUX_inst_X), .B0_f (new_AGEMA_signal_18374), .B1_t (new_AGEMA_signal_18375), .B1_f (new_AGEMA_signal_18376), .Z0_t (RoundReg_Inst_ff_SDE_126_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18926), .Z1_t (new_AGEMA_signal_18927), .Z1_f (new_AGEMA_signal_18928) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_126_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_126_MUX_inst_Y), .A0_f (new_AGEMA_signal_18926), .A1_t (new_AGEMA_signal_18927), .A1_f (new_AGEMA_signal_18928), .B0_t (RoundOutput[126]), .B0_f (new_AGEMA_signal_17333), .B1_t (new_AGEMA_signal_17334), .B1_f (new_AGEMA_signal_17335), .Z0_t (RoundInput[126]), .Z0_f (new_AGEMA_signal_5321), .Z1_t (new_AGEMA_signal_5322), .Z1_f (new_AGEMA_signal_5323) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_127_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[127]), .A0_f (new_AGEMA_signal_17336), .A1_t (new_AGEMA_signal_17337), .A1_f (new_AGEMA_signal_17338), .B0_t (plaintext_s0_t[127]), .B0_f (plaintext_s0_f[127]), .B1_t (plaintext_s1_t[127]), .B1_f (plaintext_s1_f[127]), .Z0_t (RoundReg_Inst_ff_SDE_127_MUX_inst_X), .Z0_f (new_AGEMA_signal_18380), .Z1_t (new_AGEMA_signal_18381), .Z1_f (new_AGEMA_signal_18382) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_127_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (RoundReg_Inst_ff_SDE_127_MUX_inst_X), .B0_f (new_AGEMA_signal_18380), .B1_t (new_AGEMA_signal_18381), .B1_f (new_AGEMA_signal_18382), .Z0_t (RoundReg_Inst_ff_SDE_127_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18929), .Z1_t (new_AGEMA_signal_18930), .Z1_f (new_AGEMA_signal_18931) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_127_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_127_MUX_inst_Y), .A0_f (new_AGEMA_signal_18929), .A1_t (new_AGEMA_signal_18930), .A1_f (new_AGEMA_signal_18931), .B0_t (RoundOutput[127]), .B0_f (new_AGEMA_signal_17336), .B1_t (new_AGEMA_signal_17337), .B1_f (new_AGEMA_signal_17338), .Z0_t (RoundInput[127]), .Z0_f (new_AGEMA_signal_5330), .Z1_t (new_AGEMA_signal_5331), .Z1_f (new_AGEMA_signal_5332) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[7]), .A0_f (ciphertext_s0_f[7]), .A1_t (ciphertext_s1_t[7]), .A1_f (ciphertext_s1_f[7]), .B0_t (ciphertext_s0_t[4]), .B0_f (ciphertext_s0_f[4]), .B1_t (ciphertext_s1_t[4]), .B1_f (ciphertext_s1_f[4]), .Z0_t (SubBytesIns_Inst_Sbox_0_T1), .Z0_f (new_AGEMA_signal_6346), .Z1_t (new_AGEMA_signal_6347), .Z1_f (new_AGEMA_signal_6348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[7]), .A0_f (ciphertext_s0_f[7]), .A1_t (ciphertext_s1_t[7]), .A1_f (ciphertext_s1_f[7]), .B0_t (ciphertext_s0_t[2]), .B0_f (ciphertext_s0_f[2]), .B1_t (ciphertext_s1_t[2]), .B1_f (ciphertext_s1_f[2]), .Z0_t (SubBytesIns_Inst_Sbox_0_T2), .Z0_f (new_AGEMA_signal_6349), .Z1_t (new_AGEMA_signal_6350), .Z1_f (new_AGEMA_signal_6351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[7]), .A0_f (ciphertext_s0_f[7]), .A1_t (ciphertext_s1_t[7]), .A1_f (ciphertext_s1_f[7]), .B0_t (ciphertext_s0_t[1]), .B0_f (ciphertext_s0_f[1]), .B1_t (ciphertext_s1_t[1]), .B1_f (ciphertext_s1_f[1]), .Z0_t (SubBytesIns_Inst_Sbox_0_T3), .Z0_f (new_AGEMA_signal_6352), .Z1_t (new_AGEMA_signal_6353), .Z1_f (new_AGEMA_signal_6354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[4]), .A0_f (ciphertext_s0_f[4]), .A1_t (ciphertext_s1_t[4]), .A1_f (ciphertext_s1_f[4]), .B0_t (ciphertext_s0_t[2]), .B0_f (ciphertext_s0_f[2]), .B1_t (ciphertext_s1_t[2]), .B1_f (ciphertext_s1_f[2]), .Z0_t (SubBytesIns_Inst_Sbox_0_T4), .Z0_f (new_AGEMA_signal_6355), .Z1_t (new_AGEMA_signal_6356), .Z1_f (new_AGEMA_signal_6357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[3]), .A0_f (ciphertext_s0_f[3]), .A1_t (ciphertext_s1_t[3]), .A1_f (ciphertext_s1_f[3]), .B0_t (ciphertext_s0_t[1]), .B0_f (ciphertext_s0_f[1]), .B1_t (ciphertext_s1_t[1]), .B1_f (ciphertext_s1_f[1]), .Z0_t (SubBytesIns_Inst_Sbox_0_T5), .Z0_f (new_AGEMA_signal_6358), .Z1_t (new_AGEMA_signal_6359), .Z1_f (new_AGEMA_signal_6360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T1), .A0_f (new_AGEMA_signal_6346), .A1_t (new_AGEMA_signal_6347), .A1_f (new_AGEMA_signal_6348), .B0_t (SubBytesIns_Inst_Sbox_0_T5), .B0_f (new_AGEMA_signal_6358), .B1_t (new_AGEMA_signal_6359), .B1_f (new_AGEMA_signal_6360), .Z0_t (SubBytesIns_Inst_Sbox_0_T6), .Z0_f (new_AGEMA_signal_6928), .Z1_t (new_AGEMA_signal_6929), .Z1_f (new_AGEMA_signal_6930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[6]), .A0_f (ciphertext_s0_f[6]), .A1_t (ciphertext_s1_t[6]), .A1_f (ciphertext_s1_f[6]), .B0_t (ciphertext_s0_t[5]), .B0_f (ciphertext_s0_f[5]), .B1_t (ciphertext_s1_t[5]), .B1_f (ciphertext_s1_f[5]), .Z0_t (SubBytesIns_Inst_Sbox_0_T7), .Z0_f (new_AGEMA_signal_6361), .Z1_t (new_AGEMA_signal_6362), .Z1_f (new_AGEMA_signal_6363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[0]), .A0_f (ciphertext_s0_f[0]), .A1_t (ciphertext_s1_t[0]), .A1_f (ciphertext_s1_f[0]), .B0_t (SubBytesIns_Inst_Sbox_0_T6), .B0_f (new_AGEMA_signal_6928), .B1_t (new_AGEMA_signal_6929), .B1_f (new_AGEMA_signal_6930), .Z0_t (SubBytesIns_Inst_Sbox_0_T8), .Z0_f (new_AGEMA_signal_7472), .Z1_t (new_AGEMA_signal_7473), .Z1_f (new_AGEMA_signal_7474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[0]), .A0_f (ciphertext_s0_f[0]), .A1_t (ciphertext_s1_t[0]), .A1_f (ciphertext_s1_f[0]), .B0_t (SubBytesIns_Inst_Sbox_0_T7), .B0_f (new_AGEMA_signal_6361), .B1_t (new_AGEMA_signal_6362), .B1_f (new_AGEMA_signal_6363), .Z0_t (SubBytesIns_Inst_Sbox_0_T9), .Z0_f (new_AGEMA_signal_6931), .Z1_t (new_AGEMA_signal_6932), .Z1_f (new_AGEMA_signal_6933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T6), .A0_f (new_AGEMA_signal_6928), .A1_t (new_AGEMA_signal_6929), .A1_f (new_AGEMA_signal_6930), .B0_t (SubBytesIns_Inst_Sbox_0_T7), .B0_f (new_AGEMA_signal_6361), .B1_t (new_AGEMA_signal_6362), .B1_f (new_AGEMA_signal_6363), .Z0_t (SubBytesIns_Inst_Sbox_0_T10), .Z0_f (new_AGEMA_signal_7475), .Z1_t (new_AGEMA_signal_7476), .Z1_f (new_AGEMA_signal_7477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[6]), .A0_f (ciphertext_s0_f[6]), .A1_t (ciphertext_s1_t[6]), .A1_f (ciphertext_s1_f[6]), .B0_t (ciphertext_s0_t[2]), .B0_f (ciphertext_s0_f[2]), .B1_t (ciphertext_s1_t[2]), .B1_f (ciphertext_s1_f[2]), .Z0_t (SubBytesIns_Inst_Sbox_0_T11), .Z0_f (new_AGEMA_signal_6364), .Z1_t (new_AGEMA_signal_6365), .Z1_f (new_AGEMA_signal_6366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[5]), .A0_f (ciphertext_s0_f[5]), .A1_t (ciphertext_s1_t[5]), .A1_f (ciphertext_s1_f[5]), .B0_t (ciphertext_s0_t[2]), .B0_f (ciphertext_s0_f[2]), .B1_t (ciphertext_s1_t[2]), .B1_f (ciphertext_s1_f[2]), .Z0_t (SubBytesIns_Inst_Sbox_0_T12), .Z0_f (new_AGEMA_signal_6367), .Z1_t (new_AGEMA_signal_6368), .Z1_f (new_AGEMA_signal_6369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T3), .A0_f (new_AGEMA_signal_6352), .A1_t (new_AGEMA_signal_6353), .A1_f (new_AGEMA_signal_6354), .B0_t (SubBytesIns_Inst_Sbox_0_T4), .B0_f (new_AGEMA_signal_6355), .B1_t (new_AGEMA_signal_6356), .B1_f (new_AGEMA_signal_6357), .Z0_t (SubBytesIns_Inst_Sbox_0_T13), .Z0_f (new_AGEMA_signal_6934), .Z1_t (new_AGEMA_signal_6935), .Z1_f (new_AGEMA_signal_6936) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T6), .A0_f (new_AGEMA_signal_6928), .A1_t (new_AGEMA_signal_6929), .A1_f (new_AGEMA_signal_6930), .B0_t (SubBytesIns_Inst_Sbox_0_T11), .B0_f (new_AGEMA_signal_6364), .B1_t (new_AGEMA_signal_6365), .B1_f (new_AGEMA_signal_6366), .Z0_t (SubBytesIns_Inst_Sbox_0_T14), .Z0_f (new_AGEMA_signal_7478), .Z1_t (new_AGEMA_signal_7479), .Z1_f (new_AGEMA_signal_7480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T5), .A0_f (new_AGEMA_signal_6358), .A1_t (new_AGEMA_signal_6359), .A1_f (new_AGEMA_signal_6360), .B0_t (SubBytesIns_Inst_Sbox_0_T11), .B0_f (new_AGEMA_signal_6364), .B1_t (new_AGEMA_signal_6365), .B1_f (new_AGEMA_signal_6366), .Z0_t (SubBytesIns_Inst_Sbox_0_T15), .Z0_f (new_AGEMA_signal_6937), .Z1_t (new_AGEMA_signal_6938), .Z1_f (new_AGEMA_signal_6939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T5), .A0_f (new_AGEMA_signal_6358), .A1_t (new_AGEMA_signal_6359), .A1_f (new_AGEMA_signal_6360), .B0_t (SubBytesIns_Inst_Sbox_0_T12), .B0_f (new_AGEMA_signal_6367), .B1_t (new_AGEMA_signal_6368), .B1_f (new_AGEMA_signal_6369), .Z0_t (SubBytesIns_Inst_Sbox_0_T16), .Z0_f (new_AGEMA_signal_6940), .Z1_t (new_AGEMA_signal_6941), .Z1_f (new_AGEMA_signal_6942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T9), .A0_f (new_AGEMA_signal_6931), .A1_t (new_AGEMA_signal_6932), .A1_f (new_AGEMA_signal_6933), .B0_t (SubBytesIns_Inst_Sbox_0_T16), .B0_f (new_AGEMA_signal_6940), .B1_t (new_AGEMA_signal_6941), .B1_f (new_AGEMA_signal_6942), .Z0_t (SubBytesIns_Inst_Sbox_0_T17), .Z0_f (new_AGEMA_signal_7481), .Z1_t (new_AGEMA_signal_7482), .Z1_f (new_AGEMA_signal_7483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[4]), .A0_f (ciphertext_s0_f[4]), .A1_t (ciphertext_s1_t[4]), .A1_f (ciphertext_s1_f[4]), .B0_t (ciphertext_s0_t[0]), .B0_f (ciphertext_s0_f[0]), .B1_t (ciphertext_s1_t[0]), .B1_f (ciphertext_s1_f[0]), .Z0_t (SubBytesIns_Inst_Sbox_0_T18), .Z0_f (new_AGEMA_signal_6370), .Z1_t (new_AGEMA_signal_6371), .Z1_f (new_AGEMA_signal_6372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T7), .A0_f (new_AGEMA_signal_6361), .A1_t (new_AGEMA_signal_6362), .A1_f (new_AGEMA_signal_6363), .B0_t (SubBytesIns_Inst_Sbox_0_T18), .B0_f (new_AGEMA_signal_6370), .B1_t (new_AGEMA_signal_6371), .B1_f (new_AGEMA_signal_6372), .Z0_t (SubBytesIns_Inst_Sbox_0_T19), .Z0_f (new_AGEMA_signal_6943), .Z1_t (new_AGEMA_signal_6944), .Z1_f (new_AGEMA_signal_6945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T1), .A0_f (new_AGEMA_signal_6346), .A1_t (new_AGEMA_signal_6347), .A1_f (new_AGEMA_signal_6348), .B0_t (SubBytesIns_Inst_Sbox_0_T19), .B0_f (new_AGEMA_signal_6943), .B1_t (new_AGEMA_signal_6944), .B1_f (new_AGEMA_signal_6945), .Z0_t (SubBytesIns_Inst_Sbox_0_T20), .Z0_f (new_AGEMA_signal_7484), .Z1_t (new_AGEMA_signal_7485), .Z1_f (new_AGEMA_signal_7486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[1]), .A0_f (ciphertext_s0_f[1]), .A1_t (ciphertext_s1_t[1]), .A1_f (ciphertext_s1_f[1]), .B0_t (ciphertext_s0_t[0]), .B0_f (ciphertext_s0_f[0]), .B1_t (ciphertext_s1_t[0]), .B1_f (ciphertext_s1_f[0]), .Z0_t (SubBytesIns_Inst_Sbox_0_T21), .Z0_f (new_AGEMA_signal_6373), .Z1_t (new_AGEMA_signal_6374), .Z1_f (new_AGEMA_signal_6375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T7), .A0_f (new_AGEMA_signal_6361), .A1_t (new_AGEMA_signal_6362), .A1_f (new_AGEMA_signal_6363), .B0_t (SubBytesIns_Inst_Sbox_0_T21), .B0_f (new_AGEMA_signal_6373), .B1_t (new_AGEMA_signal_6374), .B1_f (new_AGEMA_signal_6375), .Z0_t (SubBytesIns_Inst_Sbox_0_T22), .Z0_f (new_AGEMA_signal_6946), .Z1_t (new_AGEMA_signal_6947), .Z1_f (new_AGEMA_signal_6948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T2), .A0_f (new_AGEMA_signal_6349), .A1_t (new_AGEMA_signal_6350), .A1_f (new_AGEMA_signal_6351), .B0_t (SubBytesIns_Inst_Sbox_0_T22), .B0_f (new_AGEMA_signal_6946), .B1_t (new_AGEMA_signal_6947), .B1_f (new_AGEMA_signal_6948), .Z0_t (SubBytesIns_Inst_Sbox_0_T23), .Z0_f (new_AGEMA_signal_7487), .Z1_t (new_AGEMA_signal_7488), .Z1_f (new_AGEMA_signal_7489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T2), .A0_f (new_AGEMA_signal_6349), .A1_t (new_AGEMA_signal_6350), .A1_f (new_AGEMA_signal_6351), .B0_t (SubBytesIns_Inst_Sbox_0_T10), .B0_f (new_AGEMA_signal_7475), .B1_t (new_AGEMA_signal_7476), .B1_f (new_AGEMA_signal_7477), .Z0_t (SubBytesIns_Inst_Sbox_0_T24), .Z0_f (new_AGEMA_signal_8204), .Z1_t (new_AGEMA_signal_8205), .Z1_f (new_AGEMA_signal_8206) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T20), .A0_f (new_AGEMA_signal_7484), .A1_t (new_AGEMA_signal_7485), .A1_f (new_AGEMA_signal_7486), .B0_t (SubBytesIns_Inst_Sbox_0_T17), .B0_f (new_AGEMA_signal_7481), .B1_t (new_AGEMA_signal_7482), .B1_f (new_AGEMA_signal_7483), .Z0_t (SubBytesIns_Inst_Sbox_0_T25), .Z0_f (new_AGEMA_signal_8207), .Z1_t (new_AGEMA_signal_8208), .Z1_f (new_AGEMA_signal_8209) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T3), .A0_f (new_AGEMA_signal_6352), .A1_t (new_AGEMA_signal_6353), .A1_f (new_AGEMA_signal_6354), .B0_t (SubBytesIns_Inst_Sbox_0_T16), .B0_f (new_AGEMA_signal_6940), .B1_t (new_AGEMA_signal_6941), .B1_f (new_AGEMA_signal_6942), .Z0_t (SubBytesIns_Inst_Sbox_0_T26), .Z0_f (new_AGEMA_signal_7490), .Z1_t (new_AGEMA_signal_7491), .Z1_f (new_AGEMA_signal_7492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T1), .A0_f (new_AGEMA_signal_6346), .A1_t (new_AGEMA_signal_6347), .A1_f (new_AGEMA_signal_6348), .B0_t (SubBytesIns_Inst_Sbox_0_T12), .B0_f (new_AGEMA_signal_6367), .B1_t (new_AGEMA_signal_6368), .B1_f (new_AGEMA_signal_6369), .Z0_t (SubBytesIns_Inst_Sbox_0_T27), .Z0_f (new_AGEMA_signal_6949), .Z1_t (new_AGEMA_signal_6950), .Z1_f (new_AGEMA_signal_6951) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T13), .A0_f (new_AGEMA_signal_6934), .A1_t (new_AGEMA_signal_6935), .A1_f (new_AGEMA_signal_6936), .B0_t (SubBytesIns_Inst_Sbox_0_T6), .B0_f (new_AGEMA_signal_6928), .B1_t (new_AGEMA_signal_6929), .B1_f (new_AGEMA_signal_6930), .Z0_t (SubBytesIns_Inst_Sbox_0_M1), .Z0_f (new_AGEMA_signal_7493), .Z1_t (new_AGEMA_signal_7494), .Z1_f (new_AGEMA_signal_7495) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T23), .A0_f (new_AGEMA_signal_7487), .A1_t (new_AGEMA_signal_7488), .A1_f (new_AGEMA_signal_7489), .B0_t (SubBytesIns_Inst_Sbox_0_T8), .B0_f (new_AGEMA_signal_7472), .B1_t (new_AGEMA_signal_7473), .B1_f (new_AGEMA_signal_7474), .Z0_t (SubBytesIns_Inst_Sbox_0_M2), .Z0_f (new_AGEMA_signal_8210), .Z1_t (new_AGEMA_signal_8211), .Z1_f (new_AGEMA_signal_8212) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T14), .A0_f (new_AGEMA_signal_7478), .A1_t (new_AGEMA_signal_7479), .A1_f (new_AGEMA_signal_7480), .B0_t (SubBytesIns_Inst_Sbox_0_M1), .B0_f (new_AGEMA_signal_7493), .B1_t (new_AGEMA_signal_7494), .B1_f (new_AGEMA_signal_7495), .Z0_t (SubBytesIns_Inst_Sbox_0_M3), .Z0_f (new_AGEMA_signal_8213), .Z1_t (new_AGEMA_signal_8214), .Z1_f (new_AGEMA_signal_8215) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T19), .A0_f (new_AGEMA_signal_6943), .A1_t (new_AGEMA_signal_6944), .A1_f (new_AGEMA_signal_6945), .B0_t (ciphertext_s0_t[0]), .B0_f (ciphertext_s0_f[0]), .B1_t (ciphertext_s1_t[0]), .B1_f (ciphertext_s1_f[0]), .Z0_t (SubBytesIns_Inst_Sbox_0_M4), .Z0_f (new_AGEMA_signal_7496), .Z1_t (new_AGEMA_signal_7497), .Z1_f (new_AGEMA_signal_7498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M4), .A0_f (new_AGEMA_signal_7496), .A1_t (new_AGEMA_signal_7497), .A1_f (new_AGEMA_signal_7498), .B0_t (SubBytesIns_Inst_Sbox_0_M1), .B0_f (new_AGEMA_signal_7493), .B1_t (new_AGEMA_signal_7494), .B1_f (new_AGEMA_signal_7495), .Z0_t (SubBytesIns_Inst_Sbox_0_M5), .Z0_f (new_AGEMA_signal_8216), .Z1_t (new_AGEMA_signal_8217), .Z1_f (new_AGEMA_signal_8218) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T3), .A0_f (new_AGEMA_signal_6352), .A1_t (new_AGEMA_signal_6353), .A1_f (new_AGEMA_signal_6354), .B0_t (SubBytesIns_Inst_Sbox_0_T16), .B0_f (new_AGEMA_signal_6940), .B1_t (new_AGEMA_signal_6941), .B1_f (new_AGEMA_signal_6942), .Z0_t (SubBytesIns_Inst_Sbox_0_M6), .Z0_f (new_AGEMA_signal_7499), .Z1_t (new_AGEMA_signal_7500), .Z1_f (new_AGEMA_signal_7501) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T22), .A0_f (new_AGEMA_signal_6946), .A1_t (new_AGEMA_signal_6947), .A1_f (new_AGEMA_signal_6948), .B0_t (SubBytesIns_Inst_Sbox_0_T9), .B0_f (new_AGEMA_signal_6931), .B1_t (new_AGEMA_signal_6932), .B1_f (new_AGEMA_signal_6933), .Z0_t (SubBytesIns_Inst_Sbox_0_M7), .Z0_f (new_AGEMA_signal_7502), .Z1_t (new_AGEMA_signal_7503), .Z1_f (new_AGEMA_signal_7504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T26), .A0_f (new_AGEMA_signal_7490), .A1_t (new_AGEMA_signal_7491), .A1_f (new_AGEMA_signal_7492), .B0_t (SubBytesIns_Inst_Sbox_0_M6), .B0_f (new_AGEMA_signal_7499), .B1_t (new_AGEMA_signal_7500), .B1_f (new_AGEMA_signal_7501), .Z0_t (SubBytesIns_Inst_Sbox_0_M8), .Z0_f (new_AGEMA_signal_8219), .Z1_t (new_AGEMA_signal_8220), .Z1_f (new_AGEMA_signal_8221) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T20), .A0_f (new_AGEMA_signal_7484), .A1_t (new_AGEMA_signal_7485), .A1_f (new_AGEMA_signal_7486), .B0_t (SubBytesIns_Inst_Sbox_0_T17), .B0_f (new_AGEMA_signal_7481), .B1_t (new_AGEMA_signal_7482), .B1_f (new_AGEMA_signal_7483), .Z0_t (SubBytesIns_Inst_Sbox_0_M9), .Z0_f (new_AGEMA_signal_8222), .Z1_t (new_AGEMA_signal_8223), .Z1_f (new_AGEMA_signal_8224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M9), .A0_f (new_AGEMA_signal_8222), .A1_t (new_AGEMA_signal_8223), .A1_f (new_AGEMA_signal_8224), .B0_t (SubBytesIns_Inst_Sbox_0_M6), .B0_f (new_AGEMA_signal_7499), .B1_t (new_AGEMA_signal_7500), .B1_f (new_AGEMA_signal_7501), .Z0_t (SubBytesIns_Inst_Sbox_0_M10), .Z0_f (new_AGEMA_signal_8696), .Z1_t (new_AGEMA_signal_8697), .Z1_f (new_AGEMA_signal_8698) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T1), .A0_f (new_AGEMA_signal_6346), .A1_t (new_AGEMA_signal_6347), .A1_f (new_AGEMA_signal_6348), .B0_t (SubBytesIns_Inst_Sbox_0_T15), .B0_f (new_AGEMA_signal_6937), .B1_t (new_AGEMA_signal_6938), .B1_f (new_AGEMA_signal_6939), .Z0_t (SubBytesIns_Inst_Sbox_0_M11), .Z0_f (new_AGEMA_signal_7505), .Z1_t (new_AGEMA_signal_7506), .Z1_f (new_AGEMA_signal_7507) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T4), .A0_f (new_AGEMA_signal_6355), .A1_t (new_AGEMA_signal_6356), .A1_f (new_AGEMA_signal_6357), .B0_t (SubBytesIns_Inst_Sbox_0_T27), .B0_f (new_AGEMA_signal_6949), .B1_t (new_AGEMA_signal_6950), .B1_f (new_AGEMA_signal_6951), .Z0_t (SubBytesIns_Inst_Sbox_0_M12), .Z0_f (new_AGEMA_signal_7508), .Z1_t (new_AGEMA_signal_7509), .Z1_f (new_AGEMA_signal_7510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M12), .A0_f (new_AGEMA_signal_7508), .A1_t (new_AGEMA_signal_7509), .A1_f (new_AGEMA_signal_7510), .B0_t (SubBytesIns_Inst_Sbox_0_M11), .B0_f (new_AGEMA_signal_7505), .B1_t (new_AGEMA_signal_7506), .B1_f (new_AGEMA_signal_7507), .Z0_t (SubBytesIns_Inst_Sbox_0_M13), .Z0_f (new_AGEMA_signal_8225), .Z1_t (new_AGEMA_signal_8226), .Z1_f (new_AGEMA_signal_8227) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T2), .A0_f (new_AGEMA_signal_6349), .A1_t (new_AGEMA_signal_6350), .A1_f (new_AGEMA_signal_6351), .B0_t (SubBytesIns_Inst_Sbox_0_T10), .B0_f (new_AGEMA_signal_7475), .B1_t (new_AGEMA_signal_7476), .B1_f (new_AGEMA_signal_7477), .Z0_t (SubBytesIns_Inst_Sbox_0_M14), .Z0_f (new_AGEMA_signal_8228), .Z1_t (new_AGEMA_signal_8229), .Z1_f (new_AGEMA_signal_8230) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M14), .A0_f (new_AGEMA_signal_8228), .A1_t (new_AGEMA_signal_8229), .A1_f (new_AGEMA_signal_8230), .B0_t (SubBytesIns_Inst_Sbox_0_M11), .B0_f (new_AGEMA_signal_7505), .B1_t (new_AGEMA_signal_7506), .B1_f (new_AGEMA_signal_7507), .Z0_t (SubBytesIns_Inst_Sbox_0_M15), .Z0_f (new_AGEMA_signal_8699), .Z1_t (new_AGEMA_signal_8700), .Z1_f (new_AGEMA_signal_8701) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M3), .A0_f (new_AGEMA_signal_8213), .A1_t (new_AGEMA_signal_8214), .A1_f (new_AGEMA_signal_8215), .B0_t (SubBytesIns_Inst_Sbox_0_M2), .B0_f (new_AGEMA_signal_8210), .B1_t (new_AGEMA_signal_8211), .B1_f (new_AGEMA_signal_8212), .Z0_t (SubBytesIns_Inst_Sbox_0_M16), .Z0_f (new_AGEMA_signal_8702), .Z1_t (new_AGEMA_signal_8703), .Z1_f (new_AGEMA_signal_8704) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M5), .A0_f (new_AGEMA_signal_8216), .A1_t (new_AGEMA_signal_8217), .A1_f (new_AGEMA_signal_8218), .B0_t (SubBytesIns_Inst_Sbox_0_T24), .B0_f (new_AGEMA_signal_8204), .B1_t (new_AGEMA_signal_8205), .B1_f (new_AGEMA_signal_8206), .Z0_t (SubBytesIns_Inst_Sbox_0_M17), .Z0_f (new_AGEMA_signal_8705), .Z1_t (new_AGEMA_signal_8706), .Z1_f (new_AGEMA_signal_8707) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M8), .A0_f (new_AGEMA_signal_8219), .A1_t (new_AGEMA_signal_8220), .A1_f (new_AGEMA_signal_8221), .B0_t (SubBytesIns_Inst_Sbox_0_M7), .B0_f (new_AGEMA_signal_7502), .B1_t (new_AGEMA_signal_7503), .B1_f (new_AGEMA_signal_7504), .Z0_t (SubBytesIns_Inst_Sbox_0_M18), .Z0_f (new_AGEMA_signal_8708), .Z1_t (new_AGEMA_signal_8709), .Z1_f (new_AGEMA_signal_8710) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M10), .A0_f (new_AGEMA_signal_8696), .A1_t (new_AGEMA_signal_8697), .A1_f (new_AGEMA_signal_8698), .B0_t (SubBytesIns_Inst_Sbox_0_M15), .B0_f (new_AGEMA_signal_8699), .B1_t (new_AGEMA_signal_8700), .B1_f (new_AGEMA_signal_8701), .Z0_t (SubBytesIns_Inst_Sbox_0_M19), .Z0_f (new_AGEMA_signal_8984), .Z1_t (new_AGEMA_signal_8985), .Z1_f (new_AGEMA_signal_8986) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M16), .A0_f (new_AGEMA_signal_8702), .A1_t (new_AGEMA_signal_8703), .A1_f (new_AGEMA_signal_8704), .B0_t (SubBytesIns_Inst_Sbox_0_M13), .B0_f (new_AGEMA_signal_8225), .B1_t (new_AGEMA_signal_8226), .B1_f (new_AGEMA_signal_8227), .Z0_t (SubBytesIns_Inst_Sbox_0_M20), .Z0_f (new_AGEMA_signal_8987), .Z1_t (new_AGEMA_signal_8988), .Z1_f (new_AGEMA_signal_8989) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M17), .A0_f (new_AGEMA_signal_8705), .A1_t (new_AGEMA_signal_8706), .A1_f (new_AGEMA_signal_8707), .B0_t (SubBytesIns_Inst_Sbox_0_M15), .B0_f (new_AGEMA_signal_8699), .B1_t (new_AGEMA_signal_8700), .B1_f (new_AGEMA_signal_8701), .Z0_t (SubBytesIns_Inst_Sbox_0_M21), .Z0_f (new_AGEMA_signal_8990), .Z1_t (new_AGEMA_signal_8991), .Z1_f (new_AGEMA_signal_8992) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M18), .A0_f (new_AGEMA_signal_8708), .A1_t (new_AGEMA_signal_8709), .A1_f (new_AGEMA_signal_8710), .B0_t (SubBytesIns_Inst_Sbox_0_M13), .B0_f (new_AGEMA_signal_8225), .B1_t (new_AGEMA_signal_8226), .B1_f (new_AGEMA_signal_8227), .Z0_t (SubBytesIns_Inst_Sbox_0_M22), .Z0_f (new_AGEMA_signal_8993), .Z1_t (new_AGEMA_signal_8994), .Z1_f (new_AGEMA_signal_8995) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M19), .A0_f (new_AGEMA_signal_8984), .A1_t (new_AGEMA_signal_8985), .A1_f (new_AGEMA_signal_8986), .B0_t (SubBytesIns_Inst_Sbox_0_T25), .B0_f (new_AGEMA_signal_8207), .B1_t (new_AGEMA_signal_8208), .B1_f (new_AGEMA_signal_8209), .Z0_t (SubBytesIns_Inst_Sbox_0_M23), .Z0_f (new_AGEMA_signal_9224), .Z1_t (new_AGEMA_signal_9225), .Z1_f (new_AGEMA_signal_9226) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M22), .A0_f (new_AGEMA_signal_8993), .A1_t (new_AGEMA_signal_8994), .A1_f (new_AGEMA_signal_8995), .B0_t (SubBytesIns_Inst_Sbox_0_M23), .B0_f (new_AGEMA_signal_9224), .B1_t (new_AGEMA_signal_9225), .B1_f (new_AGEMA_signal_9226), .Z0_t (SubBytesIns_Inst_Sbox_0_M24), .Z0_f (new_AGEMA_signal_9476), .Z1_t (new_AGEMA_signal_9477), .Z1_f (new_AGEMA_signal_9478) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M22), .A0_f (new_AGEMA_signal_8993), .A1_t (new_AGEMA_signal_8994), .A1_f (new_AGEMA_signal_8995), .B0_t (SubBytesIns_Inst_Sbox_0_M20), .B0_f (new_AGEMA_signal_8987), .B1_t (new_AGEMA_signal_8988), .B1_f (new_AGEMA_signal_8989), .Z0_t (SubBytesIns_Inst_Sbox_0_M25), .Z0_f (new_AGEMA_signal_9227), .Z1_t (new_AGEMA_signal_9228), .Z1_f (new_AGEMA_signal_9229) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M21), .A0_f (new_AGEMA_signal_8990), .A1_t (new_AGEMA_signal_8991), .A1_f (new_AGEMA_signal_8992), .B0_t (SubBytesIns_Inst_Sbox_0_M25), .B0_f (new_AGEMA_signal_9227), .B1_t (new_AGEMA_signal_9228), .B1_f (new_AGEMA_signal_9229), .Z0_t (SubBytesIns_Inst_Sbox_0_M26), .Z0_f (new_AGEMA_signal_9479), .Z1_t (new_AGEMA_signal_9480), .Z1_f (new_AGEMA_signal_9481) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M20), .A0_f (new_AGEMA_signal_8987), .A1_t (new_AGEMA_signal_8988), .A1_f (new_AGEMA_signal_8989), .B0_t (SubBytesIns_Inst_Sbox_0_M21), .B0_f (new_AGEMA_signal_8990), .B1_t (new_AGEMA_signal_8991), .B1_f (new_AGEMA_signal_8992), .Z0_t (SubBytesIns_Inst_Sbox_0_M27), .Z0_f (new_AGEMA_signal_9230), .Z1_t (new_AGEMA_signal_9231), .Z1_f (new_AGEMA_signal_9232) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M23), .A0_f (new_AGEMA_signal_9224), .A1_t (new_AGEMA_signal_9225), .A1_f (new_AGEMA_signal_9226), .B0_t (SubBytesIns_Inst_Sbox_0_M25), .B0_f (new_AGEMA_signal_9227), .B1_t (new_AGEMA_signal_9228), .B1_f (new_AGEMA_signal_9229), .Z0_t (SubBytesIns_Inst_Sbox_0_M28), .Z0_f (new_AGEMA_signal_9482), .Z1_t (new_AGEMA_signal_9483), .Z1_f (new_AGEMA_signal_9484) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M28), .A0_f (new_AGEMA_signal_9482), .A1_t (new_AGEMA_signal_9483), .A1_f (new_AGEMA_signal_9484), .B0_t (SubBytesIns_Inst_Sbox_0_M27), .B0_f (new_AGEMA_signal_9230), .B1_t (new_AGEMA_signal_9231), .B1_f (new_AGEMA_signal_9232), .Z0_t (SubBytesIns_Inst_Sbox_0_M29), .Z0_f (new_AGEMA_signal_9776), .Z1_t (new_AGEMA_signal_9777), .Z1_f (new_AGEMA_signal_9778) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M26), .A0_f (new_AGEMA_signal_9479), .A1_t (new_AGEMA_signal_9480), .A1_f (new_AGEMA_signal_9481), .B0_t (SubBytesIns_Inst_Sbox_0_M24), .B0_f (new_AGEMA_signal_9476), .B1_t (new_AGEMA_signal_9477), .B1_f (new_AGEMA_signal_9478), .Z0_t (SubBytesIns_Inst_Sbox_0_M30), .Z0_f (new_AGEMA_signal_9779), .Z1_t (new_AGEMA_signal_9780), .Z1_f (new_AGEMA_signal_9781) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M20), .A0_f (new_AGEMA_signal_8987), .A1_t (new_AGEMA_signal_8988), .A1_f (new_AGEMA_signal_8989), .B0_t (SubBytesIns_Inst_Sbox_0_M23), .B0_f (new_AGEMA_signal_9224), .B1_t (new_AGEMA_signal_9225), .B1_f (new_AGEMA_signal_9226), .Z0_t (SubBytesIns_Inst_Sbox_0_M31), .Z0_f (new_AGEMA_signal_9485), .Z1_t (new_AGEMA_signal_9486), .Z1_f (new_AGEMA_signal_9487) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M27), .A0_f (new_AGEMA_signal_9230), .A1_t (new_AGEMA_signal_9231), .A1_f (new_AGEMA_signal_9232), .B0_t (SubBytesIns_Inst_Sbox_0_M31), .B0_f (new_AGEMA_signal_9485), .B1_t (new_AGEMA_signal_9486), .B1_f (new_AGEMA_signal_9487), .Z0_t (SubBytesIns_Inst_Sbox_0_M32), .Z0_f (new_AGEMA_signal_9782), .Z1_t (new_AGEMA_signal_9783), .Z1_f (new_AGEMA_signal_9784) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M27), .A0_f (new_AGEMA_signal_9230), .A1_t (new_AGEMA_signal_9231), .A1_f (new_AGEMA_signal_9232), .B0_t (SubBytesIns_Inst_Sbox_0_M25), .B0_f (new_AGEMA_signal_9227), .B1_t (new_AGEMA_signal_9228), .B1_f (new_AGEMA_signal_9229), .Z0_t (SubBytesIns_Inst_Sbox_0_M33), .Z0_f (new_AGEMA_signal_9488), .Z1_t (new_AGEMA_signal_9489), .Z1_f (new_AGEMA_signal_9490) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M21), .A0_f (new_AGEMA_signal_8990), .A1_t (new_AGEMA_signal_8991), .A1_f (new_AGEMA_signal_8992), .B0_t (SubBytesIns_Inst_Sbox_0_M22), .B0_f (new_AGEMA_signal_8993), .B1_t (new_AGEMA_signal_8994), .B1_f (new_AGEMA_signal_8995), .Z0_t (SubBytesIns_Inst_Sbox_0_M34), .Z0_f (new_AGEMA_signal_9233), .Z1_t (new_AGEMA_signal_9234), .Z1_f (new_AGEMA_signal_9235) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M24), .A0_f (new_AGEMA_signal_9476), .A1_t (new_AGEMA_signal_9477), .A1_f (new_AGEMA_signal_9478), .B0_t (SubBytesIns_Inst_Sbox_0_M34), .B0_f (new_AGEMA_signal_9233), .B1_t (new_AGEMA_signal_9234), .B1_f (new_AGEMA_signal_9235), .Z0_t (SubBytesIns_Inst_Sbox_0_M35), .Z0_f (new_AGEMA_signal_9785), .Z1_t (new_AGEMA_signal_9786), .Z1_f (new_AGEMA_signal_9787) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M24), .A0_f (new_AGEMA_signal_9476), .A1_t (new_AGEMA_signal_9477), .A1_f (new_AGEMA_signal_9478), .B0_t (SubBytesIns_Inst_Sbox_0_M25), .B0_f (new_AGEMA_signal_9227), .B1_t (new_AGEMA_signal_9228), .B1_f (new_AGEMA_signal_9229), .Z0_t (SubBytesIns_Inst_Sbox_0_M36), .Z0_f (new_AGEMA_signal_9788), .Z1_t (new_AGEMA_signal_9789), .Z1_f (new_AGEMA_signal_9790) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M21), .A0_f (new_AGEMA_signal_8990), .A1_t (new_AGEMA_signal_8991), .A1_f (new_AGEMA_signal_8992), .B0_t (SubBytesIns_Inst_Sbox_0_M29), .B0_f (new_AGEMA_signal_9776), .B1_t (new_AGEMA_signal_9777), .B1_f (new_AGEMA_signal_9778), .Z0_t (SubBytesIns_Inst_Sbox_0_M37), .Z0_f (new_AGEMA_signal_10064), .Z1_t (new_AGEMA_signal_10065), .Z1_f (new_AGEMA_signal_10066) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M32), .A0_f (new_AGEMA_signal_9782), .A1_t (new_AGEMA_signal_9783), .A1_f (new_AGEMA_signal_9784), .B0_t (SubBytesIns_Inst_Sbox_0_M33), .B0_f (new_AGEMA_signal_9488), .B1_t (new_AGEMA_signal_9489), .B1_f (new_AGEMA_signal_9490), .Z0_t (SubBytesIns_Inst_Sbox_0_M38), .Z0_f (new_AGEMA_signal_10067), .Z1_t (new_AGEMA_signal_10068), .Z1_f (new_AGEMA_signal_10069) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M23), .A0_f (new_AGEMA_signal_9224), .A1_t (new_AGEMA_signal_9225), .A1_f (new_AGEMA_signal_9226), .B0_t (SubBytesIns_Inst_Sbox_0_M30), .B0_f (new_AGEMA_signal_9779), .B1_t (new_AGEMA_signal_9780), .B1_f (new_AGEMA_signal_9781), .Z0_t (SubBytesIns_Inst_Sbox_0_M39), .Z0_f (new_AGEMA_signal_10070), .Z1_t (new_AGEMA_signal_10071), .Z1_f (new_AGEMA_signal_10072) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M35), .A0_f (new_AGEMA_signal_9785), .A1_t (new_AGEMA_signal_9786), .A1_f (new_AGEMA_signal_9787), .B0_t (SubBytesIns_Inst_Sbox_0_M36), .B0_f (new_AGEMA_signal_9788), .B1_t (new_AGEMA_signal_9789), .B1_f (new_AGEMA_signal_9790), .Z0_t (SubBytesIns_Inst_Sbox_0_M40), .Z0_f (new_AGEMA_signal_10073), .Z1_t (new_AGEMA_signal_10074), .Z1_f (new_AGEMA_signal_10075) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M38), .A0_f (new_AGEMA_signal_10067), .A1_t (new_AGEMA_signal_10068), .A1_f (new_AGEMA_signal_10069), .B0_t (SubBytesIns_Inst_Sbox_0_M40), .B0_f (new_AGEMA_signal_10073), .B1_t (new_AGEMA_signal_10074), .B1_f (new_AGEMA_signal_10075), .Z0_t (SubBytesIns_Inst_Sbox_0_M41), .Z0_f (new_AGEMA_signal_10400), .Z1_t (new_AGEMA_signal_10401), .Z1_f (new_AGEMA_signal_10402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M37), .A0_f (new_AGEMA_signal_10064), .A1_t (new_AGEMA_signal_10065), .A1_f (new_AGEMA_signal_10066), .B0_t (SubBytesIns_Inst_Sbox_0_M39), .B0_f (new_AGEMA_signal_10070), .B1_t (new_AGEMA_signal_10071), .B1_f (new_AGEMA_signal_10072), .Z0_t (SubBytesIns_Inst_Sbox_0_M42), .Z0_f (new_AGEMA_signal_10403), .Z1_t (new_AGEMA_signal_10404), .Z1_f (new_AGEMA_signal_10405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M37), .A0_f (new_AGEMA_signal_10064), .A1_t (new_AGEMA_signal_10065), .A1_f (new_AGEMA_signal_10066), .B0_t (SubBytesIns_Inst_Sbox_0_M38), .B0_f (new_AGEMA_signal_10067), .B1_t (new_AGEMA_signal_10068), .B1_f (new_AGEMA_signal_10069), .Z0_t (SubBytesIns_Inst_Sbox_0_M43), .Z0_f (new_AGEMA_signal_10406), .Z1_t (new_AGEMA_signal_10407), .Z1_f (new_AGEMA_signal_10408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M39), .A0_f (new_AGEMA_signal_10070), .A1_t (new_AGEMA_signal_10071), .A1_f (new_AGEMA_signal_10072), .B0_t (SubBytesIns_Inst_Sbox_0_M40), .B0_f (new_AGEMA_signal_10073), .B1_t (new_AGEMA_signal_10074), .B1_f (new_AGEMA_signal_10075), .Z0_t (SubBytesIns_Inst_Sbox_0_M44), .Z0_f (new_AGEMA_signal_10409), .Z1_t (new_AGEMA_signal_10410), .Z1_f (new_AGEMA_signal_10411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M42), .A0_f (new_AGEMA_signal_10403), .A1_t (new_AGEMA_signal_10404), .A1_f (new_AGEMA_signal_10405), .B0_t (SubBytesIns_Inst_Sbox_0_M41), .B0_f (new_AGEMA_signal_10400), .B1_t (new_AGEMA_signal_10401), .B1_f (new_AGEMA_signal_10402), .Z0_t (SubBytesIns_Inst_Sbox_0_M45), .Z0_f (new_AGEMA_signal_11120), .Z1_t (new_AGEMA_signal_11121), .Z1_f (new_AGEMA_signal_11122) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M44), .A0_f (new_AGEMA_signal_10409), .A1_t (new_AGEMA_signal_10410), .A1_f (new_AGEMA_signal_10411), .B0_t (SubBytesIns_Inst_Sbox_0_T6), .B0_f (new_AGEMA_signal_6928), .B1_t (new_AGEMA_signal_6929), .B1_f (new_AGEMA_signal_6930), .Z0_t (SubBytesIns_Inst_Sbox_0_M46), .Z0_f (new_AGEMA_signal_11123), .Z1_t (new_AGEMA_signal_11124), .Z1_f (new_AGEMA_signal_11125) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M40), .A0_f (new_AGEMA_signal_10073), .A1_t (new_AGEMA_signal_10074), .A1_f (new_AGEMA_signal_10075), .B0_t (SubBytesIns_Inst_Sbox_0_T8), .B0_f (new_AGEMA_signal_7472), .B1_t (new_AGEMA_signal_7473), .B1_f (new_AGEMA_signal_7474), .Z0_t (SubBytesIns_Inst_Sbox_0_M47), .Z0_f (new_AGEMA_signal_10412), .Z1_t (new_AGEMA_signal_10413), .Z1_f (new_AGEMA_signal_10414) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M39), .A0_f (new_AGEMA_signal_10070), .A1_t (new_AGEMA_signal_10071), .A1_f (new_AGEMA_signal_10072), .B0_t (ciphertext_s0_t[0]), .B0_f (ciphertext_s0_f[0]), .B1_t (ciphertext_s1_t[0]), .B1_f (ciphertext_s1_f[0]), .Z0_t (SubBytesIns_Inst_Sbox_0_M48), .Z0_f (new_AGEMA_signal_10415), .Z1_t (new_AGEMA_signal_10416), .Z1_f (new_AGEMA_signal_10417) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M43), .A0_f (new_AGEMA_signal_10406), .A1_t (new_AGEMA_signal_10407), .A1_f (new_AGEMA_signal_10408), .B0_t (SubBytesIns_Inst_Sbox_0_T16), .B0_f (new_AGEMA_signal_6940), .B1_t (new_AGEMA_signal_6941), .B1_f (new_AGEMA_signal_6942), .Z0_t (SubBytesIns_Inst_Sbox_0_M49), .Z0_f (new_AGEMA_signal_11126), .Z1_t (new_AGEMA_signal_11127), .Z1_f (new_AGEMA_signal_11128) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M38), .A0_f (new_AGEMA_signal_10067), .A1_t (new_AGEMA_signal_10068), .A1_f (new_AGEMA_signal_10069), .B0_t (SubBytesIns_Inst_Sbox_0_T9), .B0_f (new_AGEMA_signal_6931), .B1_t (new_AGEMA_signal_6932), .B1_f (new_AGEMA_signal_6933), .Z0_t (SubBytesIns_Inst_Sbox_0_M50), .Z0_f (new_AGEMA_signal_10418), .Z1_t (new_AGEMA_signal_10419), .Z1_f (new_AGEMA_signal_10420) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M37), .A0_f (new_AGEMA_signal_10064), .A1_t (new_AGEMA_signal_10065), .A1_f (new_AGEMA_signal_10066), .B0_t (SubBytesIns_Inst_Sbox_0_T17), .B0_f (new_AGEMA_signal_7481), .B1_t (new_AGEMA_signal_7482), .B1_f (new_AGEMA_signal_7483), .Z0_t (SubBytesIns_Inst_Sbox_0_M51), .Z0_f (new_AGEMA_signal_10421), .Z1_t (new_AGEMA_signal_10422), .Z1_f (new_AGEMA_signal_10423) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M42), .A0_f (new_AGEMA_signal_10403), .A1_t (new_AGEMA_signal_10404), .A1_f (new_AGEMA_signal_10405), .B0_t (SubBytesIns_Inst_Sbox_0_T15), .B0_f (new_AGEMA_signal_6937), .B1_t (new_AGEMA_signal_6938), .B1_f (new_AGEMA_signal_6939), .Z0_t (SubBytesIns_Inst_Sbox_0_M52), .Z0_f (new_AGEMA_signal_11129), .Z1_t (new_AGEMA_signal_11130), .Z1_f (new_AGEMA_signal_11131) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M45), .A0_f (new_AGEMA_signal_11120), .A1_t (new_AGEMA_signal_11121), .A1_f (new_AGEMA_signal_11122), .B0_t (SubBytesIns_Inst_Sbox_0_T27), .B0_f (new_AGEMA_signal_6949), .B1_t (new_AGEMA_signal_6950), .B1_f (new_AGEMA_signal_6951), .Z0_t (SubBytesIns_Inst_Sbox_0_M53), .Z0_f (new_AGEMA_signal_11816), .Z1_t (new_AGEMA_signal_11817), .Z1_f (new_AGEMA_signal_11818) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M41), .A0_f (new_AGEMA_signal_10400), .A1_t (new_AGEMA_signal_10401), .A1_f (new_AGEMA_signal_10402), .B0_t (SubBytesIns_Inst_Sbox_0_T10), .B0_f (new_AGEMA_signal_7475), .B1_t (new_AGEMA_signal_7476), .B1_f (new_AGEMA_signal_7477), .Z0_t (SubBytesIns_Inst_Sbox_0_M54), .Z0_f (new_AGEMA_signal_11132), .Z1_t (new_AGEMA_signal_11133), .Z1_f (new_AGEMA_signal_11134) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M44), .A0_f (new_AGEMA_signal_10409), .A1_t (new_AGEMA_signal_10410), .A1_f (new_AGEMA_signal_10411), .B0_t (SubBytesIns_Inst_Sbox_0_T13), .B0_f (new_AGEMA_signal_6934), .B1_t (new_AGEMA_signal_6935), .B1_f (new_AGEMA_signal_6936), .Z0_t (SubBytesIns_Inst_Sbox_0_M55), .Z0_f (new_AGEMA_signal_11135), .Z1_t (new_AGEMA_signal_11136), .Z1_f (new_AGEMA_signal_11137) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M40), .A0_f (new_AGEMA_signal_10073), .A1_t (new_AGEMA_signal_10074), .A1_f (new_AGEMA_signal_10075), .B0_t (SubBytesIns_Inst_Sbox_0_T23), .B0_f (new_AGEMA_signal_7487), .B1_t (new_AGEMA_signal_7488), .B1_f (new_AGEMA_signal_7489), .Z0_t (SubBytesIns_Inst_Sbox_0_M56), .Z0_f (new_AGEMA_signal_10424), .Z1_t (new_AGEMA_signal_10425), .Z1_f (new_AGEMA_signal_10426) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M39), .A0_f (new_AGEMA_signal_10070), .A1_t (new_AGEMA_signal_10071), .A1_f (new_AGEMA_signal_10072), .B0_t (SubBytesIns_Inst_Sbox_0_T19), .B0_f (new_AGEMA_signal_6943), .B1_t (new_AGEMA_signal_6944), .B1_f (new_AGEMA_signal_6945), .Z0_t (SubBytesIns_Inst_Sbox_0_M57), .Z0_f (new_AGEMA_signal_10427), .Z1_t (new_AGEMA_signal_10428), .Z1_f (new_AGEMA_signal_10429) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M43), .A0_f (new_AGEMA_signal_10406), .A1_t (new_AGEMA_signal_10407), .A1_f (new_AGEMA_signal_10408), .B0_t (SubBytesIns_Inst_Sbox_0_T3), .B0_f (new_AGEMA_signal_6352), .B1_t (new_AGEMA_signal_6353), .B1_f (new_AGEMA_signal_6354), .Z0_t (SubBytesIns_Inst_Sbox_0_M58), .Z0_f (new_AGEMA_signal_11138), .Z1_t (new_AGEMA_signal_11139), .Z1_f (new_AGEMA_signal_11140) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M38), .A0_f (new_AGEMA_signal_10067), .A1_t (new_AGEMA_signal_10068), .A1_f (new_AGEMA_signal_10069), .B0_t (SubBytesIns_Inst_Sbox_0_T22), .B0_f (new_AGEMA_signal_6946), .B1_t (new_AGEMA_signal_6947), .B1_f (new_AGEMA_signal_6948), .Z0_t (SubBytesIns_Inst_Sbox_0_M59), .Z0_f (new_AGEMA_signal_10430), .Z1_t (new_AGEMA_signal_10431), .Z1_f (new_AGEMA_signal_10432) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M37), .A0_f (new_AGEMA_signal_10064), .A1_t (new_AGEMA_signal_10065), .A1_f (new_AGEMA_signal_10066), .B0_t (SubBytesIns_Inst_Sbox_0_T20), .B0_f (new_AGEMA_signal_7484), .B1_t (new_AGEMA_signal_7485), .B1_f (new_AGEMA_signal_7486), .Z0_t (SubBytesIns_Inst_Sbox_0_M60), .Z0_f (new_AGEMA_signal_10433), .Z1_t (new_AGEMA_signal_10434), .Z1_f (new_AGEMA_signal_10435) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M42), .A0_f (new_AGEMA_signal_10403), .A1_t (new_AGEMA_signal_10404), .A1_f (new_AGEMA_signal_10405), .B0_t (SubBytesIns_Inst_Sbox_0_T1), .B0_f (new_AGEMA_signal_6346), .B1_t (new_AGEMA_signal_6347), .B1_f (new_AGEMA_signal_6348), .Z0_t (SubBytesIns_Inst_Sbox_0_M61), .Z0_f (new_AGEMA_signal_11141), .Z1_t (new_AGEMA_signal_11142), .Z1_f (new_AGEMA_signal_11143) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M45), .A0_f (new_AGEMA_signal_11120), .A1_t (new_AGEMA_signal_11121), .A1_f (new_AGEMA_signal_11122), .B0_t (SubBytesIns_Inst_Sbox_0_T4), .B0_f (new_AGEMA_signal_6355), .B1_t (new_AGEMA_signal_6356), .B1_f (new_AGEMA_signal_6357), .Z0_t (SubBytesIns_Inst_Sbox_0_M62), .Z0_f (new_AGEMA_signal_11819), .Z1_t (new_AGEMA_signal_11820), .Z1_f (new_AGEMA_signal_11821) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M41), .A0_f (new_AGEMA_signal_10400), .A1_t (new_AGEMA_signal_10401), .A1_f (new_AGEMA_signal_10402), .B0_t (SubBytesIns_Inst_Sbox_0_T2), .B0_f (new_AGEMA_signal_6349), .B1_t (new_AGEMA_signal_6350), .B1_f (new_AGEMA_signal_6351), .Z0_t (SubBytesIns_Inst_Sbox_0_M63), .Z0_f (new_AGEMA_signal_11144), .Z1_t (new_AGEMA_signal_11145), .Z1_f (new_AGEMA_signal_11146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M61), .A0_f (new_AGEMA_signal_11141), .A1_t (new_AGEMA_signal_11142), .A1_f (new_AGEMA_signal_11143), .B0_t (SubBytesIns_Inst_Sbox_0_M62), .B0_f (new_AGEMA_signal_11819), .B1_t (new_AGEMA_signal_11820), .B1_f (new_AGEMA_signal_11821), .Z0_t (SubBytesIns_Inst_Sbox_0_L0), .Z0_f (new_AGEMA_signal_12404), .Z1_t (new_AGEMA_signal_12405), .Z1_f (new_AGEMA_signal_12406) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M50), .A0_f (new_AGEMA_signal_10418), .A1_t (new_AGEMA_signal_10419), .A1_f (new_AGEMA_signal_10420), .B0_t (SubBytesIns_Inst_Sbox_0_M56), .B0_f (new_AGEMA_signal_10424), .B1_t (new_AGEMA_signal_10425), .B1_f (new_AGEMA_signal_10426), .Z0_t (SubBytesIns_Inst_Sbox_0_L1), .Z0_f (new_AGEMA_signal_11147), .Z1_t (new_AGEMA_signal_11148), .Z1_f (new_AGEMA_signal_11149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M46), .A0_f (new_AGEMA_signal_11123), .A1_t (new_AGEMA_signal_11124), .A1_f (new_AGEMA_signal_11125), .B0_t (SubBytesIns_Inst_Sbox_0_M48), .B0_f (new_AGEMA_signal_10415), .B1_t (new_AGEMA_signal_10416), .B1_f (new_AGEMA_signal_10417), .Z0_t (SubBytesIns_Inst_Sbox_0_L2), .Z0_f (new_AGEMA_signal_11822), .Z1_t (new_AGEMA_signal_11823), .Z1_f (new_AGEMA_signal_11824) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M47), .A0_f (new_AGEMA_signal_10412), .A1_t (new_AGEMA_signal_10413), .A1_f (new_AGEMA_signal_10414), .B0_t (SubBytesIns_Inst_Sbox_0_M55), .B0_f (new_AGEMA_signal_11135), .B1_t (new_AGEMA_signal_11136), .B1_f (new_AGEMA_signal_11137), .Z0_t (SubBytesIns_Inst_Sbox_0_L3), .Z0_f (new_AGEMA_signal_11825), .Z1_t (new_AGEMA_signal_11826), .Z1_f (new_AGEMA_signal_11827) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M54), .A0_f (new_AGEMA_signal_11132), .A1_t (new_AGEMA_signal_11133), .A1_f (new_AGEMA_signal_11134), .B0_t (SubBytesIns_Inst_Sbox_0_M58), .B0_f (new_AGEMA_signal_11138), .B1_t (new_AGEMA_signal_11139), .B1_f (new_AGEMA_signal_11140), .Z0_t (SubBytesIns_Inst_Sbox_0_L4), .Z0_f (new_AGEMA_signal_11828), .Z1_t (new_AGEMA_signal_11829), .Z1_f (new_AGEMA_signal_11830) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M49), .A0_f (new_AGEMA_signal_11126), .A1_t (new_AGEMA_signal_11127), .A1_f (new_AGEMA_signal_11128), .B0_t (SubBytesIns_Inst_Sbox_0_M61), .B0_f (new_AGEMA_signal_11141), .B1_t (new_AGEMA_signal_11142), .B1_f (new_AGEMA_signal_11143), .Z0_t (SubBytesIns_Inst_Sbox_0_L5), .Z0_f (new_AGEMA_signal_11831), .Z1_t (new_AGEMA_signal_11832), .Z1_f (new_AGEMA_signal_11833) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M62), .A0_f (new_AGEMA_signal_11819), .A1_t (new_AGEMA_signal_11820), .A1_f (new_AGEMA_signal_11821), .B0_t (SubBytesIns_Inst_Sbox_0_L5), .B0_f (new_AGEMA_signal_11831), .B1_t (new_AGEMA_signal_11832), .B1_f (new_AGEMA_signal_11833), .Z0_t (SubBytesIns_Inst_Sbox_0_L6), .Z0_f (new_AGEMA_signal_12407), .Z1_t (new_AGEMA_signal_12408), .Z1_f (new_AGEMA_signal_12409) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M46), .A0_f (new_AGEMA_signal_11123), .A1_t (new_AGEMA_signal_11124), .A1_f (new_AGEMA_signal_11125), .B0_t (SubBytesIns_Inst_Sbox_0_L3), .B0_f (new_AGEMA_signal_11825), .B1_t (new_AGEMA_signal_11826), .B1_f (new_AGEMA_signal_11827), .Z0_t (SubBytesIns_Inst_Sbox_0_L7), .Z0_f (new_AGEMA_signal_12410), .Z1_t (new_AGEMA_signal_12411), .Z1_f (new_AGEMA_signal_12412) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M51), .A0_f (new_AGEMA_signal_10421), .A1_t (new_AGEMA_signal_10422), .A1_f (new_AGEMA_signal_10423), .B0_t (SubBytesIns_Inst_Sbox_0_M59), .B0_f (new_AGEMA_signal_10430), .B1_t (new_AGEMA_signal_10431), .B1_f (new_AGEMA_signal_10432), .Z0_t (SubBytesIns_Inst_Sbox_0_L8), .Z0_f (new_AGEMA_signal_11150), .Z1_t (new_AGEMA_signal_11151), .Z1_f (new_AGEMA_signal_11152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M52), .A0_f (new_AGEMA_signal_11129), .A1_t (new_AGEMA_signal_11130), .A1_f (new_AGEMA_signal_11131), .B0_t (SubBytesIns_Inst_Sbox_0_M53), .B0_f (new_AGEMA_signal_11816), .B1_t (new_AGEMA_signal_11817), .B1_f (new_AGEMA_signal_11818), .Z0_t (SubBytesIns_Inst_Sbox_0_L9), .Z0_f (new_AGEMA_signal_12413), .Z1_t (new_AGEMA_signal_12414), .Z1_f (new_AGEMA_signal_12415) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M53), .A0_f (new_AGEMA_signal_11816), .A1_t (new_AGEMA_signal_11817), .A1_f (new_AGEMA_signal_11818), .B0_t (SubBytesIns_Inst_Sbox_0_L4), .B0_f (new_AGEMA_signal_11828), .B1_t (new_AGEMA_signal_11829), .B1_f (new_AGEMA_signal_11830), .Z0_t (SubBytesIns_Inst_Sbox_0_L10), .Z0_f (new_AGEMA_signal_12416), .Z1_t (new_AGEMA_signal_12417), .Z1_f (new_AGEMA_signal_12418) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M60), .A0_f (new_AGEMA_signal_10433), .A1_t (new_AGEMA_signal_10434), .A1_f (new_AGEMA_signal_10435), .B0_t (SubBytesIns_Inst_Sbox_0_L2), .B0_f (new_AGEMA_signal_11822), .B1_t (new_AGEMA_signal_11823), .B1_f (new_AGEMA_signal_11824), .Z0_t (SubBytesIns_Inst_Sbox_0_L11), .Z0_f (new_AGEMA_signal_12419), .Z1_t (new_AGEMA_signal_12420), .Z1_f (new_AGEMA_signal_12421) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M48), .A0_f (new_AGEMA_signal_10415), .A1_t (new_AGEMA_signal_10416), .A1_f (new_AGEMA_signal_10417), .B0_t (SubBytesIns_Inst_Sbox_0_M51), .B0_f (new_AGEMA_signal_10421), .B1_t (new_AGEMA_signal_10422), .B1_f (new_AGEMA_signal_10423), .Z0_t (SubBytesIns_Inst_Sbox_0_L12), .Z0_f (new_AGEMA_signal_11153), .Z1_t (new_AGEMA_signal_11154), .Z1_f (new_AGEMA_signal_11155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M50), .A0_f (new_AGEMA_signal_10418), .A1_t (new_AGEMA_signal_10419), .A1_f (new_AGEMA_signal_10420), .B0_t (SubBytesIns_Inst_Sbox_0_L0), .B0_f (new_AGEMA_signal_12404), .B1_t (new_AGEMA_signal_12405), .B1_f (new_AGEMA_signal_12406), .Z0_t (SubBytesIns_Inst_Sbox_0_L13), .Z0_f (new_AGEMA_signal_12968), .Z1_t (new_AGEMA_signal_12969), .Z1_f (new_AGEMA_signal_12970) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M52), .A0_f (new_AGEMA_signal_11129), .A1_t (new_AGEMA_signal_11130), .A1_f (new_AGEMA_signal_11131), .B0_t (SubBytesIns_Inst_Sbox_0_M61), .B0_f (new_AGEMA_signal_11141), .B1_t (new_AGEMA_signal_11142), .B1_f (new_AGEMA_signal_11143), .Z0_t (SubBytesIns_Inst_Sbox_0_L14), .Z0_f (new_AGEMA_signal_11834), .Z1_t (new_AGEMA_signal_11835), .Z1_f (new_AGEMA_signal_11836) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M55), .A0_f (new_AGEMA_signal_11135), .A1_t (new_AGEMA_signal_11136), .A1_f (new_AGEMA_signal_11137), .B0_t (SubBytesIns_Inst_Sbox_0_L1), .B0_f (new_AGEMA_signal_11147), .B1_t (new_AGEMA_signal_11148), .B1_f (new_AGEMA_signal_11149), .Z0_t (SubBytesIns_Inst_Sbox_0_L15), .Z0_f (new_AGEMA_signal_11837), .Z1_t (new_AGEMA_signal_11838), .Z1_f (new_AGEMA_signal_11839) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M56), .A0_f (new_AGEMA_signal_10424), .A1_t (new_AGEMA_signal_10425), .A1_f (new_AGEMA_signal_10426), .B0_t (SubBytesIns_Inst_Sbox_0_L0), .B0_f (new_AGEMA_signal_12404), .B1_t (new_AGEMA_signal_12405), .B1_f (new_AGEMA_signal_12406), .Z0_t (SubBytesIns_Inst_Sbox_0_L16), .Z0_f (new_AGEMA_signal_12971), .Z1_t (new_AGEMA_signal_12972), .Z1_f (new_AGEMA_signal_12973) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M57), .A0_f (new_AGEMA_signal_10427), .A1_t (new_AGEMA_signal_10428), .A1_f (new_AGEMA_signal_10429), .B0_t (SubBytesIns_Inst_Sbox_0_L1), .B0_f (new_AGEMA_signal_11147), .B1_t (new_AGEMA_signal_11148), .B1_f (new_AGEMA_signal_11149), .Z0_t (SubBytesIns_Inst_Sbox_0_L17), .Z0_f (new_AGEMA_signal_11840), .Z1_t (new_AGEMA_signal_11841), .Z1_f (new_AGEMA_signal_11842) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M58), .A0_f (new_AGEMA_signal_11138), .A1_t (new_AGEMA_signal_11139), .A1_f (new_AGEMA_signal_11140), .B0_t (SubBytesIns_Inst_Sbox_0_L8), .B0_f (new_AGEMA_signal_11150), .B1_t (new_AGEMA_signal_11151), .B1_f (new_AGEMA_signal_11152), .Z0_t (SubBytesIns_Inst_Sbox_0_L18), .Z0_f (new_AGEMA_signal_11843), .Z1_t (new_AGEMA_signal_11844), .Z1_f (new_AGEMA_signal_11845) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M63), .A0_f (new_AGEMA_signal_11144), .A1_t (new_AGEMA_signal_11145), .A1_f (new_AGEMA_signal_11146), .B0_t (SubBytesIns_Inst_Sbox_0_L4), .B0_f (new_AGEMA_signal_11828), .B1_t (new_AGEMA_signal_11829), .B1_f (new_AGEMA_signal_11830), .Z0_t (SubBytesIns_Inst_Sbox_0_L19), .Z0_f (new_AGEMA_signal_12422), .Z1_t (new_AGEMA_signal_12423), .Z1_f (new_AGEMA_signal_12424) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L0), .A0_f (new_AGEMA_signal_12404), .A1_t (new_AGEMA_signal_12405), .A1_f (new_AGEMA_signal_12406), .B0_t (SubBytesIns_Inst_Sbox_0_L1), .B0_f (new_AGEMA_signal_11147), .B1_t (new_AGEMA_signal_11148), .B1_f (new_AGEMA_signal_11149), .Z0_t (SubBytesIns_Inst_Sbox_0_L20), .Z0_f (new_AGEMA_signal_12974), .Z1_t (new_AGEMA_signal_12975), .Z1_f (new_AGEMA_signal_12976) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L1), .A0_f (new_AGEMA_signal_11147), .A1_t (new_AGEMA_signal_11148), .A1_f (new_AGEMA_signal_11149), .B0_t (SubBytesIns_Inst_Sbox_0_L7), .B0_f (new_AGEMA_signal_12410), .B1_t (new_AGEMA_signal_12411), .B1_f (new_AGEMA_signal_12412), .Z0_t (SubBytesIns_Inst_Sbox_0_L21), .Z0_f (new_AGEMA_signal_12977), .Z1_t (new_AGEMA_signal_12978), .Z1_f (new_AGEMA_signal_12979) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L3), .A0_f (new_AGEMA_signal_11825), .A1_t (new_AGEMA_signal_11826), .A1_f (new_AGEMA_signal_11827), .B0_t (SubBytesIns_Inst_Sbox_0_L12), .B0_f (new_AGEMA_signal_11153), .B1_t (new_AGEMA_signal_11154), .B1_f (new_AGEMA_signal_11155), .Z0_t (SubBytesIns_Inst_Sbox_0_L22), .Z0_f (new_AGEMA_signal_12425), .Z1_t (new_AGEMA_signal_12426), .Z1_f (new_AGEMA_signal_12427) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L18), .A0_f (new_AGEMA_signal_11843), .A1_t (new_AGEMA_signal_11844), .A1_f (new_AGEMA_signal_11845), .B0_t (SubBytesIns_Inst_Sbox_0_L2), .B0_f (new_AGEMA_signal_11822), .B1_t (new_AGEMA_signal_11823), .B1_f (new_AGEMA_signal_11824), .Z0_t (SubBytesIns_Inst_Sbox_0_L23), .Z0_f (new_AGEMA_signal_12428), .Z1_t (new_AGEMA_signal_12429), .Z1_f (new_AGEMA_signal_12430) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L15), .A0_f (new_AGEMA_signal_11837), .A1_t (new_AGEMA_signal_11838), .A1_f (new_AGEMA_signal_11839), .B0_t (SubBytesIns_Inst_Sbox_0_L9), .B0_f (new_AGEMA_signal_12413), .B1_t (new_AGEMA_signal_12414), .B1_f (new_AGEMA_signal_12415), .Z0_t (SubBytesIns_Inst_Sbox_0_L24), .Z0_f (new_AGEMA_signal_12980), .Z1_t (new_AGEMA_signal_12981), .Z1_f (new_AGEMA_signal_12982) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L6), .A0_f (new_AGEMA_signal_12407), .A1_t (new_AGEMA_signal_12408), .A1_f (new_AGEMA_signal_12409), .B0_t (SubBytesIns_Inst_Sbox_0_L10), .B0_f (new_AGEMA_signal_12416), .B1_t (new_AGEMA_signal_12417), .B1_f (new_AGEMA_signal_12418), .Z0_t (SubBytesIns_Inst_Sbox_0_L25), .Z0_f (new_AGEMA_signal_12983), .Z1_t (new_AGEMA_signal_12984), .Z1_f (new_AGEMA_signal_12985) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L7), .A0_f (new_AGEMA_signal_12410), .A1_t (new_AGEMA_signal_12411), .A1_f (new_AGEMA_signal_12412), .B0_t (SubBytesIns_Inst_Sbox_0_L9), .B0_f (new_AGEMA_signal_12413), .B1_t (new_AGEMA_signal_12414), .B1_f (new_AGEMA_signal_12415), .Z0_t (SubBytesIns_Inst_Sbox_0_L26), .Z0_f (new_AGEMA_signal_12986), .Z1_t (new_AGEMA_signal_12987), .Z1_f (new_AGEMA_signal_12988) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L8), .A0_f (new_AGEMA_signal_11150), .A1_t (new_AGEMA_signal_11151), .A1_f (new_AGEMA_signal_11152), .B0_t (SubBytesIns_Inst_Sbox_0_L10), .B0_f (new_AGEMA_signal_12416), .B1_t (new_AGEMA_signal_12417), .B1_f (new_AGEMA_signal_12418), .Z0_t (SubBytesIns_Inst_Sbox_0_L27), .Z0_f (new_AGEMA_signal_12989), .Z1_t (new_AGEMA_signal_12990), .Z1_f (new_AGEMA_signal_12991) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L11), .A0_f (new_AGEMA_signal_12419), .A1_t (new_AGEMA_signal_12420), .A1_f (new_AGEMA_signal_12421), .B0_t (SubBytesIns_Inst_Sbox_0_L14), .B0_f (new_AGEMA_signal_11834), .B1_t (new_AGEMA_signal_11835), .B1_f (new_AGEMA_signal_11836), .Z0_t (SubBytesIns_Inst_Sbox_0_L28), .Z0_f (new_AGEMA_signal_12992), .Z1_t (new_AGEMA_signal_12993), .Z1_f (new_AGEMA_signal_12994) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L11), .A0_f (new_AGEMA_signal_12419), .A1_t (new_AGEMA_signal_12420), .A1_f (new_AGEMA_signal_12421), .B0_t (SubBytesIns_Inst_Sbox_0_L17), .B0_f (new_AGEMA_signal_11840), .B1_t (new_AGEMA_signal_11841), .B1_f (new_AGEMA_signal_11842), .Z0_t (SubBytesIns_Inst_Sbox_0_L29), .Z0_f (new_AGEMA_signal_12995), .Z1_t (new_AGEMA_signal_12996), .Z1_f (new_AGEMA_signal_12997) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L6), .A0_f (new_AGEMA_signal_12407), .A1_t (new_AGEMA_signal_12408), .A1_f (new_AGEMA_signal_12409), .B0_t (SubBytesIns_Inst_Sbox_0_L24), .B0_f (new_AGEMA_signal_12980), .B1_t (new_AGEMA_signal_12981), .B1_f (new_AGEMA_signal_12982), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .Z0_f (new_AGEMA_signal_13640), .Z1_t (new_AGEMA_signal_13641), .Z1_f (new_AGEMA_signal_13642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L16), .A0_f (new_AGEMA_signal_12971), .A1_t (new_AGEMA_signal_12972), .A1_f (new_AGEMA_signal_12973), .B0_t (SubBytesIns_Inst_Sbox_0_L26), .B0_f (new_AGEMA_signal_12986), .B1_t (new_AGEMA_signal_12987), .B1_f (new_AGEMA_signal_12988), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .Z0_f (new_AGEMA_signal_13643), .Z1_t (new_AGEMA_signal_13644), .Z1_f (new_AGEMA_signal_13645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L19), .A0_f (new_AGEMA_signal_12422), .A1_t (new_AGEMA_signal_12423), .A1_f (new_AGEMA_signal_12424), .B0_t (SubBytesIns_Inst_Sbox_0_L28), .B0_f (new_AGEMA_signal_12992), .B1_t (new_AGEMA_signal_12993), .B1_f (new_AGEMA_signal_12994), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .Z0_f (new_AGEMA_signal_13646), .Z1_t (new_AGEMA_signal_13647), .Z1_f (new_AGEMA_signal_13648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L6), .A0_f (new_AGEMA_signal_12407), .A1_t (new_AGEMA_signal_12408), .A1_f (new_AGEMA_signal_12409), .B0_t (SubBytesIns_Inst_Sbox_0_L21), .B0_f (new_AGEMA_signal_12977), .B1_t (new_AGEMA_signal_12978), .B1_f (new_AGEMA_signal_12979), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .Z0_f (new_AGEMA_signal_13649), .Z1_t (new_AGEMA_signal_13650), .Z1_f (new_AGEMA_signal_13651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L20), .A0_f (new_AGEMA_signal_12974), .A1_t (new_AGEMA_signal_12975), .A1_f (new_AGEMA_signal_12976), .B0_t (SubBytesIns_Inst_Sbox_0_L22), .B0_f (new_AGEMA_signal_12425), .B1_t (new_AGEMA_signal_12426), .B1_f (new_AGEMA_signal_12427), .Z0_t (MixColumnsInput[99]), .Z0_f (new_AGEMA_signal_13652), .Z1_t (new_AGEMA_signal_13653), .Z1_f (new_AGEMA_signal_13654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L25), .A0_f (new_AGEMA_signal_12983), .A1_t (new_AGEMA_signal_12984), .A1_f (new_AGEMA_signal_12985), .B0_t (SubBytesIns_Inst_Sbox_0_L29), .B0_f (new_AGEMA_signal_12995), .B1_t (new_AGEMA_signal_12996), .B1_f (new_AGEMA_signal_12997), .Z0_t (MixColumnsInput[98]), .Z0_f (new_AGEMA_signal_13655), .Z1_t (new_AGEMA_signal_13656), .Z1_f (new_AGEMA_signal_13657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L13), .A0_f (new_AGEMA_signal_12968), .A1_t (new_AGEMA_signal_12969), .A1_f (new_AGEMA_signal_12970), .B0_t (SubBytesIns_Inst_Sbox_0_L27), .B0_f (new_AGEMA_signal_12989), .B1_t (new_AGEMA_signal_12990), .B1_f (new_AGEMA_signal_12991), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .Z0_f (new_AGEMA_signal_13658), .Z1_t (new_AGEMA_signal_13659), .Z1_f (new_AGEMA_signal_13660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L6), .A0_f (new_AGEMA_signal_12407), .A1_t (new_AGEMA_signal_12408), .A1_f (new_AGEMA_signal_12409), .B0_t (SubBytesIns_Inst_Sbox_0_L23), .B0_f (new_AGEMA_signal_12428), .B1_t (new_AGEMA_signal_12429), .B1_f (new_AGEMA_signal_12430), .Z0_t (MixColumnsInput[96]), .Z0_f (new_AGEMA_signal_12998), .Z1_t (new_AGEMA_signal_12999), .Z1_f (new_AGEMA_signal_13000) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[15]), .A0_f (ciphertext_s0_f[15]), .A1_t (ciphertext_s1_t[15]), .A1_f (ciphertext_s1_f[15]), .B0_t (ciphertext_s0_t[12]), .B0_f (ciphertext_s0_f[12]), .B1_t (ciphertext_s1_t[12]), .B1_f (ciphertext_s1_f[12]), .Z0_t (SubBytesIns_Inst_Sbox_1_T1), .Z0_f (new_AGEMA_signal_6376), .Z1_t (new_AGEMA_signal_6377), .Z1_f (new_AGEMA_signal_6378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[15]), .A0_f (ciphertext_s0_f[15]), .A1_t (ciphertext_s1_t[15]), .A1_f (ciphertext_s1_f[15]), .B0_t (ciphertext_s0_t[10]), .B0_f (ciphertext_s0_f[10]), .B1_t (ciphertext_s1_t[10]), .B1_f (ciphertext_s1_f[10]), .Z0_t (SubBytesIns_Inst_Sbox_1_T2), .Z0_f (new_AGEMA_signal_6379), .Z1_t (new_AGEMA_signal_6380), .Z1_f (new_AGEMA_signal_6381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[15]), .A0_f (ciphertext_s0_f[15]), .A1_t (ciphertext_s1_t[15]), .A1_f (ciphertext_s1_f[15]), .B0_t (ciphertext_s0_t[9]), .B0_f (ciphertext_s0_f[9]), .B1_t (ciphertext_s1_t[9]), .B1_f (ciphertext_s1_f[9]), .Z0_t (SubBytesIns_Inst_Sbox_1_T3), .Z0_f (new_AGEMA_signal_6382), .Z1_t (new_AGEMA_signal_6383), .Z1_f (new_AGEMA_signal_6384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[12]), .A0_f (ciphertext_s0_f[12]), .A1_t (ciphertext_s1_t[12]), .A1_f (ciphertext_s1_f[12]), .B0_t (ciphertext_s0_t[10]), .B0_f (ciphertext_s0_f[10]), .B1_t (ciphertext_s1_t[10]), .B1_f (ciphertext_s1_f[10]), .Z0_t (SubBytesIns_Inst_Sbox_1_T4), .Z0_f (new_AGEMA_signal_6385), .Z1_t (new_AGEMA_signal_6386), .Z1_f (new_AGEMA_signal_6387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[11]), .A0_f (ciphertext_s0_f[11]), .A1_t (ciphertext_s1_t[11]), .A1_f (ciphertext_s1_f[11]), .B0_t (ciphertext_s0_t[9]), .B0_f (ciphertext_s0_f[9]), .B1_t (ciphertext_s1_t[9]), .B1_f (ciphertext_s1_f[9]), .Z0_t (SubBytesIns_Inst_Sbox_1_T5), .Z0_f (new_AGEMA_signal_6388), .Z1_t (new_AGEMA_signal_6389), .Z1_f (new_AGEMA_signal_6390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T1), .A0_f (new_AGEMA_signal_6376), .A1_t (new_AGEMA_signal_6377), .A1_f (new_AGEMA_signal_6378), .B0_t (SubBytesIns_Inst_Sbox_1_T5), .B0_f (new_AGEMA_signal_6388), .B1_t (new_AGEMA_signal_6389), .B1_f (new_AGEMA_signal_6390), .Z0_t (SubBytesIns_Inst_Sbox_1_T6), .Z0_f (new_AGEMA_signal_6952), .Z1_t (new_AGEMA_signal_6953), .Z1_f (new_AGEMA_signal_6954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[14]), .A0_f (ciphertext_s0_f[14]), .A1_t (ciphertext_s1_t[14]), .A1_f (ciphertext_s1_f[14]), .B0_t (ciphertext_s0_t[13]), .B0_f (ciphertext_s0_f[13]), .B1_t (ciphertext_s1_t[13]), .B1_f (ciphertext_s1_f[13]), .Z0_t (SubBytesIns_Inst_Sbox_1_T7), .Z0_f (new_AGEMA_signal_6391), .Z1_t (new_AGEMA_signal_6392), .Z1_f (new_AGEMA_signal_6393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[8]), .A0_f (ciphertext_s0_f[8]), .A1_t (ciphertext_s1_t[8]), .A1_f (ciphertext_s1_f[8]), .B0_t (SubBytesIns_Inst_Sbox_1_T6), .B0_f (new_AGEMA_signal_6952), .B1_t (new_AGEMA_signal_6953), .B1_f (new_AGEMA_signal_6954), .Z0_t (SubBytesIns_Inst_Sbox_1_T8), .Z0_f (new_AGEMA_signal_7511), .Z1_t (new_AGEMA_signal_7512), .Z1_f (new_AGEMA_signal_7513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[8]), .A0_f (ciphertext_s0_f[8]), .A1_t (ciphertext_s1_t[8]), .A1_f (ciphertext_s1_f[8]), .B0_t (SubBytesIns_Inst_Sbox_1_T7), .B0_f (new_AGEMA_signal_6391), .B1_t (new_AGEMA_signal_6392), .B1_f (new_AGEMA_signal_6393), .Z0_t (SubBytesIns_Inst_Sbox_1_T9), .Z0_f (new_AGEMA_signal_6955), .Z1_t (new_AGEMA_signal_6956), .Z1_f (new_AGEMA_signal_6957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T6), .A0_f (new_AGEMA_signal_6952), .A1_t (new_AGEMA_signal_6953), .A1_f (new_AGEMA_signal_6954), .B0_t (SubBytesIns_Inst_Sbox_1_T7), .B0_f (new_AGEMA_signal_6391), .B1_t (new_AGEMA_signal_6392), .B1_f (new_AGEMA_signal_6393), .Z0_t (SubBytesIns_Inst_Sbox_1_T10), .Z0_f (new_AGEMA_signal_7514), .Z1_t (new_AGEMA_signal_7515), .Z1_f (new_AGEMA_signal_7516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[14]), .A0_f (ciphertext_s0_f[14]), .A1_t (ciphertext_s1_t[14]), .A1_f (ciphertext_s1_f[14]), .B0_t (ciphertext_s0_t[10]), .B0_f (ciphertext_s0_f[10]), .B1_t (ciphertext_s1_t[10]), .B1_f (ciphertext_s1_f[10]), .Z0_t (SubBytesIns_Inst_Sbox_1_T11), .Z0_f (new_AGEMA_signal_6394), .Z1_t (new_AGEMA_signal_6395), .Z1_f (new_AGEMA_signal_6396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[13]), .A0_f (ciphertext_s0_f[13]), .A1_t (ciphertext_s1_t[13]), .A1_f (ciphertext_s1_f[13]), .B0_t (ciphertext_s0_t[10]), .B0_f (ciphertext_s0_f[10]), .B1_t (ciphertext_s1_t[10]), .B1_f (ciphertext_s1_f[10]), .Z0_t (SubBytesIns_Inst_Sbox_1_T12), .Z0_f (new_AGEMA_signal_6397), .Z1_t (new_AGEMA_signal_6398), .Z1_f (new_AGEMA_signal_6399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T3), .A0_f (new_AGEMA_signal_6382), .A1_t (new_AGEMA_signal_6383), .A1_f (new_AGEMA_signal_6384), .B0_t (SubBytesIns_Inst_Sbox_1_T4), .B0_f (new_AGEMA_signal_6385), .B1_t (new_AGEMA_signal_6386), .B1_f (new_AGEMA_signal_6387), .Z0_t (SubBytesIns_Inst_Sbox_1_T13), .Z0_f (new_AGEMA_signal_6958), .Z1_t (new_AGEMA_signal_6959), .Z1_f (new_AGEMA_signal_6960) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T6), .A0_f (new_AGEMA_signal_6952), .A1_t (new_AGEMA_signal_6953), .A1_f (new_AGEMA_signal_6954), .B0_t (SubBytesIns_Inst_Sbox_1_T11), .B0_f (new_AGEMA_signal_6394), .B1_t (new_AGEMA_signal_6395), .B1_f (new_AGEMA_signal_6396), .Z0_t (SubBytesIns_Inst_Sbox_1_T14), .Z0_f (new_AGEMA_signal_7517), .Z1_t (new_AGEMA_signal_7518), .Z1_f (new_AGEMA_signal_7519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T5), .A0_f (new_AGEMA_signal_6388), .A1_t (new_AGEMA_signal_6389), .A1_f (new_AGEMA_signal_6390), .B0_t (SubBytesIns_Inst_Sbox_1_T11), .B0_f (new_AGEMA_signal_6394), .B1_t (new_AGEMA_signal_6395), .B1_f (new_AGEMA_signal_6396), .Z0_t (SubBytesIns_Inst_Sbox_1_T15), .Z0_f (new_AGEMA_signal_6961), .Z1_t (new_AGEMA_signal_6962), .Z1_f (new_AGEMA_signal_6963) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T5), .A0_f (new_AGEMA_signal_6388), .A1_t (new_AGEMA_signal_6389), .A1_f (new_AGEMA_signal_6390), .B0_t (SubBytesIns_Inst_Sbox_1_T12), .B0_f (new_AGEMA_signal_6397), .B1_t (new_AGEMA_signal_6398), .B1_f (new_AGEMA_signal_6399), .Z0_t (SubBytesIns_Inst_Sbox_1_T16), .Z0_f (new_AGEMA_signal_6964), .Z1_t (new_AGEMA_signal_6965), .Z1_f (new_AGEMA_signal_6966) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T9), .A0_f (new_AGEMA_signal_6955), .A1_t (new_AGEMA_signal_6956), .A1_f (new_AGEMA_signal_6957), .B0_t (SubBytesIns_Inst_Sbox_1_T16), .B0_f (new_AGEMA_signal_6964), .B1_t (new_AGEMA_signal_6965), .B1_f (new_AGEMA_signal_6966), .Z0_t (SubBytesIns_Inst_Sbox_1_T17), .Z0_f (new_AGEMA_signal_7520), .Z1_t (new_AGEMA_signal_7521), .Z1_f (new_AGEMA_signal_7522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[12]), .A0_f (ciphertext_s0_f[12]), .A1_t (ciphertext_s1_t[12]), .A1_f (ciphertext_s1_f[12]), .B0_t (ciphertext_s0_t[8]), .B0_f (ciphertext_s0_f[8]), .B1_t (ciphertext_s1_t[8]), .B1_f (ciphertext_s1_f[8]), .Z0_t (SubBytesIns_Inst_Sbox_1_T18), .Z0_f (new_AGEMA_signal_6400), .Z1_t (new_AGEMA_signal_6401), .Z1_f (new_AGEMA_signal_6402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T7), .A0_f (new_AGEMA_signal_6391), .A1_t (new_AGEMA_signal_6392), .A1_f (new_AGEMA_signal_6393), .B0_t (SubBytesIns_Inst_Sbox_1_T18), .B0_f (new_AGEMA_signal_6400), .B1_t (new_AGEMA_signal_6401), .B1_f (new_AGEMA_signal_6402), .Z0_t (SubBytesIns_Inst_Sbox_1_T19), .Z0_f (new_AGEMA_signal_6967), .Z1_t (new_AGEMA_signal_6968), .Z1_f (new_AGEMA_signal_6969) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T1), .A0_f (new_AGEMA_signal_6376), .A1_t (new_AGEMA_signal_6377), .A1_f (new_AGEMA_signal_6378), .B0_t (SubBytesIns_Inst_Sbox_1_T19), .B0_f (new_AGEMA_signal_6967), .B1_t (new_AGEMA_signal_6968), .B1_f (new_AGEMA_signal_6969), .Z0_t (SubBytesIns_Inst_Sbox_1_T20), .Z0_f (new_AGEMA_signal_7523), .Z1_t (new_AGEMA_signal_7524), .Z1_f (new_AGEMA_signal_7525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[9]), .A0_f (ciphertext_s0_f[9]), .A1_t (ciphertext_s1_t[9]), .A1_f (ciphertext_s1_f[9]), .B0_t (ciphertext_s0_t[8]), .B0_f (ciphertext_s0_f[8]), .B1_t (ciphertext_s1_t[8]), .B1_f (ciphertext_s1_f[8]), .Z0_t (SubBytesIns_Inst_Sbox_1_T21), .Z0_f (new_AGEMA_signal_6403), .Z1_t (new_AGEMA_signal_6404), .Z1_f (new_AGEMA_signal_6405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T7), .A0_f (new_AGEMA_signal_6391), .A1_t (new_AGEMA_signal_6392), .A1_f (new_AGEMA_signal_6393), .B0_t (SubBytesIns_Inst_Sbox_1_T21), .B0_f (new_AGEMA_signal_6403), .B1_t (new_AGEMA_signal_6404), .B1_f (new_AGEMA_signal_6405), .Z0_t (SubBytesIns_Inst_Sbox_1_T22), .Z0_f (new_AGEMA_signal_6970), .Z1_t (new_AGEMA_signal_6971), .Z1_f (new_AGEMA_signal_6972) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T2), .A0_f (new_AGEMA_signal_6379), .A1_t (new_AGEMA_signal_6380), .A1_f (new_AGEMA_signal_6381), .B0_t (SubBytesIns_Inst_Sbox_1_T22), .B0_f (new_AGEMA_signal_6970), .B1_t (new_AGEMA_signal_6971), .B1_f (new_AGEMA_signal_6972), .Z0_t (SubBytesIns_Inst_Sbox_1_T23), .Z0_f (new_AGEMA_signal_7526), .Z1_t (new_AGEMA_signal_7527), .Z1_f (new_AGEMA_signal_7528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T2), .A0_f (new_AGEMA_signal_6379), .A1_t (new_AGEMA_signal_6380), .A1_f (new_AGEMA_signal_6381), .B0_t (SubBytesIns_Inst_Sbox_1_T10), .B0_f (new_AGEMA_signal_7514), .B1_t (new_AGEMA_signal_7515), .B1_f (new_AGEMA_signal_7516), .Z0_t (SubBytesIns_Inst_Sbox_1_T24), .Z0_f (new_AGEMA_signal_8231), .Z1_t (new_AGEMA_signal_8232), .Z1_f (new_AGEMA_signal_8233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T20), .A0_f (new_AGEMA_signal_7523), .A1_t (new_AGEMA_signal_7524), .A1_f (new_AGEMA_signal_7525), .B0_t (SubBytesIns_Inst_Sbox_1_T17), .B0_f (new_AGEMA_signal_7520), .B1_t (new_AGEMA_signal_7521), .B1_f (new_AGEMA_signal_7522), .Z0_t (SubBytesIns_Inst_Sbox_1_T25), .Z0_f (new_AGEMA_signal_8234), .Z1_t (new_AGEMA_signal_8235), .Z1_f (new_AGEMA_signal_8236) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T3), .A0_f (new_AGEMA_signal_6382), .A1_t (new_AGEMA_signal_6383), .A1_f (new_AGEMA_signal_6384), .B0_t (SubBytesIns_Inst_Sbox_1_T16), .B0_f (new_AGEMA_signal_6964), .B1_t (new_AGEMA_signal_6965), .B1_f (new_AGEMA_signal_6966), .Z0_t (SubBytesIns_Inst_Sbox_1_T26), .Z0_f (new_AGEMA_signal_7529), .Z1_t (new_AGEMA_signal_7530), .Z1_f (new_AGEMA_signal_7531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T1), .A0_f (new_AGEMA_signal_6376), .A1_t (new_AGEMA_signal_6377), .A1_f (new_AGEMA_signal_6378), .B0_t (SubBytesIns_Inst_Sbox_1_T12), .B0_f (new_AGEMA_signal_6397), .B1_t (new_AGEMA_signal_6398), .B1_f (new_AGEMA_signal_6399), .Z0_t (SubBytesIns_Inst_Sbox_1_T27), .Z0_f (new_AGEMA_signal_6973), .Z1_t (new_AGEMA_signal_6974), .Z1_f (new_AGEMA_signal_6975) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T13), .A0_f (new_AGEMA_signal_6958), .A1_t (new_AGEMA_signal_6959), .A1_f (new_AGEMA_signal_6960), .B0_t (SubBytesIns_Inst_Sbox_1_T6), .B0_f (new_AGEMA_signal_6952), .B1_t (new_AGEMA_signal_6953), .B1_f (new_AGEMA_signal_6954), .Z0_t (SubBytesIns_Inst_Sbox_1_M1), .Z0_f (new_AGEMA_signal_7532), .Z1_t (new_AGEMA_signal_7533), .Z1_f (new_AGEMA_signal_7534) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T23), .A0_f (new_AGEMA_signal_7526), .A1_t (new_AGEMA_signal_7527), .A1_f (new_AGEMA_signal_7528), .B0_t (SubBytesIns_Inst_Sbox_1_T8), .B0_f (new_AGEMA_signal_7511), .B1_t (new_AGEMA_signal_7512), .B1_f (new_AGEMA_signal_7513), .Z0_t (SubBytesIns_Inst_Sbox_1_M2), .Z0_f (new_AGEMA_signal_8237), .Z1_t (new_AGEMA_signal_8238), .Z1_f (new_AGEMA_signal_8239) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T14), .A0_f (new_AGEMA_signal_7517), .A1_t (new_AGEMA_signal_7518), .A1_f (new_AGEMA_signal_7519), .B0_t (SubBytesIns_Inst_Sbox_1_M1), .B0_f (new_AGEMA_signal_7532), .B1_t (new_AGEMA_signal_7533), .B1_f (new_AGEMA_signal_7534), .Z0_t (SubBytesIns_Inst_Sbox_1_M3), .Z0_f (new_AGEMA_signal_8240), .Z1_t (new_AGEMA_signal_8241), .Z1_f (new_AGEMA_signal_8242) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T19), .A0_f (new_AGEMA_signal_6967), .A1_t (new_AGEMA_signal_6968), .A1_f (new_AGEMA_signal_6969), .B0_t (ciphertext_s0_t[8]), .B0_f (ciphertext_s0_f[8]), .B1_t (ciphertext_s1_t[8]), .B1_f (ciphertext_s1_f[8]), .Z0_t (SubBytesIns_Inst_Sbox_1_M4), .Z0_f (new_AGEMA_signal_7535), .Z1_t (new_AGEMA_signal_7536), .Z1_f (new_AGEMA_signal_7537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M4), .A0_f (new_AGEMA_signal_7535), .A1_t (new_AGEMA_signal_7536), .A1_f (new_AGEMA_signal_7537), .B0_t (SubBytesIns_Inst_Sbox_1_M1), .B0_f (new_AGEMA_signal_7532), .B1_t (new_AGEMA_signal_7533), .B1_f (new_AGEMA_signal_7534), .Z0_t (SubBytesIns_Inst_Sbox_1_M5), .Z0_f (new_AGEMA_signal_8243), .Z1_t (new_AGEMA_signal_8244), .Z1_f (new_AGEMA_signal_8245) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T3), .A0_f (new_AGEMA_signal_6382), .A1_t (new_AGEMA_signal_6383), .A1_f (new_AGEMA_signal_6384), .B0_t (SubBytesIns_Inst_Sbox_1_T16), .B0_f (new_AGEMA_signal_6964), .B1_t (new_AGEMA_signal_6965), .B1_f (new_AGEMA_signal_6966), .Z0_t (SubBytesIns_Inst_Sbox_1_M6), .Z0_f (new_AGEMA_signal_7538), .Z1_t (new_AGEMA_signal_7539), .Z1_f (new_AGEMA_signal_7540) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T22), .A0_f (new_AGEMA_signal_6970), .A1_t (new_AGEMA_signal_6971), .A1_f (new_AGEMA_signal_6972), .B0_t (SubBytesIns_Inst_Sbox_1_T9), .B0_f (new_AGEMA_signal_6955), .B1_t (new_AGEMA_signal_6956), .B1_f (new_AGEMA_signal_6957), .Z0_t (SubBytesIns_Inst_Sbox_1_M7), .Z0_f (new_AGEMA_signal_7541), .Z1_t (new_AGEMA_signal_7542), .Z1_f (new_AGEMA_signal_7543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T26), .A0_f (new_AGEMA_signal_7529), .A1_t (new_AGEMA_signal_7530), .A1_f (new_AGEMA_signal_7531), .B0_t (SubBytesIns_Inst_Sbox_1_M6), .B0_f (new_AGEMA_signal_7538), .B1_t (new_AGEMA_signal_7539), .B1_f (new_AGEMA_signal_7540), .Z0_t (SubBytesIns_Inst_Sbox_1_M8), .Z0_f (new_AGEMA_signal_8246), .Z1_t (new_AGEMA_signal_8247), .Z1_f (new_AGEMA_signal_8248) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T20), .A0_f (new_AGEMA_signal_7523), .A1_t (new_AGEMA_signal_7524), .A1_f (new_AGEMA_signal_7525), .B0_t (SubBytesIns_Inst_Sbox_1_T17), .B0_f (new_AGEMA_signal_7520), .B1_t (new_AGEMA_signal_7521), .B1_f (new_AGEMA_signal_7522), .Z0_t (SubBytesIns_Inst_Sbox_1_M9), .Z0_f (new_AGEMA_signal_8249), .Z1_t (new_AGEMA_signal_8250), .Z1_f (new_AGEMA_signal_8251) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M9), .A0_f (new_AGEMA_signal_8249), .A1_t (new_AGEMA_signal_8250), .A1_f (new_AGEMA_signal_8251), .B0_t (SubBytesIns_Inst_Sbox_1_M6), .B0_f (new_AGEMA_signal_7538), .B1_t (new_AGEMA_signal_7539), .B1_f (new_AGEMA_signal_7540), .Z0_t (SubBytesIns_Inst_Sbox_1_M10), .Z0_f (new_AGEMA_signal_8711), .Z1_t (new_AGEMA_signal_8712), .Z1_f (new_AGEMA_signal_8713) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T1), .A0_f (new_AGEMA_signal_6376), .A1_t (new_AGEMA_signal_6377), .A1_f (new_AGEMA_signal_6378), .B0_t (SubBytesIns_Inst_Sbox_1_T15), .B0_f (new_AGEMA_signal_6961), .B1_t (new_AGEMA_signal_6962), .B1_f (new_AGEMA_signal_6963), .Z0_t (SubBytesIns_Inst_Sbox_1_M11), .Z0_f (new_AGEMA_signal_7544), .Z1_t (new_AGEMA_signal_7545), .Z1_f (new_AGEMA_signal_7546) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T4), .A0_f (new_AGEMA_signal_6385), .A1_t (new_AGEMA_signal_6386), .A1_f (new_AGEMA_signal_6387), .B0_t (SubBytesIns_Inst_Sbox_1_T27), .B0_f (new_AGEMA_signal_6973), .B1_t (new_AGEMA_signal_6974), .B1_f (new_AGEMA_signal_6975), .Z0_t (SubBytesIns_Inst_Sbox_1_M12), .Z0_f (new_AGEMA_signal_7547), .Z1_t (new_AGEMA_signal_7548), .Z1_f (new_AGEMA_signal_7549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M12), .A0_f (new_AGEMA_signal_7547), .A1_t (new_AGEMA_signal_7548), .A1_f (new_AGEMA_signal_7549), .B0_t (SubBytesIns_Inst_Sbox_1_M11), .B0_f (new_AGEMA_signal_7544), .B1_t (new_AGEMA_signal_7545), .B1_f (new_AGEMA_signal_7546), .Z0_t (SubBytesIns_Inst_Sbox_1_M13), .Z0_f (new_AGEMA_signal_8252), .Z1_t (new_AGEMA_signal_8253), .Z1_f (new_AGEMA_signal_8254) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T2), .A0_f (new_AGEMA_signal_6379), .A1_t (new_AGEMA_signal_6380), .A1_f (new_AGEMA_signal_6381), .B0_t (SubBytesIns_Inst_Sbox_1_T10), .B0_f (new_AGEMA_signal_7514), .B1_t (new_AGEMA_signal_7515), .B1_f (new_AGEMA_signal_7516), .Z0_t (SubBytesIns_Inst_Sbox_1_M14), .Z0_f (new_AGEMA_signal_8255), .Z1_t (new_AGEMA_signal_8256), .Z1_f (new_AGEMA_signal_8257) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M14), .A0_f (new_AGEMA_signal_8255), .A1_t (new_AGEMA_signal_8256), .A1_f (new_AGEMA_signal_8257), .B0_t (SubBytesIns_Inst_Sbox_1_M11), .B0_f (new_AGEMA_signal_7544), .B1_t (new_AGEMA_signal_7545), .B1_f (new_AGEMA_signal_7546), .Z0_t (SubBytesIns_Inst_Sbox_1_M15), .Z0_f (new_AGEMA_signal_8714), .Z1_t (new_AGEMA_signal_8715), .Z1_f (new_AGEMA_signal_8716) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M3), .A0_f (new_AGEMA_signal_8240), .A1_t (new_AGEMA_signal_8241), .A1_f (new_AGEMA_signal_8242), .B0_t (SubBytesIns_Inst_Sbox_1_M2), .B0_f (new_AGEMA_signal_8237), .B1_t (new_AGEMA_signal_8238), .B1_f (new_AGEMA_signal_8239), .Z0_t (SubBytesIns_Inst_Sbox_1_M16), .Z0_f (new_AGEMA_signal_8717), .Z1_t (new_AGEMA_signal_8718), .Z1_f (new_AGEMA_signal_8719) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M5), .A0_f (new_AGEMA_signal_8243), .A1_t (new_AGEMA_signal_8244), .A1_f (new_AGEMA_signal_8245), .B0_t (SubBytesIns_Inst_Sbox_1_T24), .B0_f (new_AGEMA_signal_8231), .B1_t (new_AGEMA_signal_8232), .B1_f (new_AGEMA_signal_8233), .Z0_t (SubBytesIns_Inst_Sbox_1_M17), .Z0_f (new_AGEMA_signal_8720), .Z1_t (new_AGEMA_signal_8721), .Z1_f (new_AGEMA_signal_8722) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M8), .A0_f (new_AGEMA_signal_8246), .A1_t (new_AGEMA_signal_8247), .A1_f (new_AGEMA_signal_8248), .B0_t (SubBytesIns_Inst_Sbox_1_M7), .B0_f (new_AGEMA_signal_7541), .B1_t (new_AGEMA_signal_7542), .B1_f (new_AGEMA_signal_7543), .Z0_t (SubBytesIns_Inst_Sbox_1_M18), .Z0_f (new_AGEMA_signal_8723), .Z1_t (new_AGEMA_signal_8724), .Z1_f (new_AGEMA_signal_8725) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M10), .A0_f (new_AGEMA_signal_8711), .A1_t (new_AGEMA_signal_8712), .A1_f (new_AGEMA_signal_8713), .B0_t (SubBytesIns_Inst_Sbox_1_M15), .B0_f (new_AGEMA_signal_8714), .B1_t (new_AGEMA_signal_8715), .B1_f (new_AGEMA_signal_8716), .Z0_t (SubBytesIns_Inst_Sbox_1_M19), .Z0_f (new_AGEMA_signal_8996), .Z1_t (new_AGEMA_signal_8997), .Z1_f (new_AGEMA_signal_8998) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M16), .A0_f (new_AGEMA_signal_8717), .A1_t (new_AGEMA_signal_8718), .A1_f (new_AGEMA_signal_8719), .B0_t (SubBytesIns_Inst_Sbox_1_M13), .B0_f (new_AGEMA_signal_8252), .B1_t (new_AGEMA_signal_8253), .B1_f (new_AGEMA_signal_8254), .Z0_t (SubBytesIns_Inst_Sbox_1_M20), .Z0_f (new_AGEMA_signal_8999), .Z1_t (new_AGEMA_signal_9000), .Z1_f (new_AGEMA_signal_9001) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M17), .A0_f (new_AGEMA_signal_8720), .A1_t (new_AGEMA_signal_8721), .A1_f (new_AGEMA_signal_8722), .B0_t (SubBytesIns_Inst_Sbox_1_M15), .B0_f (new_AGEMA_signal_8714), .B1_t (new_AGEMA_signal_8715), .B1_f (new_AGEMA_signal_8716), .Z0_t (SubBytesIns_Inst_Sbox_1_M21), .Z0_f (new_AGEMA_signal_9002), .Z1_t (new_AGEMA_signal_9003), .Z1_f (new_AGEMA_signal_9004) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M18), .A0_f (new_AGEMA_signal_8723), .A1_t (new_AGEMA_signal_8724), .A1_f (new_AGEMA_signal_8725), .B0_t (SubBytesIns_Inst_Sbox_1_M13), .B0_f (new_AGEMA_signal_8252), .B1_t (new_AGEMA_signal_8253), .B1_f (new_AGEMA_signal_8254), .Z0_t (SubBytesIns_Inst_Sbox_1_M22), .Z0_f (new_AGEMA_signal_9005), .Z1_t (new_AGEMA_signal_9006), .Z1_f (new_AGEMA_signal_9007) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M19), .A0_f (new_AGEMA_signal_8996), .A1_t (new_AGEMA_signal_8997), .A1_f (new_AGEMA_signal_8998), .B0_t (SubBytesIns_Inst_Sbox_1_T25), .B0_f (new_AGEMA_signal_8234), .B1_t (new_AGEMA_signal_8235), .B1_f (new_AGEMA_signal_8236), .Z0_t (SubBytesIns_Inst_Sbox_1_M23), .Z0_f (new_AGEMA_signal_9236), .Z1_t (new_AGEMA_signal_9237), .Z1_f (new_AGEMA_signal_9238) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M22), .A0_f (new_AGEMA_signal_9005), .A1_t (new_AGEMA_signal_9006), .A1_f (new_AGEMA_signal_9007), .B0_t (SubBytesIns_Inst_Sbox_1_M23), .B0_f (new_AGEMA_signal_9236), .B1_t (new_AGEMA_signal_9237), .B1_f (new_AGEMA_signal_9238), .Z0_t (SubBytesIns_Inst_Sbox_1_M24), .Z0_f (new_AGEMA_signal_9491), .Z1_t (new_AGEMA_signal_9492), .Z1_f (new_AGEMA_signal_9493) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M22), .A0_f (new_AGEMA_signal_9005), .A1_t (new_AGEMA_signal_9006), .A1_f (new_AGEMA_signal_9007), .B0_t (SubBytesIns_Inst_Sbox_1_M20), .B0_f (new_AGEMA_signal_8999), .B1_t (new_AGEMA_signal_9000), .B1_f (new_AGEMA_signal_9001), .Z0_t (SubBytesIns_Inst_Sbox_1_M25), .Z0_f (new_AGEMA_signal_9239), .Z1_t (new_AGEMA_signal_9240), .Z1_f (new_AGEMA_signal_9241) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M21), .A0_f (new_AGEMA_signal_9002), .A1_t (new_AGEMA_signal_9003), .A1_f (new_AGEMA_signal_9004), .B0_t (SubBytesIns_Inst_Sbox_1_M25), .B0_f (new_AGEMA_signal_9239), .B1_t (new_AGEMA_signal_9240), .B1_f (new_AGEMA_signal_9241), .Z0_t (SubBytesIns_Inst_Sbox_1_M26), .Z0_f (new_AGEMA_signal_9494), .Z1_t (new_AGEMA_signal_9495), .Z1_f (new_AGEMA_signal_9496) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M20), .A0_f (new_AGEMA_signal_8999), .A1_t (new_AGEMA_signal_9000), .A1_f (new_AGEMA_signal_9001), .B0_t (SubBytesIns_Inst_Sbox_1_M21), .B0_f (new_AGEMA_signal_9002), .B1_t (new_AGEMA_signal_9003), .B1_f (new_AGEMA_signal_9004), .Z0_t (SubBytesIns_Inst_Sbox_1_M27), .Z0_f (new_AGEMA_signal_9242), .Z1_t (new_AGEMA_signal_9243), .Z1_f (new_AGEMA_signal_9244) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M23), .A0_f (new_AGEMA_signal_9236), .A1_t (new_AGEMA_signal_9237), .A1_f (new_AGEMA_signal_9238), .B0_t (SubBytesIns_Inst_Sbox_1_M25), .B0_f (new_AGEMA_signal_9239), .B1_t (new_AGEMA_signal_9240), .B1_f (new_AGEMA_signal_9241), .Z0_t (SubBytesIns_Inst_Sbox_1_M28), .Z0_f (new_AGEMA_signal_9497), .Z1_t (new_AGEMA_signal_9498), .Z1_f (new_AGEMA_signal_9499) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M28), .A0_f (new_AGEMA_signal_9497), .A1_t (new_AGEMA_signal_9498), .A1_f (new_AGEMA_signal_9499), .B0_t (SubBytesIns_Inst_Sbox_1_M27), .B0_f (new_AGEMA_signal_9242), .B1_t (new_AGEMA_signal_9243), .B1_f (new_AGEMA_signal_9244), .Z0_t (SubBytesIns_Inst_Sbox_1_M29), .Z0_f (new_AGEMA_signal_9791), .Z1_t (new_AGEMA_signal_9792), .Z1_f (new_AGEMA_signal_9793) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M26), .A0_f (new_AGEMA_signal_9494), .A1_t (new_AGEMA_signal_9495), .A1_f (new_AGEMA_signal_9496), .B0_t (SubBytesIns_Inst_Sbox_1_M24), .B0_f (new_AGEMA_signal_9491), .B1_t (new_AGEMA_signal_9492), .B1_f (new_AGEMA_signal_9493), .Z0_t (SubBytesIns_Inst_Sbox_1_M30), .Z0_f (new_AGEMA_signal_9794), .Z1_t (new_AGEMA_signal_9795), .Z1_f (new_AGEMA_signal_9796) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M20), .A0_f (new_AGEMA_signal_8999), .A1_t (new_AGEMA_signal_9000), .A1_f (new_AGEMA_signal_9001), .B0_t (SubBytesIns_Inst_Sbox_1_M23), .B0_f (new_AGEMA_signal_9236), .B1_t (new_AGEMA_signal_9237), .B1_f (new_AGEMA_signal_9238), .Z0_t (SubBytesIns_Inst_Sbox_1_M31), .Z0_f (new_AGEMA_signal_9500), .Z1_t (new_AGEMA_signal_9501), .Z1_f (new_AGEMA_signal_9502) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M27), .A0_f (new_AGEMA_signal_9242), .A1_t (new_AGEMA_signal_9243), .A1_f (new_AGEMA_signal_9244), .B0_t (SubBytesIns_Inst_Sbox_1_M31), .B0_f (new_AGEMA_signal_9500), .B1_t (new_AGEMA_signal_9501), .B1_f (new_AGEMA_signal_9502), .Z0_t (SubBytesIns_Inst_Sbox_1_M32), .Z0_f (new_AGEMA_signal_9797), .Z1_t (new_AGEMA_signal_9798), .Z1_f (new_AGEMA_signal_9799) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M27), .A0_f (new_AGEMA_signal_9242), .A1_t (new_AGEMA_signal_9243), .A1_f (new_AGEMA_signal_9244), .B0_t (SubBytesIns_Inst_Sbox_1_M25), .B0_f (new_AGEMA_signal_9239), .B1_t (new_AGEMA_signal_9240), .B1_f (new_AGEMA_signal_9241), .Z0_t (SubBytesIns_Inst_Sbox_1_M33), .Z0_f (new_AGEMA_signal_9503), .Z1_t (new_AGEMA_signal_9504), .Z1_f (new_AGEMA_signal_9505) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M21), .A0_f (new_AGEMA_signal_9002), .A1_t (new_AGEMA_signal_9003), .A1_f (new_AGEMA_signal_9004), .B0_t (SubBytesIns_Inst_Sbox_1_M22), .B0_f (new_AGEMA_signal_9005), .B1_t (new_AGEMA_signal_9006), .B1_f (new_AGEMA_signal_9007), .Z0_t (SubBytesIns_Inst_Sbox_1_M34), .Z0_f (new_AGEMA_signal_9245), .Z1_t (new_AGEMA_signal_9246), .Z1_f (new_AGEMA_signal_9247) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M24), .A0_f (new_AGEMA_signal_9491), .A1_t (new_AGEMA_signal_9492), .A1_f (new_AGEMA_signal_9493), .B0_t (SubBytesIns_Inst_Sbox_1_M34), .B0_f (new_AGEMA_signal_9245), .B1_t (new_AGEMA_signal_9246), .B1_f (new_AGEMA_signal_9247), .Z0_t (SubBytesIns_Inst_Sbox_1_M35), .Z0_f (new_AGEMA_signal_9800), .Z1_t (new_AGEMA_signal_9801), .Z1_f (new_AGEMA_signal_9802) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M24), .A0_f (new_AGEMA_signal_9491), .A1_t (new_AGEMA_signal_9492), .A1_f (new_AGEMA_signal_9493), .B0_t (SubBytesIns_Inst_Sbox_1_M25), .B0_f (new_AGEMA_signal_9239), .B1_t (new_AGEMA_signal_9240), .B1_f (new_AGEMA_signal_9241), .Z0_t (SubBytesIns_Inst_Sbox_1_M36), .Z0_f (new_AGEMA_signal_9803), .Z1_t (new_AGEMA_signal_9804), .Z1_f (new_AGEMA_signal_9805) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M21), .A0_f (new_AGEMA_signal_9002), .A1_t (new_AGEMA_signal_9003), .A1_f (new_AGEMA_signal_9004), .B0_t (SubBytesIns_Inst_Sbox_1_M29), .B0_f (new_AGEMA_signal_9791), .B1_t (new_AGEMA_signal_9792), .B1_f (new_AGEMA_signal_9793), .Z0_t (SubBytesIns_Inst_Sbox_1_M37), .Z0_f (new_AGEMA_signal_10076), .Z1_t (new_AGEMA_signal_10077), .Z1_f (new_AGEMA_signal_10078) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M32), .A0_f (new_AGEMA_signal_9797), .A1_t (new_AGEMA_signal_9798), .A1_f (new_AGEMA_signal_9799), .B0_t (SubBytesIns_Inst_Sbox_1_M33), .B0_f (new_AGEMA_signal_9503), .B1_t (new_AGEMA_signal_9504), .B1_f (new_AGEMA_signal_9505), .Z0_t (SubBytesIns_Inst_Sbox_1_M38), .Z0_f (new_AGEMA_signal_10079), .Z1_t (new_AGEMA_signal_10080), .Z1_f (new_AGEMA_signal_10081) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M23), .A0_f (new_AGEMA_signal_9236), .A1_t (new_AGEMA_signal_9237), .A1_f (new_AGEMA_signal_9238), .B0_t (SubBytesIns_Inst_Sbox_1_M30), .B0_f (new_AGEMA_signal_9794), .B1_t (new_AGEMA_signal_9795), .B1_f (new_AGEMA_signal_9796), .Z0_t (SubBytesIns_Inst_Sbox_1_M39), .Z0_f (new_AGEMA_signal_10082), .Z1_t (new_AGEMA_signal_10083), .Z1_f (new_AGEMA_signal_10084) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M35), .A0_f (new_AGEMA_signal_9800), .A1_t (new_AGEMA_signal_9801), .A1_f (new_AGEMA_signal_9802), .B0_t (SubBytesIns_Inst_Sbox_1_M36), .B0_f (new_AGEMA_signal_9803), .B1_t (new_AGEMA_signal_9804), .B1_f (new_AGEMA_signal_9805), .Z0_t (SubBytesIns_Inst_Sbox_1_M40), .Z0_f (new_AGEMA_signal_10085), .Z1_t (new_AGEMA_signal_10086), .Z1_f (new_AGEMA_signal_10087) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M38), .A0_f (new_AGEMA_signal_10079), .A1_t (new_AGEMA_signal_10080), .A1_f (new_AGEMA_signal_10081), .B0_t (SubBytesIns_Inst_Sbox_1_M40), .B0_f (new_AGEMA_signal_10085), .B1_t (new_AGEMA_signal_10086), .B1_f (new_AGEMA_signal_10087), .Z0_t (SubBytesIns_Inst_Sbox_1_M41), .Z0_f (new_AGEMA_signal_10436), .Z1_t (new_AGEMA_signal_10437), .Z1_f (new_AGEMA_signal_10438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M37), .A0_f (new_AGEMA_signal_10076), .A1_t (new_AGEMA_signal_10077), .A1_f (new_AGEMA_signal_10078), .B0_t (SubBytesIns_Inst_Sbox_1_M39), .B0_f (new_AGEMA_signal_10082), .B1_t (new_AGEMA_signal_10083), .B1_f (new_AGEMA_signal_10084), .Z0_t (SubBytesIns_Inst_Sbox_1_M42), .Z0_f (new_AGEMA_signal_10439), .Z1_t (new_AGEMA_signal_10440), .Z1_f (new_AGEMA_signal_10441) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M37), .A0_f (new_AGEMA_signal_10076), .A1_t (new_AGEMA_signal_10077), .A1_f (new_AGEMA_signal_10078), .B0_t (SubBytesIns_Inst_Sbox_1_M38), .B0_f (new_AGEMA_signal_10079), .B1_t (new_AGEMA_signal_10080), .B1_f (new_AGEMA_signal_10081), .Z0_t (SubBytesIns_Inst_Sbox_1_M43), .Z0_f (new_AGEMA_signal_10442), .Z1_t (new_AGEMA_signal_10443), .Z1_f (new_AGEMA_signal_10444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M39), .A0_f (new_AGEMA_signal_10082), .A1_t (new_AGEMA_signal_10083), .A1_f (new_AGEMA_signal_10084), .B0_t (SubBytesIns_Inst_Sbox_1_M40), .B0_f (new_AGEMA_signal_10085), .B1_t (new_AGEMA_signal_10086), .B1_f (new_AGEMA_signal_10087), .Z0_t (SubBytesIns_Inst_Sbox_1_M44), .Z0_f (new_AGEMA_signal_10445), .Z1_t (new_AGEMA_signal_10446), .Z1_f (new_AGEMA_signal_10447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M42), .A0_f (new_AGEMA_signal_10439), .A1_t (new_AGEMA_signal_10440), .A1_f (new_AGEMA_signal_10441), .B0_t (SubBytesIns_Inst_Sbox_1_M41), .B0_f (new_AGEMA_signal_10436), .B1_t (new_AGEMA_signal_10437), .B1_f (new_AGEMA_signal_10438), .Z0_t (SubBytesIns_Inst_Sbox_1_M45), .Z0_f (new_AGEMA_signal_11156), .Z1_t (new_AGEMA_signal_11157), .Z1_f (new_AGEMA_signal_11158) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M44), .A0_f (new_AGEMA_signal_10445), .A1_t (new_AGEMA_signal_10446), .A1_f (new_AGEMA_signal_10447), .B0_t (SubBytesIns_Inst_Sbox_1_T6), .B0_f (new_AGEMA_signal_6952), .B1_t (new_AGEMA_signal_6953), .B1_f (new_AGEMA_signal_6954), .Z0_t (SubBytesIns_Inst_Sbox_1_M46), .Z0_f (new_AGEMA_signal_11159), .Z1_t (new_AGEMA_signal_11160), .Z1_f (new_AGEMA_signal_11161) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M40), .A0_f (new_AGEMA_signal_10085), .A1_t (new_AGEMA_signal_10086), .A1_f (new_AGEMA_signal_10087), .B0_t (SubBytesIns_Inst_Sbox_1_T8), .B0_f (new_AGEMA_signal_7511), .B1_t (new_AGEMA_signal_7512), .B1_f (new_AGEMA_signal_7513), .Z0_t (SubBytesIns_Inst_Sbox_1_M47), .Z0_f (new_AGEMA_signal_10448), .Z1_t (new_AGEMA_signal_10449), .Z1_f (new_AGEMA_signal_10450) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M39), .A0_f (new_AGEMA_signal_10082), .A1_t (new_AGEMA_signal_10083), .A1_f (new_AGEMA_signal_10084), .B0_t (ciphertext_s0_t[8]), .B0_f (ciphertext_s0_f[8]), .B1_t (ciphertext_s1_t[8]), .B1_f (ciphertext_s1_f[8]), .Z0_t (SubBytesIns_Inst_Sbox_1_M48), .Z0_f (new_AGEMA_signal_10451), .Z1_t (new_AGEMA_signal_10452), .Z1_f (new_AGEMA_signal_10453) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M43), .A0_f (new_AGEMA_signal_10442), .A1_t (new_AGEMA_signal_10443), .A1_f (new_AGEMA_signal_10444), .B0_t (SubBytesIns_Inst_Sbox_1_T16), .B0_f (new_AGEMA_signal_6964), .B1_t (new_AGEMA_signal_6965), .B1_f (new_AGEMA_signal_6966), .Z0_t (SubBytesIns_Inst_Sbox_1_M49), .Z0_f (new_AGEMA_signal_11162), .Z1_t (new_AGEMA_signal_11163), .Z1_f (new_AGEMA_signal_11164) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M38), .A0_f (new_AGEMA_signal_10079), .A1_t (new_AGEMA_signal_10080), .A1_f (new_AGEMA_signal_10081), .B0_t (SubBytesIns_Inst_Sbox_1_T9), .B0_f (new_AGEMA_signal_6955), .B1_t (new_AGEMA_signal_6956), .B1_f (new_AGEMA_signal_6957), .Z0_t (SubBytesIns_Inst_Sbox_1_M50), .Z0_f (new_AGEMA_signal_10454), .Z1_t (new_AGEMA_signal_10455), .Z1_f (new_AGEMA_signal_10456) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M37), .A0_f (new_AGEMA_signal_10076), .A1_t (new_AGEMA_signal_10077), .A1_f (new_AGEMA_signal_10078), .B0_t (SubBytesIns_Inst_Sbox_1_T17), .B0_f (new_AGEMA_signal_7520), .B1_t (new_AGEMA_signal_7521), .B1_f (new_AGEMA_signal_7522), .Z0_t (SubBytesIns_Inst_Sbox_1_M51), .Z0_f (new_AGEMA_signal_10457), .Z1_t (new_AGEMA_signal_10458), .Z1_f (new_AGEMA_signal_10459) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M42), .A0_f (new_AGEMA_signal_10439), .A1_t (new_AGEMA_signal_10440), .A1_f (new_AGEMA_signal_10441), .B0_t (SubBytesIns_Inst_Sbox_1_T15), .B0_f (new_AGEMA_signal_6961), .B1_t (new_AGEMA_signal_6962), .B1_f (new_AGEMA_signal_6963), .Z0_t (SubBytesIns_Inst_Sbox_1_M52), .Z0_f (new_AGEMA_signal_11165), .Z1_t (new_AGEMA_signal_11166), .Z1_f (new_AGEMA_signal_11167) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M45), .A0_f (new_AGEMA_signal_11156), .A1_t (new_AGEMA_signal_11157), .A1_f (new_AGEMA_signal_11158), .B0_t (SubBytesIns_Inst_Sbox_1_T27), .B0_f (new_AGEMA_signal_6973), .B1_t (new_AGEMA_signal_6974), .B1_f (new_AGEMA_signal_6975), .Z0_t (SubBytesIns_Inst_Sbox_1_M53), .Z0_f (new_AGEMA_signal_11846), .Z1_t (new_AGEMA_signal_11847), .Z1_f (new_AGEMA_signal_11848) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M41), .A0_f (new_AGEMA_signal_10436), .A1_t (new_AGEMA_signal_10437), .A1_f (new_AGEMA_signal_10438), .B0_t (SubBytesIns_Inst_Sbox_1_T10), .B0_f (new_AGEMA_signal_7514), .B1_t (new_AGEMA_signal_7515), .B1_f (new_AGEMA_signal_7516), .Z0_t (SubBytesIns_Inst_Sbox_1_M54), .Z0_f (new_AGEMA_signal_11168), .Z1_t (new_AGEMA_signal_11169), .Z1_f (new_AGEMA_signal_11170) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M44), .A0_f (new_AGEMA_signal_10445), .A1_t (new_AGEMA_signal_10446), .A1_f (new_AGEMA_signal_10447), .B0_t (SubBytesIns_Inst_Sbox_1_T13), .B0_f (new_AGEMA_signal_6958), .B1_t (new_AGEMA_signal_6959), .B1_f (new_AGEMA_signal_6960), .Z0_t (SubBytesIns_Inst_Sbox_1_M55), .Z0_f (new_AGEMA_signal_11171), .Z1_t (new_AGEMA_signal_11172), .Z1_f (new_AGEMA_signal_11173) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M40), .A0_f (new_AGEMA_signal_10085), .A1_t (new_AGEMA_signal_10086), .A1_f (new_AGEMA_signal_10087), .B0_t (SubBytesIns_Inst_Sbox_1_T23), .B0_f (new_AGEMA_signal_7526), .B1_t (new_AGEMA_signal_7527), .B1_f (new_AGEMA_signal_7528), .Z0_t (SubBytesIns_Inst_Sbox_1_M56), .Z0_f (new_AGEMA_signal_10460), .Z1_t (new_AGEMA_signal_10461), .Z1_f (new_AGEMA_signal_10462) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M39), .A0_f (new_AGEMA_signal_10082), .A1_t (new_AGEMA_signal_10083), .A1_f (new_AGEMA_signal_10084), .B0_t (SubBytesIns_Inst_Sbox_1_T19), .B0_f (new_AGEMA_signal_6967), .B1_t (new_AGEMA_signal_6968), .B1_f (new_AGEMA_signal_6969), .Z0_t (SubBytesIns_Inst_Sbox_1_M57), .Z0_f (new_AGEMA_signal_10463), .Z1_t (new_AGEMA_signal_10464), .Z1_f (new_AGEMA_signal_10465) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M43), .A0_f (new_AGEMA_signal_10442), .A1_t (new_AGEMA_signal_10443), .A1_f (new_AGEMA_signal_10444), .B0_t (SubBytesIns_Inst_Sbox_1_T3), .B0_f (new_AGEMA_signal_6382), .B1_t (new_AGEMA_signal_6383), .B1_f (new_AGEMA_signal_6384), .Z0_t (SubBytesIns_Inst_Sbox_1_M58), .Z0_f (new_AGEMA_signal_11174), .Z1_t (new_AGEMA_signal_11175), .Z1_f (new_AGEMA_signal_11176) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M38), .A0_f (new_AGEMA_signal_10079), .A1_t (new_AGEMA_signal_10080), .A1_f (new_AGEMA_signal_10081), .B0_t (SubBytesIns_Inst_Sbox_1_T22), .B0_f (new_AGEMA_signal_6970), .B1_t (new_AGEMA_signal_6971), .B1_f (new_AGEMA_signal_6972), .Z0_t (SubBytesIns_Inst_Sbox_1_M59), .Z0_f (new_AGEMA_signal_10466), .Z1_t (new_AGEMA_signal_10467), .Z1_f (new_AGEMA_signal_10468) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M37), .A0_f (new_AGEMA_signal_10076), .A1_t (new_AGEMA_signal_10077), .A1_f (new_AGEMA_signal_10078), .B0_t (SubBytesIns_Inst_Sbox_1_T20), .B0_f (new_AGEMA_signal_7523), .B1_t (new_AGEMA_signal_7524), .B1_f (new_AGEMA_signal_7525), .Z0_t (SubBytesIns_Inst_Sbox_1_M60), .Z0_f (new_AGEMA_signal_10469), .Z1_t (new_AGEMA_signal_10470), .Z1_f (new_AGEMA_signal_10471) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M42), .A0_f (new_AGEMA_signal_10439), .A1_t (new_AGEMA_signal_10440), .A1_f (new_AGEMA_signal_10441), .B0_t (SubBytesIns_Inst_Sbox_1_T1), .B0_f (new_AGEMA_signal_6376), .B1_t (new_AGEMA_signal_6377), .B1_f (new_AGEMA_signal_6378), .Z0_t (SubBytesIns_Inst_Sbox_1_M61), .Z0_f (new_AGEMA_signal_11177), .Z1_t (new_AGEMA_signal_11178), .Z1_f (new_AGEMA_signal_11179) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M45), .A0_f (new_AGEMA_signal_11156), .A1_t (new_AGEMA_signal_11157), .A1_f (new_AGEMA_signal_11158), .B0_t (SubBytesIns_Inst_Sbox_1_T4), .B0_f (new_AGEMA_signal_6385), .B1_t (new_AGEMA_signal_6386), .B1_f (new_AGEMA_signal_6387), .Z0_t (SubBytesIns_Inst_Sbox_1_M62), .Z0_f (new_AGEMA_signal_11849), .Z1_t (new_AGEMA_signal_11850), .Z1_f (new_AGEMA_signal_11851) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M41), .A0_f (new_AGEMA_signal_10436), .A1_t (new_AGEMA_signal_10437), .A1_f (new_AGEMA_signal_10438), .B0_t (SubBytesIns_Inst_Sbox_1_T2), .B0_f (new_AGEMA_signal_6379), .B1_t (new_AGEMA_signal_6380), .B1_f (new_AGEMA_signal_6381), .Z0_t (SubBytesIns_Inst_Sbox_1_M63), .Z0_f (new_AGEMA_signal_11180), .Z1_t (new_AGEMA_signal_11181), .Z1_f (new_AGEMA_signal_11182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M61), .A0_f (new_AGEMA_signal_11177), .A1_t (new_AGEMA_signal_11178), .A1_f (new_AGEMA_signal_11179), .B0_t (SubBytesIns_Inst_Sbox_1_M62), .B0_f (new_AGEMA_signal_11849), .B1_t (new_AGEMA_signal_11850), .B1_f (new_AGEMA_signal_11851), .Z0_t (SubBytesIns_Inst_Sbox_1_L0), .Z0_f (new_AGEMA_signal_12431), .Z1_t (new_AGEMA_signal_12432), .Z1_f (new_AGEMA_signal_12433) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M50), .A0_f (new_AGEMA_signal_10454), .A1_t (new_AGEMA_signal_10455), .A1_f (new_AGEMA_signal_10456), .B0_t (SubBytesIns_Inst_Sbox_1_M56), .B0_f (new_AGEMA_signal_10460), .B1_t (new_AGEMA_signal_10461), .B1_f (new_AGEMA_signal_10462), .Z0_t (SubBytesIns_Inst_Sbox_1_L1), .Z0_f (new_AGEMA_signal_11183), .Z1_t (new_AGEMA_signal_11184), .Z1_f (new_AGEMA_signal_11185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M46), .A0_f (new_AGEMA_signal_11159), .A1_t (new_AGEMA_signal_11160), .A1_f (new_AGEMA_signal_11161), .B0_t (SubBytesIns_Inst_Sbox_1_M48), .B0_f (new_AGEMA_signal_10451), .B1_t (new_AGEMA_signal_10452), .B1_f (new_AGEMA_signal_10453), .Z0_t (SubBytesIns_Inst_Sbox_1_L2), .Z0_f (new_AGEMA_signal_11852), .Z1_t (new_AGEMA_signal_11853), .Z1_f (new_AGEMA_signal_11854) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M47), .A0_f (new_AGEMA_signal_10448), .A1_t (new_AGEMA_signal_10449), .A1_f (new_AGEMA_signal_10450), .B0_t (SubBytesIns_Inst_Sbox_1_M55), .B0_f (new_AGEMA_signal_11171), .B1_t (new_AGEMA_signal_11172), .B1_f (new_AGEMA_signal_11173), .Z0_t (SubBytesIns_Inst_Sbox_1_L3), .Z0_f (new_AGEMA_signal_11855), .Z1_t (new_AGEMA_signal_11856), .Z1_f (new_AGEMA_signal_11857) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M54), .A0_f (new_AGEMA_signal_11168), .A1_t (new_AGEMA_signal_11169), .A1_f (new_AGEMA_signal_11170), .B0_t (SubBytesIns_Inst_Sbox_1_M58), .B0_f (new_AGEMA_signal_11174), .B1_t (new_AGEMA_signal_11175), .B1_f (new_AGEMA_signal_11176), .Z0_t (SubBytesIns_Inst_Sbox_1_L4), .Z0_f (new_AGEMA_signal_11858), .Z1_t (new_AGEMA_signal_11859), .Z1_f (new_AGEMA_signal_11860) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M49), .A0_f (new_AGEMA_signal_11162), .A1_t (new_AGEMA_signal_11163), .A1_f (new_AGEMA_signal_11164), .B0_t (SubBytesIns_Inst_Sbox_1_M61), .B0_f (new_AGEMA_signal_11177), .B1_t (new_AGEMA_signal_11178), .B1_f (new_AGEMA_signal_11179), .Z0_t (SubBytesIns_Inst_Sbox_1_L5), .Z0_f (new_AGEMA_signal_11861), .Z1_t (new_AGEMA_signal_11862), .Z1_f (new_AGEMA_signal_11863) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M62), .A0_f (new_AGEMA_signal_11849), .A1_t (new_AGEMA_signal_11850), .A1_f (new_AGEMA_signal_11851), .B0_t (SubBytesIns_Inst_Sbox_1_L5), .B0_f (new_AGEMA_signal_11861), .B1_t (new_AGEMA_signal_11862), .B1_f (new_AGEMA_signal_11863), .Z0_t (SubBytesIns_Inst_Sbox_1_L6), .Z0_f (new_AGEMA_signal_12434), .Z1_t (new_AGEMA_signal_12435), .Z1_f (new_AGEMA_signal_12436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M46), .A0_f (new_AGEMA_signal_11159), .A1_t (new_AGEMA_signal_11160), .A1_f (new_AGEMA_signal_11161), .B0_t (SubBytesIns_Inst_Sbox_1_L3), .B0_f (new_AGEMA_signal_11855), .B1_t (new_AGEMA_signal_11856), .B1_f (new_AGEMA_signal_11857), .Z0_t (SubBytesIns_Inst_Sbox_1_L7), .Z0_f (new_AGEMA_signal_12437), .Z1_t (new_AGEMA_signal_12438), .Z1_f (new_AGEMA_signal_12439) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M51), .A0_f (new_AGEMA_signal_10457), .A1_t (new_AGEMA_signal_10458), .A1_f (new_AGEMA_signal_10459), .B0_t (SubBytesIns_Inst_Sbox_1_M59), .B0_f (new_AGEMA_signal_10466), .B1_t (new_AGEMA_signal_10467), .B1_f (new_AGEMA_signal_10468), .Z0_t (SubBytesIns_Inst_Sbox_1_L8), .Z0_f (new_AGEMA_signal_11186), .Z1_t (new_AGEMA_signal_11187), .Z1_f (new_AGEMA_signal_11188) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M52), .A0_f (new_AGEMA_signal_11165), .A1_t (new_AGEMA_signal_11166), .A1_f (new_AGEMA_signal_11167), .B0_t (SubBytesIns_Inst_Sbox_1_M53), .B0_f (new_AGEMA_signal_11846), .B1_t (new_AGEMA_signal_11847), .B1_f (new_AGEMA_signal_11848), .Z0_t (SubBytesIns_Inst_Sbox_1_L9), .Z0_f (new_AGEMA_signal_12440), .Z1_t (new_AGEMA_signal_12441), .Z1_f (new_AGEMA_signal_12442) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M53), .A0_f (new_AGEMA_signal_11846), .A1_t (new_AGEMA_signal_11847), .A1_f (new_AGEMA_signal_11848), .B0_t (SubBytesIns_Inst_Sbox_1_L4), .B0_f (new_AGEMA_signal_11858), .B1_t (new_AGEMA_signal_11859), .B1_f (new_AGEMA_signal_11860), .Z0_t (SubBytesIns_Inst_Sbox_1_L10), .Z0_f (new_AGEMA_signal_12443), .Z1_t (new_AGEMA_signal_12444), .Z1_f (new_AGEMA_signal_12445) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M60), .A0_f (new_AGEMA_signal_10469), .A1_t (new_AGEMA_signal_10470), .A1_f (new_AGEMA_signal_10471), .B0_t (SubBytesIns_Inst_Sbox_1_L2), .B0_f (new_AGEMA_signal_11852), .B1_t (new_AGEMA_signal_11853), .B1_f (new_AGEMA_signal_11854), .Z0_t (SubBytesIns_Inst_Sbox_1_L11), .Z0_f (new_AGEMA_signal_12446), .Z1_t (new_AGEMA_signal_12447), .Z1_f (new_AGEMA_signal_12448) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M48), .A0_f (new_AGEMA_signal_10451), .A1_t (new_AGEMA_signal_10452), .A1_f (new_AGEMA_signal_10453), .B0_t (SubBytesIns_Inst_Sbox_1_M51), .B0_f (new_AGEMA_signal_10457), .B1_t (new_AGEMA_signal_10458), .B1_f (new_AGEMA_signal_10459), .Z0_t (SubBytesIns_Inst_Sbox_1_L12), .Z0_f (new_AGEMA_signal_11189), .Z1_t (new_AGEMA_signal_11190), .Z1_f (new_AGEMA_signal_11191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M50), .A0_f (new_AGEMA_signal_10454), .A1_t (new_AGEMA_signal_10455), .A1_f (new_AGEMA_signal_10456), .B0_t (SubBytesIns_Inst_Sbox_1_L0), .B0_f (new_AGEMA_signal_12431), .B1_t (new_AGEMA_signal_12432), .B1_f (new_AGEMA_signal_12433), .Z0_t (SubBytesIns_Inst_Sbox_1_L13), .Z0_f (new_AGEMA_signal_13001), .Z1_t (new_AGEMA_signal_13002), .Z1_f (new_AGEMA_signal_13003) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M52), .A0_f (new_AGEMA_signal_11165), .A1_t (new_AGEMA_signal_11166), .A1_f (new_AGEMA_signal_11167), .B0_t (SubBytesIns_Inst_Sbox_1_M61), .B0_f (new_AGEMA_signal_11177), .B1_t (new_AGEMA_signal_11178), .B1_f (new_AGEMA_signal_11179), .Z0_t (SubBytesIns_Inst_Sbox_1_L14), .Z0_f (new_AGEMA_signal_11864), .Z1_t (new_AGEMA_signal_11865), .Z1_f (new_AGEMA_signal_11866) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M55), .A0_f (new_AGEMA_signal_11171), .A1_t (new_AGEMA_signal_11172), .A1_f (new_AGEMA_signal_11173), .B0_t (SubBytesIns_Inst_Sbox_1_L1), .B0_f (new_AGEMA_signal_11183), .B1_t (new_AGEMA_signal_11184), .B1_f (new_AGEMA_signal_11185), .Z0_t (SubBytesIns_Inst_Sbox_1_L15), .Z0_f (new_AGEMA_signal_11867), .Z1_t (new_AGEMA_signal_11868), .Z1_f (new_AGEMA_signal_11869) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M56), .A0_f (new_AGEMA_signal_10460), .A1_t (new_AGEMA_signal_10461), .A1_f (new_AGEMA_signal_10462), .B0_t (SubBytesIns_Inst_Sbox_1_L0), .B0_f (new_AGEMA_signal_12431), .B1_t (new_AGEMA_signal_12432), .B1_f (new_AGEMA_signal_12433), .Z0_t (SubBytesIns_Inst_Sbox_1_L16), .Z0_f (new_AGEMA_signal_13004), .Z1_t (new_AGEMA_signal_13005), .Z1_f (new_AGEMA_signal_13006) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M57), .A0_f (new_AGEMA_signal_10463), .A1_t (new_AGEMA_signal_10464), .A1_f (new_AGEMA_signal_10465), .B0_t (SubBytesIns_Inst_Sbox_1_L1), .B0_f (new_AGEMA_signal_11183), .B1_t (new_AGEMA_signal_11184), .B1_f (new_AGEMA_signal_11185), .Z0_t (SubBytesIns_Inst_Sbox_1_L17), .Z0_f (new_AGEMA_signal_11870), .Z1_t (new_AGEMA_signal_11871), .Z1_f (new_AGEMA_signal_11872) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M58), .A0_f (new_AGEMA_signal_11174), .A1_t (new_AGEMA_signal_11175), .A1_f (new_AGEMA_signal_11176), .B0_t (SubBytesIns_Inst_Sbox_1_L8), .B0_f (new_AGEMA_signal_11186), .B1_t (new_AGEMA_signal_11187), .B1_f (new_AGEMA_signal_11188), .Z0_t (SubBytesIns_Inst_Sbox_1_L18), .Z0_f (new_AGEMA_signal_11873), .Z1_t (new_AGEMA_signal_11874), .Z1_f (new_AGEMA_signal_11875) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M63), .A0_f (new_AGEMA_signal_11180), .A1_t (new_AGEMA_signal_11181), .A1_f (new_AGEMA_signal_11182), .B0_t (SubBytesIns_Inst_Sbox_1_L4), .B0_f (new_AGEMA_signal_11858), .B1_t (new_AGEMA_signal_11859), .B1_f (new_AGEMA_signal_11860), .Z0_t (SubBytesIns_Inst_Sbox_1_L19), .Z0_f (new_AGEMA_signal_12449), .Z1_t (new_AGEMA_signal_12450), .Z1_f (new_AGEMA_signal_12451) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L0), .A0_f (new_AGEMA_signal_12431), .A1_t (new_AGEMA_signal_12432), .A1_f (new_AGEMA_signal_12433), .B0_t (SubBytesIns_Inst_Sbox_1_L1), .B0_f (new_AGEMA_signal_11183), .B1_t (new_AGEMA_signal_11184), .B1_f (new_AGEMA_signal_11185), .Z0_t (SubBytesIns_Inst_Sbox_1_L20), .Z0_f (new_AGEMA_signal_13007), .Z1_t (new_AGEMA_signal_13008), .Z1_f (new_AGEMA_signal_13009) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L1), .A0_f (new_AGEMA_signal_11183), .A1_t (new_AGEMA_signal_11184), .A1_f (new_AGEMA_signal_11185), .B0_t (SubBytesIns_Inst_Sbox_1_L7), .B0_f (new_AGEMA_signal_12437), .B1_t (new_AGEMA_signal_12438), .B1_f (new_AGEMA_signal_12439), .Z0_t (SubBytesIns_Inst_Sbox_1_L21), .Z0_f (new_AGEMA_signal_13010), .Z1_t (new_AGEMA_signal_13011), .Z1_f (new_AGEMA_signal_13012) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L3), .A0_f (new_AGEMA_signal_11855), .A1_t (new_AGEMA_signal_11856), .A1_f (new_AGEMA_signal_11857), .B0_t (SubBytesIns_Inst_Sbox_1_L12), .B0_f (new_AGEMA_signal_11189), .B1_t (new_AGEMA_signal_11190), .B1_f (new_AGEMA_signal_11191), .Z0_t (SubBytesIns_Inst_Sbox_1_L22), .Z0_f (new_AGEMA_signal_12452), .Z1_t (new_AGEMA_signal_12453), .Z1_f (new_AGEMA_signal_12454) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L18), .A0_f (new_AGEMA_signal_11873), .A1_t (new_AGEMA_signal_11874), .A1_f (new_AGEMA_signal_11875), .B0_t (SubBytesIns_Inst_Sbox_1_L2), .B0_f (new_AGEMA_signal_11852), .B1_t (new_AGEMA_signal_11853), .B1_f (new_AGEMA_signal_11854), .Z0_t (SubBytesIns_Inst_Sbox_1_L23), .Z0_f (new_AGEMA_signal_12455), .Z1_t (new_AGEMA_signal_12456), .Z1_f (new_AGEMA_signal_12457) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L15), .A0_f (new_AGEMA_signal_11867), .A1_t (new_AGEMA_signal_11868), .A1_f (new_AGEMA_signal_11869), .B0_t (SubBytesIns_Inst_Sbox_1_L9), .B0_f (new_AGEMA_signal_12440), .B1_t (new_AGEMA_signal_12441), .B1_f (new_AGEMA_signal_12442), .Z0_t (SubBytesIns_Inst_Sbox_1_L24), .Z0_f (new_AGEMA_signal_13013), .Z1_t (new_AGEMA_signal_13014), .Z1_f (new_AGEMA_signal_13015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L6), .A0_f (new_AGEMA_signal_12434), .A1_t (new_AGEMA_signal_12435), .A1_f (new_AGEMA_signal_12436), .B0_t (SubBytesIns_Inst_Sbox_1_L10), .B0_f (new_AGEMA_signal_12443), .B1_t (new_AGEMA_signal_12444), .B1_f (new_AGEMA_signal_12445), .Z0_t (SubBytesIns_Inst_Sbox_1_L25), .Z0_f (new_AGEMA_signal_13016), .Z1_t (new_AGEMA_signal_13017), .Z1_f (new_AGEMA_signal_13018) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L7), .A0_f (new_AGEMA_signal_12437), .A1_t (new_AGEMA_signal_12438), .A1_f (new_AGEMA_signal_12439), .B0_t (SubBytesIns_Inst_Sbox_1_L9), .B0_f (new_AGEMA_signal_12440), .B1_t (new_AGEMA_signal_12441), .B1_f (new_AGEMA_signal_12442), .Z0_t (SubBytesIns_Inst_Sbox_1_L26), .Z0_f (new_AGEMA_signal_13019), .Z1_t (new_AGEMA_signal_13020), .Z1_f (new_AGEMA_signal_13021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L8), .A0_f (new_AGEMA_signal_11186), .A1_t (new_AGEMA_signal_11187), .A1_f (new_AGEMA_signal_11188), .B0_t (SubBytesIns_Inst_Sbox_1_L10), .B0_f (new_AGEMA_signal_12443), .B1_t (new_AGEMA_signal_12444), .B1_f (new_AGEMA_signal_12445), .Z0_t (SubBytesIns_Inst_Sbox_1_L27), .Z0_f (new_AGEMA_signal_13022), .Z1_t (new_AGEMA_signal_13023), .Z1_f (new_AGEMA_signal_13024) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L11), .A0_f (new_AGEMA_signal_12446), .A1_t (new_AGEMA_signal_12447), .A1_f (new_AGEMA_signal_12448), .B0_t (SubBytesIns_Inst_Sbox_1_L14), .B0_f (new_AGEMA_signal_11864), .B1_t (new_AGEMA_signal_11865), .B1_f (new_AGEMA_signal_11866), .Z0_t (SubBytesIns_Inst_Sbox_1_L28), .Z0_f (new_AGEMA_signal_13025), .Z1_t (new_AGEMA_signal_13026), .Z1_f (new_AGEMA_signal_13027) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L11), .A0_f (new_AGEMA_signal_12446), .A1_t (new_AGEMA_signal_12447), .A1_f (new_AGEMA_signal_12448), .B0_t (SubBytesIns_Inst_Sbox_1_L17), .B0_f (new_AGEMA_signal_11870), .B1_t (new_AGEMA_signal_11871), .B1_f (new_AGEMA_signal_11872), .Z0_t (SubBytesIns_Inst_Sbox_1_L29), .Z0_f (new_AGEMA_signal_13028), .Z1_t (new_AGEMA_signal_13029), .Z1_f (new_AGEMA_signal_13030) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L6), .A0_f (new_AGEMA_signal_12434), .A1_t (new_AGEMA_signal_12435), .A1_f (new_AGEMA_signal_12436), .B0_t (SubBytesIns_Inst_Sbox_1_L24), .B0_f (new_AGEMA_signal_13013), .B1_t (new_AGEMA_signal_13014), .B1_f (new_AGEMA_signal_13015), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .Z0_f (new_AGEMA_signal_13661), .Z1_t (new_AGEMA_signal_13662), .Z1_f (new_AGEMA_signal_13663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L16), .A0_f (new_AGEMA_signal_13004), .A1_t (new_AGEMA_signal_13005), .A1_f (new_AGEMA_signal_13006), .B0_t (SubBytesIns_Inst_Sbox_1_L26), .B0_f (new_AGEMA_signal_13019), .B1_t (new_AGEMA_signal_13020), .B1_f (new_AGEMA_signal_13021), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .Z0_f (new_AGEMA_signal_13664), .Z1_t (new_AGEMA_signal_13665), .Z1_f (new_AGEMA_signal_13666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L19), .A0_f (new_AGEMA_signal_12449), .A1_t (new_AGEMA_signal_12450), .A1_f (new_AGEMA_signal_12451), .B0_t (SubBytesIns_Inst_Sbox_1_L28), .B0_f (new_AGEMA_signal_13025), .B1_t (new_AGEMA_signal_13026), .B1_f (new_AGEMA_signal_13027), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .Z0_f (new_AGEMA_signal_13667), .Z1_t (new_AGEMA_signal_13668), .Z1_f (new_AGEMA_signal_13669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L6), .A0_f (new_AGEMA_signal_12434), .A1_t (new_AGEMA_signal_12435), .A1_f (new_AGEMA_signal_12436), .B0_t (SubBytesIns_Inst_Sbox_1_L21), .B0_f (new_AGEMA_signal_13010), .B1_t (new_AGEMA_signal_13011), .B1_f (new_AGEMA_signal_13012), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .Z0_f (new_AGEMA_signal_13670), .Z1_t (new_AGEMA_signal_13671), .Z1_f (new_AGEMA_signal_13672) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L20), .A0_f (new_AGEMA_signal_13007), .A1_t (new_AGEMA_signal_13008), .A1_f (new_AGEMA_signal_13009), .B0_t (SubBytesIns_Inst_Sbox_1_L22), .B0_f (new_AGEMA_signal_12452), .B1_t (new_AGEMA_signal_12453), .B1_f (new_AGEMA_signal_12454), .Z0_t (MixColumnsInput[75]), .Z0_f (new_AGEMA_signal_13673), .Z1_t (new_AGEMA_signal_13674), .Z1_f (new_AGEMA_signal_13675) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L25), .A0_f (new_AGEMA_signal_13016), .A1_t (new_AGEMA_signal_13017), .A1_f (new_AGEMA_signal_13018), .B0_t (SubBytesIns_Inst_Sbox_1_L29), .B0_f (new_AGEMA_signal_13028), .B1_t (new_AGEMA_signal_13029), .B1_f (new_AGEMA_signal_13030), .Z0_t (MixColumnsInput[74]), .Z0_f (new_AGEMA_signal_13676), .Z1_t (new_AGEMA_signal_13677), .Z1_f (new_AGEMA_signal_13678) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L13), .A0_f (new_AGEMA_signal_13001), .A1_t (new_AGEMA_signal_13002), .A1_f (new_AGEMA_signal_13003), .B0_t (SubBytesIns_Inst_Sbox_1_L27), .B0_f (new_AGEMA_signal_13022), .B1_t (new_AGEMA_signal_13023), .B1_f (new_AGEMA_signal_13024), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .Z0_f (new_AGEMA_signal_13679), .Z1_t (new_AGEMA_signal_13680), .Z1_f (new_AGEMA_signal_13681) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L6), .A0_f (new_AGEMA_signal_12434), .A1_t (new_AGEMA_signal_12435), .A1_f (new_AGEMA_signal_12436), .B0_t (SubBytesIns_Inst_Sbox_1_L23), .B0_f (new_AGEMA_signal_12455), .B1_t (new_AGEMA_signal_12456), .B1_f (new_AGEMA_signal_12457), .Z0_t (MixColumnsInput[72]), .Z0_f (new_AGEMA_signal_13031), .Z1_t (new_AGEMA_signal_13032), .Z1_f (new_AGEMA_signal_13033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[23]), .A0_f (ciphertext_s0_f[23]), .A1_t (ciphertext_s1_t[23]), .A1_f (ciphertext_s1_f[23]), .B0_t (ciphertext_s0_t[20]), .B0_f (ciphertext_s0_f[20]), .B1_t (ciphertext_s1_t[20]), .B1_f (ciphertext_s1_f[20]), .Z0_t (SubBytesIns_Inst_Sbox_2_T1), .Z0_f (new_AGEMA_signal_6406), .Z1_t (new_AGEMA_signal_6407), .Z1_f (new_AGEMA_signal_6408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[23]), .A0_f (ciphertext_s0_f[23]), .A1_t (ciphertext_s1_t[23]), .A1_f (ciphertext_s1_f[23]), .B0_t (ciphertext_s0_t[18]), .B0_f (ciphertext_s0_f[18]), .B1_t (ciphertext_s1_t[18]), .B1_f (ciphertext_s1_f[18]), .Z0_t (SubBytesIns_Inst_Sbox_2_T2), .Z0_f (new_AGEMA_signal_6409), .Z1_t (new_AGEMA_signal_6410), .Z1_f (new_AGEMA_signal_6411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[23]), .A0_f (ciphertext_s0_f[23]), .A1_t (ciphertext_s1_t[23]), .A1_f (ciphertext_s1_f[23]), .B0_t (ciphertext_s0_t[17]), .B0_f (ciphertext_s0_f[17]), .B1_t (ciphertext_s1_t[17]), .B1_f (ciphertext_s1_f[17]), .Z0_t (SubBytesIns_Inst_Sbox_2_T3), .Z0_f (new_AGEMA_signal_6412), .Z1_t (new_AGEMA_signal_6413), .Z1_f (new_AGEMA_signal_6414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[20]), .A0_f (ciphertext_s0_f[20]), .A1_t (ciphertext_s1_t[20]), .A1_f (ciphertext_s1_f[20]), .B0_t (ciphertext_s0_t[18]), .B0_f (ciphertext_s0_f[18]), .B1_t (ciphertext_s1_t[18]), .B1_f (ciphertext_s1_f[18]), .Z0_t (SubBytesIns_Inst_Sbox_2_T4), .Z0_f (new_AGEMA_signal_6415), .Z1_t (new_AGEMA_signal_6416), .Z1_f (new_AGEMA_signal_6417) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[19]), .A0_f (ciphertext_s0_f[19]), .A1_t (ciphertext_s1_t[19]), .A1_f (ciphertext_s1_f[19]), .B0_t (ciphertext_s0_t[17]), .B0_f (ciphertext_s0_f[17]), .B1_t (ciphertext_s1_t[17]), .B1_f (ciphertext_s1_f[17]), .Z0_t (SubBytesIns_Inst_Sbox_2_T5), .Z0_f (new_AGEMA_signal_6418), .Z1_t (new_AGEMA_signal_6419), .Z1_f (new_AGEMA_signal_6420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T1), .A0_f (new_AGEMA_signal_6406), .A1_t (new_AGEMA_signal_6407), .A1_f (new_AGEMA_signal_6408), .B0_t (SubBytesIns_Inst_Sbox_2_T5), .B0_f (new_AGEMA_signal_6418), .B1_t (new_AGEMA_signal_6419), .B1_f (new_AGEMA_signal_6420), .Z0_t (SubBytesIns_Inst_Sbox_2_T6), .Z0_f (new_AGEMA_signal_6976), .Z1_t (new_AGEMA_signal_6977), .Z1_f (new_AGEMA_signal_6978) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[22]), .A0_f (ciphertext_s0_f[22]), .A1_t (ciphertext_s1_t[22]), .A1_f (ciphertext_s1_f[22]), .B0_t (ciphertext_s0_t[21]), .B0_f (ciphertext_s0_f[21]), .B1_t (ciphertext_s1_t[21]), .B1_f (ciphertext_s1_f[21]), .Z0_t (SubBytesIns_Inst_Sbox_2_T7), .Z0_f (new_AGEMA_signal_6421), .Z1_t (new_AGEMA_signal_6422), .Z1_f (new_AGEMA_signal_6423) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[16]), .A0_f (ciphertext_s0_f[16]), .A1_t (ciphertext_s1_t[16]), .A1_f (ciphertext_s1_f[16]), .B0_t (SubBytesIns_Inst_Sbox_2_T6), .B0_f (new_AGEMA_signal_6976), .B1_t (new_AGEMA_signal_6977), .B1_f (new_AGEMA_signal_6978), .Z0_t (SubBytesIns_Inst_Sbox_2_T8), .Z0_f (new_AGEMA_signal_7550), .Z1_t (new_AGEMA_signal_7551), .Z1_f (new_AGEMA_signal_7552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[16]), .A0_f (ciphertext_s0_f[16]), .A1_t (ciphertext_s1_t[16]), .A1_f (ciphertext_s1_f[16]), .B0_t (SubBytesIns_Inst_Sbox_2_T7), .B0_f (new_AGEMA_signal_6421), .B1_t (new_AGEMA_signal_6422), .B1_f (new_AGEMA_signal_6423), .Z0_t (SubBytesIns_Inst_Sbox_2_T9), .Z0_f (new_AGEMA_signal_6979), .Z1_t (new_AGEMA_signal_6980), .Z1_f (new_AGEMA_signal_6981) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T6), .A0_f (new_AGEMA_signal_6976), .A1_t (new_AGEMA_signal_6977), .A1_f (new_AGEMA_signal_6978), .B0_t (SubBytesIns_Inst_Sbox_2_T7), .B0_f (new_AGEMA_signal_6421), .B1_t (new_AGEMA_signal_6422), .B1_f (new_AGEMA_signal_6423), .Z0_t (SubBytesIns_Inst_Sbox_2_T10), .Z0_f (new_AGEMA_signal_7553), .Z1_t (new_AGEMA_signal_7554), .Z1_f (new_AGEMA_signal_7555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[22]), .A0_f (ciphertext_s0_f[22]), .A1_t (ciphertext_s1_t[22]), .A1_f (ciphertext_s1_f[22]), .B0_t (ciphertext_s0_t[18]), .B0_f (ciphertext_s0_f[18]), .B1_t (ciphertext_s1_t[18]), .B1_f (ciphertext_s1_f[18]), .Z0_t (SubBytesIns_Inst_Sbox_2_T11), .Z0_f (new_AGEMA_signal_6424), .Z1_t (new_AGEMA_signal_6425), .Z1_f (new_AGEMA_signal_6426) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[21]), .A0_f (ciphertext_s0_f[21]), .A1_t (ciphertext_s1_t[21]), .A1_f (ciphertext_s1_f[21]), .B0_t (ciphertext_s0_t[18]), .B0_f (ciphertext_s0_f[18]), .B1_t (ciphertext_s1_t[18]), .B1_f (ciphertext_s1_f[18]), .Z0_t (SubBytesIns_Inst_Sbox_2_T12), .Z0_f (new_AGEMA_signal_6427), .Z1_t (new_AGEMA_signal_6428), .Z1_f (new_AGEMA_signal_6429) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T3), .A0_f (new_AGEMA_signal_6412), .A1_t (new_AGEMA_signal_6413), .A1_f (new_AGEMA_signal_6414), .B0_t (SubBytesIns_Inst_Sbox_2_T4), .B0_f (new_AGEMA_signal_6415), .B1_t (new_AGEMA_signal_6416), .B1_f (new_AGEMA_signal_6417), .Z0_t (SubBytesIns_Inst_Sbox_2_T13), .Z0_f (new_AGEMA_signal_6982), .Z1_t (new_AGEMA_signal_6983), .Z1_f (new_AGEMA_signal_6984) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T6), .A0_f (new_AGEMA_signal_6976), .A1_t (new_AGEMA_signal_6977), .A1_f (new_AGEMA_signal_6978), .B0_t (SubBytesIns_Inst_Sbox_2_T11), .B0_f (new_AGEMA_signal_6424), .B1_t (new_AGEMA_signal_6425), .B1_f (new_AGEMA_signal_6426), .Z0_t (SubBytesIns_Inst_Sbox_2_T14), .Z0_f (new_AGEMA_signal_7556), .Z1_t (new_AGEMA_signal_7557), .Z1_f (new_AGEMA_signal_7558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T5), .A0_f (new_AGEMA_signal_6418), .A1_t (new_AGEMA_signal_6419), .A1_f (new_AGEMA_signal_6420), .B0_t (SubBytesIns_Inst_Sbox_2_T11), .B0_f (new_AGEMA_signal_6424), .B1_t (new_AGEMA_signal_6425), .B1_f (new_AGEMA_signal_6426), .Z0_t (SubBytesIns_Inst_Sbox_2_T15), .Z0_f (new_AGEMA_signal_6985), .Z1_t (new_AGEMA_signal_6986), .Z1_f (new_AGEMA_signal_6987) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T5), .A0_f (new_AGEMA_signal_6418), .A1_t (new_AGEMA_signal_6419), .A1_f (new_AGEMA_signal_6420), .B0_t (SubBytesIns_Inst_Sbox_2_T12), .B0_f (new_AGEMA_signal_6427), .B1_t (new_AGEMA_signal_6428), .B1_f (new_AGEMA_signal_6429), .Z0_t (SubBytesIns_Inst_Sbox_2_T16), .Z0_f (new_AGEMA_signal_6988), .Z1_t (new_AGEMA_signal_6989), .Z1_f (new_AGEMA_signal_6990) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T9), .A0_f (new_AGEMA_signal_6979), .A1_t (new_AGEMA_signal_6980), .A1_f (new_AGEMA_signal_6981), .B0_t (SubBytesIns_Inst_Sbox_2_T16), .B0_f (new_AGEMA_signal_6988), .B1_t (new_AGEMA_signal_6989), .B1_f (new_AGEMA_signal_6990), .Z0_t (SubBytesIns_Inst_Sbox_2_T17), .Z0_f (new_AGEMA_signal_7559), .Z1_t (new_AGEMA_signal_7560), .Z1_f (new_AGEMA_signal_7561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[20]), .A0_f (ciphertext_s0_f[20]), .A1_t (ciphertext_s1_t[20]), .A1_f (ciphertext_s1_f[20]), .B0_t (ciphertext_s0_t[16]), .B0_f (ciphertext_s0_f[16]), .B1_t (ciphertext_s1_t[16]), .B1_f (ciphertext_s1_f[16]), .Z0_t (SubBytesIns_Inst_Sbox_2_T18), .Z0_f (new_AGEMA_signal_6430), .Z1_t (new_AGEMA_signal_6431), .Z1_f (new_AGEMA_signal_6432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T7), .A0_f (new_AGEMA_signal_6421), .A1_t (new_AGEMA_signal_6422), .A1_f (new_AGEMA_signal_6423), .B0_t (SubBytesIns_Inst_Sbox_2_T18), .B0_f (new_AGEMA_signal_6430), .B1_t (new_AGEMA_signal_6431), .B1_f (new_AGEMA_signal_6432), .Z0_t (SubBytesIns_Inst_Sbox_2_T19), .Z0_f (new_AGEMA_signal_6991), .Z1_t (new_AGEMA_signal_6992), .Z1_f (new_AGEMA_signal_6993) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T1), .A0_f (new_AGEMA_signal_6406), .A1_t (new_AGEMA_signal_6407), .A1_f (new_AGEMA_signal_6408), .B0_t (SubBytesIns_Inst_Sbox_2_T19), .B0_f (new_AGEMA_signal_6991), .B1_t (new_AGEMA_signal_6992), .B1_f (new_AGEMA_signal_6993), .Z0_t (SubBytesIns_Inst_Sbox_2_T20), .Z0_f (new_AGEMA_signal_7562), .Z1_t (new_AGEMA_signal_7563), .Z1_f (new_AGEMA_signal_7564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[17]), .A0_f (ciphertext_s0_f[17]), .A1_t (ciphertext_s1_t[17]), .A1_f (ciphertext_s1_f[17]), .B0_t (ciphertext_s0_t[16]), .B0_f (ciphertext_s0_f[16]), .B1_t (ciphertext_s1_t[16]), .B1_f (ciphertext_s1_f[16]), .Z0_t (SubBytesIns_Inst_Sbox_2_T21), .Z0_f (new_AGEMA_signal_6433), .Z1_t (new_AGEMA_signal_6434), .Z1_f (new_AGEMA_signal_6435) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T7), .A0_f (new_AGEMA_signal_6421), .A1_t (new_AGEMA_signal_6422), .A1_f (new_AGEMA_signal_6423), .B0_t (SubBytesIns_Inst_Sbox_2_T21), .B0_f (new_AGEMA_signal_6433), .B1_t (new_AGEMA_signal_6434), .B1_f (new_AGEMA_signal_6435), .Z0_t (SubBytesIns_Inst_Sbox_2_T22), .Z0_f (new_AGEMA_signal_6994), .Z1_t (new_AGEMA_signal_6995), .Z1_f (new_AGEMA_signal_6996) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T2), .A0_f (new_AGEMA_signal_6409), .A1_t (new_AGEMA_signal_6410), .A1_f (new_AGEMA_signal_6411), .B0_t (SubBytesIns_Inst_Sbox_2_T22), .B0_f (new_AGEMA_signal_6994), .B1_t (new_AGEMA_signal_6995), .B1_f (new_AGEMA_signal_6996), .Z0_t (SubBytesIns_Inst_Sbox_2_T23), .Z0_f (new_AGEMA_signal_7565), .Z1_t (new_AGEMA_signal_7566), .Z1_f (new_AGEMA_signal_7567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T2), .A0_f (new_AGEMA_signal_6409), .A1_t (new_AGEMA_signal_6410), .A1_f (new_AGEMA_signal_6411), .B0_t (SubBytesIns_Inst_Sbox_2_T10), .B0_f (new_AGEMA_signal_7553), .B1_t (new_AGEMA_signal_7554), .B1_f (new_AGEMA_signal_7555), .Z0_t (SubBytesIns_Inst_Sbox_2_T24), .Z0_f (new_AGEMA_signal_8258), .Z1_t (new_AGEMA_signal_8259), .Z1_f (new_AGEMA_signal_8260) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T20), .A0_f (new_AGEMA_signal_7562), .A1_t (new_AGEMA_signal_7563), .A1_f (new_AGEMA_signal_7564), .B0_t (SubBytesIns_Inst_Sbox_2_T17), .B0_f (new_AGEMA_signal_7559), .B1_t (new_AGEMA_signal_7560), .B1_f (new_AGEMA_signal_7561), .Z0_t (SubBytesIns_Inst_Sbox_2_T25), .Z0_f (new_AGEMA_signal_8261), .Z1_t (new_AGEMA_signal_8262), .Z1_f (new_AGEMA_signal_8263) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T3), .A0_f (new_AGEMA_signal_6412), .A1_t (new_AGEMA_signal_6413), .A1_f (new_AGEMA_signal_6414), .B0_t (SubBytesIns_Inst_Sbox_2_T16), .B0_f (new_AGEMA_signal_6988), .B1_t (new_AGEMA_signal_6989), .B1_f (new_AGEMA_signal_6990), .Z0_t (SubBytesIns_Inst_Sbox_2_T26), .Z0_f (new_AGEMA_signal_7568), .Z1_t (new_AGEMA_signal_7569), .Z1_f (new_AGEMA_signal_7570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T1), .A0_f (new_AGEMA_signal_6406), .A1_t (new_AGEMA_signal_6407), .A1_f (new_AGEMA_signal_6408), .B0_t (SubBytesIns_Inst_Sbox_2_T12), .B0_f (new_AGEMA_signal_6427), .B1_t (new_AGEMA_signal_6428), .B1_f (new_AGEMA_signal_6429), .Z0_t (SubBytesIns_Inst_Sbox_2_T27), .Z0_f (new_AGEMA_signal_6997), .Z1_t (new_AGEMA_signal_6998), .Z1_f (new_AGEMA_signal_6999) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T13), .A0_f (new_AGEMA_signal_6982), .A1_t (new_AGEMA_signal_6983), .A1_f (new_AGEMA_signal_6984), .B0_t (SubBytesIns_Inst_Sbox_2_T6), .B0_f (new_AGEMA_signal_6976), .B1_t (new_AGEMA_signal_6977), .B1_f (new_AGEMA_signal_6978), .Z0_t (SubBytesIns_Inst_Sbox_2_M1), .Z0_f (new_AGEMA_signal_7571), .Z1_t (new_AGEMA_signal_7572), .Z1_f (new_AGEMA_signal_7573) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T23), .A0_f (new_AGEMA_signal_7565), .A1_t (new_AGEMA_signal_7566), .A1_f (new_AGEMA_signal_7567), .B0_t (SubBytesIns_Inst_Sbox_2_T8), .B0_f (new_AGEMA_signal_7550), .B1_t (new_AGEMA_signal_7551), .B1_f (new_AGEMA_signal_7552), .Z0_t (SubBytesIns_Inst_Sbox_2_M2), .Z0_f (new_AGEMA_signal_8264), .Z1_t (new_AGEMA_signal_8265), .Z1_f (new_AGEMA_signal_8266) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T14), .A0_f (new_AGEMA_signal_7556), .A1_t (new_AGEMA_signal_7557), .A1_f (new_AGEMA_signal_7558), .B0_t (SubBytesIns_Inst_Sbox_2_M1), .B0_f (new_AGEMA_signal_7571), .B1_t (new_AGEMA_signal_7572), .B1_f (new_AGEMA_signal_7573), .Z0_t (SubBytesIns_Inst_Sbox_2_M3), .Z0_f (new_AGEMA_signal_8267), .Z1_t (new_AGEMA_signal_8268), .Z1_f (new_AGEMA_signal_8269) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T19), .A0_f (new_AGEMA_signal_6991), .A1_t (new_AGEMA_signal_6992), .A1_f (new_AGEMA_signal_6993), .B0_t (ciphertext_s0_t[16]), .B0_f (ciphertext_s0_f[16]), .B1_t (ciphertext_s1_t[16]), .B1_f (ciphertext_s1_f[16]), .Z0_t (SubBytesIns_Inst_Sbox_2_M4), .Z0_f (new_AGEMA_signal_7574), .Z1_t (new_AGEMA_signal_7575), .Z1_f (new_AGEMA_signal_7576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M4), .A0_f (new_AGEMA_signal_7574), .A1_t (new_AGEMA_signal_7575), .A1_f (new_AGEMA_signal_7576), .B0_t (SubBytesIns_Inst_Sbox_2_M1), .B0_f (new_AGEMA_signal_7571), .B1_t (new_AGEMA_signal_7572), .B1_f (new_AGEMA_signal_7573), .Z0_t (SubBytesIns_Inst_Sbox_2_M5), .Z0_f (new_AGEMA_signal_8270), .Z1_t (new_AGEMA_signal_8271), .Z1_f (new_AGEMA_signal_8272) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T3), .A0_f (new_AGEMA_signal_6412), .A1_t (new_AGEMA_signal_6413), .A1_f (new_AGEMA_signal_6414), .B0_t (SubBytesIns_Inst_Sbox_2_T16), .B0_f (new_AGEMA_signal_6988), .B1_t (new_AGEMA_signal_6989), .B1_f (new_AGEMA_signal_6990), .Z0_t (SubBytesIns_Inst_Sbox_2_M6), .Z0_f (new_AGEMA_signal_7577), .Z1_t (new_AGEMA_signal_7578), .Z1_f (new_AGEMA_signal_7579) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T22), .A0_f (new_AGEMA_signal_6994), .A1_t (new_AGEMA_signal_6995), .A1_f (new_AGEMA_signal_6996), .B0_t (SubBytesIns_Inst_Sbox_2_T9), .B0_f (new_AGEMA_signal_6979), .B1_t (new_AGEMA_signal_6980), .B1_f (new_AGEMA_signal_6981), .Z0_t (SubBytesIns_Inst_Sbox_2_M7), .Z0_f (new_AGEMA_signal_7580), .Z1_t (new_AGEMA_signal_7581), .Z1_f (new_AGEMA_signal_7582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T26), .A0_f (new_AGEMA_signal_7568), .A1_t (new_AGEMA_signal_7569), .A1_f (new_AGEMA_signal_7570), .B0_t (SubBytesIns_Inst_Sbox_2_M6), .B0_f (new_AGEMA_signal_7577), .B1_t (new_AGEMA_signal_7578), .B1_f (new_AGEMA_signal_7579), .Z0_t (SubBytesIns_Inst_Sbox_2_M8), .Z0_f (new_AGEMA_signal_8273), .Z1_t (new_AGEMA_signal_8274), .Z1_f (new_AGEMA_signal_8275) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T20), .A0_f (new_AGEMA_signal_7562), .A1_t (new_AGEMA_signal_7563), .A1_f (new_AGEMA_signal_7564), .B0_t (SubBytesIns_Inst_Sbox_2_T17), .B0_f (new_AGEMA_signal_7559), .B1_t (new_AGEMA_signal_7560), .B1_f (new_AGEMA_signal_7561), .Z0_t (SubBytesIns_Inst_Sbox_2_M9), .Z0_f (new_AGEMA_signal_8276), .Z1_t (new_AGEMA_signal_8277), .Z1_f (new_AGEMA_signal_8278) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M9), .A0_f (new_AGEMA_signal_8276), .A1_t (new_AGEMA_signal_8277), .A1_f (new_AGEMA_signal_8278), .B0_t (SubBytesIns_Inst_Sbox_2_M6), .B0_f (new_AGEMA_signal_7577), .B1_t (new_AGEMA_signal_7578), .B1_f (new_AGEMA_signal_7579), .Z0_t (SubBytesIns_Inst_Sbox_2_M10), .Z0_f (new_AGEMA_signal_8726), .Z1_t (new_AGEMA_signal_8727), .Z1_f (new_AGEMA_signal_8728) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T1), .A0_f (new_AGEMA_signal_6406), .A1_t (new_AGEMA_signal_6407), .A1_f (new_AGEMA_signal_6408), .B0_t (SubBytesIns_Inst_Sbox_2_T15), .B0_f (new_AGEMA_signal_6985), .B1_t (new_AGEMA_signal_6986), .B1_f (new_AGEMA_signal_6987), .Z0_t (SubBytesIns_Inst_Sbox_2_M11), .Z0_f (new_AGEMA_signal_7583), .Z1_t (new_AGEMA_signal_7584), .Z1_f (new_AGEMA_signal_7585) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T4), .A0_f (new_AGEMA_signal_6415), .A1_t (new_AGEMA_signal_6416), .A1_f (new_AGEMA_signal_6417), .B0_t (SubBytesIns_Inst_Sbox_2_T27), .B0_f (new_AGEMA_signal_6997), .B1_t (new_AGEMA_signal_6998), .B1_f (new_AGEMA_signal_6999), .Z0_t (SubBytesIns_Inst_Sbox_2_M12), .Z0_f (new_AGEMA_signal_7586), .Z1_t (new_AGEMA_signal_7587), .Z1_f (new_AGEMA_signal_7588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M12), .A0_f (new_AGEMA_signal_7586), .A1_t (new_AGEMA_signal_7587), .A1_f (new_AGEMA_signal_7588), .B0_t (SubBytesIns_Inst_Sbox_2_M11), .B0_f (new_AGEMA_signal_7583), .B1_t (new_AGEMA_signal_7584), .B1_f (new_AGEMA_signal_7585), .Z0_t (SubBytesIns_Inst_Sbox_2_M13), .Z0_f (new_AGEMA_signal_8279), .Z1_t (new_AGEMA_signal_8280), .Z1_f (new_AGEMA_signal_8281) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T2), .A0_f (new_AGEMA_signal_6409), .A1_t (new_AGEMA_signal_6410), .A1_f (new_AGEMA_signal_6411), .B0_t (SubBytesIns_Inst_Sbox_2_T10), .B0_f (new_AGEMA_signal_7553), .B1_t (new_AGEMA_signal_7554), .B1_f (new_AGEMA_signal_7555), .Z0_t (SubBytesIns_Inst_Sbox_2_M14), .Z0_f (new_AGEMA_signal_8282), .Z1_t (new_AGEMA_signal_8283), .Z1_f (new_AGEMA_signal_8284) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M14), .A0_f (new_AGEMA_signal_8282), .A1_t (new_AGEMA_signal_8283), .A1_f (new_AGEMA_signal_8284), .B0_t (SubBytesIns_Inst_Sbox_2_M11), .B0_f (new_AGEMA_signal_7583), .B1_t (new_AGEMA_signal_7584), .B1_f (new_AGEMA_signal_7585), .Z0_t (SubBytesIns_Inst_Sbox_2_M15), .Z0_f (new_AGEMA_signal_8729), .Z1_t (new_AGEMA_signal_8730), .Z1_f (new_AGEMA_signal_8731) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M3), .A0_f (new_AGEMA_signal_8267), .A1_t (new_AGEMA_signal_8268), .A1_f (new_AGEMA_signal_8269), .B0_t (SubBytesIns_Inst_Sbox_2_M2), .B0_f (new_AGEMA_signal_8264), .B1_t (new_AGEMA_signal_8265), .B1_f (new_AGEMA_signal_8266), .Z0_t (SubBytesIns_Inst_Sbox_2_M16), .Z0_f (new_AGEMA_signal_8732), .Z1_t (new_AGEMA_signal_8733), .Z1_f (new_AGEMA_signal_8734) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M5), .A0_f (new_AGEMA_signal_8270), .A1_t (new_AGEMA_signal_8271), .A1_f (new_AGEMA_signal_8272), .B0_t (SubBytesIns_Inst_Sbox_2_T24), .B0_f (new_AGEMA_signal_8258), .B1_t (new_AGEMA_signal_8259), .B1_f (new_AGEMA_signal_8260), .Z0_t (SubBytesIns_Inst_Sbox_2_M17), .Z0_f (new_AGEMA_signal_8735), .Z1_t (new_AGEMA_signal_8736), .Z1_f (new_AGEMA_signal_8737) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M8), .A0_f (new_AGEMA_signal_8273), .A1_t (new_AGEMA_signal_8274), .A1_f (new_AGEMA_signal_8275), .B0_t (SubBytesIns_Inst_Sbox_2_M7), .B0_f (new_AGEMA_signal_7580), .B1_t (new_AGEMA_signal_7581), .B1_f (new_AGEMA_signal_7582), .Z0_t (SubBytesIns_Inst_Sbox_2_M18), .Z0_f (new_AGEMA_signal_8738), .Z1_t (new_AGEMA_signal_8739), .Z1_f (new_AGEMA_signal_8740) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M10), .A0_f (new_AGEMA_signal_8726), .A1_t (new_AGEMA_signal_8727), .A1_f (new_AGEMA_signal_8728), .B0_t (SubBytesIns_Inst_Sbox_2_M15), .B0_f (new_AGEMA_signal_8729), .B1_t (new_AGEMA_signal_8730), .B1_f (new_AGEMA_signal_8731), .Z0_t (SubBytesIns_Inst_Sbox_2_M19), .Z0_f (new_AGEMA_signal_9008), .Z1_t (new_AGEMA_signal_9009), .Z1_f (new_AGEMA_signal_9010) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M16), .A0_f (new_AGEMA_signal_8732), .A1_t (new_AGEMA_signal_8733), .A1_f (new_AGEMA_signal_8734), .B0_t (SubBytesIns_Inst_Sbox_2_M13), .B0_f (new_AGEMA_signal_8279), .B1_t (new_AGEMA_signal_8280), .B1_f (new_AGEMA_signal_8281), .Z0_t (SubBytesIns_Inst_Sbox_2_M20), .Z0_f (new_AGEMA_signal_9011), .Z1_t (new_AGEMA_signal_9012), .Z1_f (new_AGEMA_signal_9013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M17), .A0_f (new_AGEMA_signal_8735), .A1_t (new_AGEMA_signal_8736), .A1_f (new_AGEMA_signal_8737), .B0_t (SubBytesIns_Inst_Sbox_2_M15), .B0_f (new_AGEMA_signal_8729), .B1_t (new_AGEMA_signal_8730), .B1_f (new_AGEMA_signal_8731), .Z0_t (SubBytesIns_Inst_Sbox_2_M21), .Z0_f (new_AGEMA_signal_9014), .Z1_t (new_AGEMA_signal_9015), .Z1_f (new_AGEMA_signal_9016) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M18), .A0_f (new_AGEMA_signal_8738), .A1_t (new_AGEMA_signal_8739), .A1_f (new_AGEMA_signal_8740), .B0_t (SubBytesIns_Inst_Sbox_2_M13), .B0_f (new_AGEMA_signal_8279), .B1_t (new_AGEMA_signal_8280), .B1_f (new_AGEMA_signal_8281), .Z0_t (SubBytesIns_Inst_Sbox_2_M22), .Z0_f (new_AGEMA_signal_9017), .Z1_t (new_AGEMA_signal_9018), .Z1_f (new_AGEMA_signal_9019) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M19), .A0_f (new_AGEMA_signal_9008), .A1_t (new_AGEMA_signal_9009), .A1_f (new_AGEMA_signal_9010), .B0_t (SubBytesIns_Inst_Sbox_2_T25), .B0_f (new_AGEMA_signal_8261), .B1_t (new_AGEMA_signal_8262), .B1_f (new_AGEMA_signal_8263), .Z0_t (SubBytesIns_Inst_Sbox_2_M23), .Z0_f (new_AGEMA_signal_9248), .Z1_t (new_AGEMA_signal_9249), .Z1_f (new_AGEMA_signal_9250) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M22), .A0_f (new_AGEMA_signal_9017), .A1_t (new_AGEMA_signal_9018), .A1_f (new_AGEMA_signal_9019), .B0_t (SubBytesIns_Inst_Sbox_2_M23), .B0_f (new_AGEMA_signal_9248), .B1_t (new_AGEMA_signal_9249), .B1_f (new_AGEMA_signal_9250), .Z0_t (SubBytesIns_Inst_Sbox_2_M24), .Z0_f (new_AGEMA_signal_9506), .Z1_t (new_AGEMA_signal_9507), .Z1_f (new_AGEMA_signal_9508) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M22), .A0_f (new_AGEMA_signal_9017), .A1_t (new_AGEMA_signal_9018), .A1_f (new_AGEMA_signal_9019), .B0_t (SubBytesIns_Inst_Sbox_2_M20), .B0_f (new_AGEMA_signal_9011), .B1_t (new_AGEMA_signal_9012), .B1_f (new_AGEMA_signal_9013), .Z0_t (SubBytesIns_Inst_Sbox_2_M25), .Z0_f (new_AGEMA_signal_9251), .Z1_t (new_AGEMA_signal_9252), .Z1_f (new_AGEMA_signal_9253) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M21), .A0_f (new_AGEMA_signal_9014), .A1_t (new_AGEMA_signal_9015), .A1_f (new_AGEMA_signal_9016), .B0_t (SubBytesIns_Inst_Sbox_2_M25), .B0_f (new_AGEMA_signal_9251), .B1_t (new_AGEMA_signal_9252), .B1_f (new_AGEMA_signal_9253), .Z0_t (SubBytesIns_Inst_Sbox_2_M26), .Z0_f (new_AGEMA_signal_9509), .Z1_t (new_AGEMA_signal_9510), .Z1_f (new_AGEMA_signal_9511) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M20), .A0_f (new_AGEMA_signal_9011), .A1_t (new_AGEMA_signal_9012), .A1_f (new_AGEMA_signal_9013), .B0_t (SubBytesIns_Inst_Sbox_2_M21), .B0_f (new_AGEMA_signal_9014), .B1_t (new_AGEMA_signal_9015), .B1_f (new_AGEMA_signal_9016), .Z0_t (SubBytesIns_Inst_Sbox_2_M27), .Z0_f (new_AGEMA_signal_9254), .Z1_t (new_AGEMA_signal_9255), .Z1_f (new_AGEMA_signal_9256) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M23), .A0_f (new_AGEMA_signal_9248), .A1_t (new_AGEMA_signal_9249), .A1_f (new_AGEMA_signal_9250), .B0_t (SubBytesIns_Inst_Sbox_2_M25), .B0_f (new_AGEMA_signal_9251), .B1_t (new_AGEMA_signal_9252), .B1_f (new_AGEMA_signal_9253), .Z0_t (SubBytesIns_Inst_Sbox_2_M28), .Z0_f (new_AGEMA_signal_9512), .Z1_t (new_AGEMA_signal_9513), .Z1_f (new_AGEMA_signal_9514) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M28), .A0_f (new_AGEMA_signal_9512), .A1_t (new_AGEMA_signal_9513), .A1_f (new_AGEMA_signal_9514), .B0_t (SubBytesIns_Inst_Sbox_2_M27), .B0_f (new_AGEMA_signal_9254), .B1_t (new_AGEMA_signal_9255), .B1_f (new_AGEMA_signal_9256), .Z0_t (SubBytesIns_Inst_Sbox_2_M29), .Z0_f (new_AGEMA_signal_9806), .Z1_t (new_AGEMA_signal_9807), .Z1_f (new_AGEMA_signal_9808) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M26), .A0_f (new_AGEMA_signal_9509), .A1_t (new_AGEMA_signal_9510), .A1_f (new_AGEMA_signal_9511), .B0_t (SubBytesIns_Inst_Sbox_2_M24), .B0_f (new_AGEMA_signal_9506), .B1_t (new_AGEMA_signal_9507), .B1_f (new_AGEMA_signal_9508), .Z0_t (SubBytesIns_Inst_Sbox_2_M30), .Z0_f (new_AGEMA_signal_9809), .Z1_t (new_AGEMA_signal_9810), .Z1_f (new_AGEMA_signal_9811) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M20), .A0_f (new_AGEMA_signal_9011), .A1_t (new_AGEMA_signal_9012), .A1_f (new_AGEMA_signal_9013), .B0_t (SubBytesIns_Inst_Sbox_2_M23), .B0_f (new_AGEMA_signal_9248), .B1_t (new_AGEMA_signal_9249), .B1_f (new_AGEMA_signal_9250), .Z0_t (SubBytesIns_Inst_Sbox_2_M31), .Z0_f (new_AGEMA_signal_9515), .Z1_t (new_AGEMA_signal_9516), .Z1_f (new_AGEMA_signal_9517) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M27), .A0_f (new_AGEMA_signal_9254), .A1_t (new_AGEMA_signal_9255), .A1_f (new_AGEMA_signal_9256), .B0_t (SubBytesIns_Inst_Sbox_2_M31), .B0_f (new_AGEMA_signal_9515), .B1_t (new_AGEMA_signal_9516), .B1_f (new_AGEMA_signal_9517), .Z0_t (SubBytesIns_Inst_Sbox_2_M32), .Z0_f (new_AGEMA_signal_9812), .Z1_t (new_AGEMA_signal_9813), .Z1_f (new_AGEMA_signal_9814) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M27), .A0_f (new_AGEMA_signal_9254), .A1_t (new_AGEMA_signal_9255), .A1_f (new_AGEMA_signal_9256), .B0_t (SubBytesIns_Inst_Sbox_2_M25), .B0_f (new_AGEMA_signal_9251), .B1_t (new_AGEMA_signal_9252), .B1_f (new_AGEMA_signal_9253), .Z0_t (SubBytesIns_Inst_Sbox_2_M33), .Z0_f (new_AGEMA_signal_9518), .Z1_t (new_AGEMA_signal_9519), .Z1_f (new_AGEMA_signal_9520) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M21), .A0_f (new_AGEMA_signal_9014), .A1_t (new_AGEMA_signal_9015), .A1_f (new_AGEMA_signal_9016), .B0_t (SubBytesIns_Inst_Sbox_2_M22), .B0_f (new_AGEMA_signal_9017), .B1_t (new_AGEMA_signal_9018), .B1_f (new_AGEMA_signal_9019), .Z0_t (SubBytesIns_Inst_Sbox_2_M34), .Z0_f (new_AGEMA_signal_9257), .Z1_t (new_AGEMA_signal_9258), .Z1_f (new_AGEMA_signal_9259) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M24), .A0_f (new_AGEMA_signal_9506), .A1_t (new_AGEMA_signal_9507), .A1_f (new_AGEMA_signal_9508), .B0_t (SubBytesIns_Inst_Sbox_2_M34), .B0_f (new_AGEMA_signal_9257), .B1_t (new_AGEMA_signal_9258), .B1_f (new_AGEMA_signal_9259), .Z0_t (SubBytesIns_Inst_Sbox_2_M35), .Z0_f (new_AGEMA_signal_9815), .Z1_t (new_AGEMA_signal_9816), .Z1_f (new_AGEMA_signal_9817) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M24), .A0_f (new_AGEMA_signal_9506), .A1_t (new_AGEMA_signal_9507), .A1_f (new_AGEMA_signal_9508), .B0_t (SubBytesIns_Inst_Sbox_2_M25), .B0_f (new_AGEMA_signal_9251), .B1_t (new_AGEMA_signal_9252), .B1_f (new_AGEMA_signal_9253), .Z0_t (SubBytesIns_Inst_Sbox_2_M36), .Z0_f (new_AGEMA_signal_9818), .Z1_t (new_AGEMA_signal_9819), .Z1_f (new_AGEMA_signal_9820) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M21), .A0_f (new_AGEMA_signal_9014), .A1_t (new_AGEMA_signal_9015), .A1_f (new_AGEMA_signal_9016), .B0_t (SubBytesIns_Inst_Sbox_2_M29), .B0_f (new_AGEMA_signal_9806), .B1_t (new_AGEMA_signal_9807), .B1_f (new_AGEMA_signal_9808), .Z0_t (SubBytesIns_Inst_Sbox_2_M37), .Z0_f (new_AGEMA_signal_10088), .Z1_t (new_AGEMA_signal_10089), .Z1_f (new_AGEMA_signal_10090) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M32), .A0_f (new_AGEMA_signal_9812), .A1_t (new_AGEMA_signal_9813), .A1_f (new_AGEMA_signal_9814), .B0_t (SubBytesIns_Inst_Sbox_2_M33), .B0_f (new_AGEMA_signal_9518), .B1_t (new_AGEMA_signal_9519), .B1_f (new_AGEMA_signal_9520), .Z0_t (SubBytesIns_Inst_Sbox_2_M38), .Z0_f (new_AGEMA_signal_10091), .Z1_t (new_AGEMA_signal_10092), .Z1_f (new_AGEMA_signal_10093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M23), .A0_f (new_AGEMA_signal_9248), .A1_t (new_AGEMA_signal_9249), .A1_f (new_AGEMA_signal_9250), .B0_t (SubBytesIns_Inst_Sbox_2_M30), .B0_f (new_AGEMA_signal_9809), .B1_t (new_AGEMA_signal_9810), .B1_f (new_AGEMA_signal_9811), .Z0_t (SubBytesIns_Inst_Sbox_2_M39), .Z0_f (new_AGEMA_signal_10094), .Z1_t (new_AGEMA_signal_10095), .Z1_f (new_AGEMA_signal_10096) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M35), .A0_f (new_AGEMA_signal_9815), .A1_t (new_AGEMA_signal_9816), .A1_f (new_AGEMA_signal_9817), .B0_t (SubBytesIns_Inst_Sbox_2_M36), .B0_f (new_AGEMA_signal_9818), .B1_t (new_AGEMA_signal_9819), .B1_f (new_AGEMA_signal_9820), .Z0_t (SubBytesIns_Inst_Sbox_2_M40), .Z0_f (new_AGEMA_signal_10097), .Z1_t (new_AGEMA_signal_10098), .Z1_f (new_AGEMA_signal_10099) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M38), .A0_f (new_AGEMA_signal_10091), .A1_t (new_AGEMA_signal_10092), .A1_f (new_AGEMA_signal_10093), .B0_t (SubBytesIns_Inst_Sbox_2_M40), .B0_f (new_AGEMA_signal_10097), .B1_t (new_AGEMA_signal_10098), .B1_f (new_AGEMA_signal_10099), .Z0_t (SubBytesIns_Inst_Sbox_2_M41), .Z0_f (new_AGEMA_signal_10472), .Z1_t (new_AGEMA_signal_10473), .Z1_f (new_AGEMA_signal_10474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M37), .A0_f (new_AGEMA_signal_10088), .A1_t (new_AGEMA_signal_10089), .A1_f (new_AGEMA_signal_10090), .B0_t (SubBytesIns_Inst_Sbox_2_M39), .B0_f (new_AGEMA_signal_10094), .B1_t (new_AGEMA_signal_10095), .B1_f (new_AGEMA_signal_10096), .Z0_t (SubBytesIns_Inst_Sbox_2_M42), .Z0_f (new_AGEMA_signal_10475), .Z1_t (new_AGEMA_signal_10476), .Z1_f (new_AGEMA_signal_10477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M37), .A0_f (new_AGEMA_signal_10088), .A1_t (new_AGEMA_signal_10089), .A1_f (new_AGEMA_signal_10090), .B0_t (SubBytesIns_Inst_Sbox_2_M38), .B0_f (new_AGEMA_signal_10091), .B1_t (new_AGEMA_signal_10092), .B1_f (new_AGEMA_signal_10093), .Z0_t (SubBytesIns_Inst_Sbox_2_M43), .Z0_f (new_AGEMA_signal_10478), .Z1_t (new_AGEMA_signal_10479), .Z1_f (new_AGEMA_signal_10480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M39), .A0_f (new_AGEMA_signal_10094), .A1_t (new_AGEMA_signal_10095), .A1_f (new_AGEMA_signal_10096), .B0_t (SubBytesIns_Inst_Sbox_2_M40), .B0_f (new_AGEMA_signal_10097), .B1_t (new_AGEMA_signal_10098), .B1_f (new_AGEMA_signal_10099), .Z0_t (SubBytesIns_Inst_Sbox_2_M44), .Z0_f (new_AGEMA_signal_10481), .Z1_t (new_AGEMA_signal_10482), .Z1_f (new_AGEMA_signal_10483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M42), .A0_f (new_AGEMA_signal_10475), .A1_t (new_AGEMA_signal_10476), .A1_f (new_AGEMA_signal_10477), .B0_t (SubBytesIns_Inst_Sbox_2_M41), .B0_f (new_AGEMA_signal_10472), .B1_t (new_AGEMA_signal_10473), .B1_f (new_AGEMA_signal_10474), .Z0_t (SubBytesIns_Inst_Sbox_2_M45), .Z0_f (new_AGEMA_signal_11192), .Z1_t (new_AGEMA_signal_11193), .Z1_f (new_AGEMA_signal_11194) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M44), .A0_f (new_AGEMA_signal_10481), .A1_t (new_AGEMA_signal_10482), .A1_f (new_AGEMA_signal_10483), .B0_t (SubBytesIns_Inst_Sbox_2_T6), .B0_f (new_AGEMA_signal_6976), .B1_t (new_AGEMA_signal_6977), .B1_f (new_AGEMA_signal_6978), .Z0_t (SubBytesIns_Inst_Sbox_2_M46), .Z0_f (new_AGEMA_signal_11195), .Z1_t (new_AGEMA_signal_11196), .Z1_f (new_AGEMA_signal_11197) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M40), .A0_f (new_AGEMA_signal_10097), .A1_t (new_AGEMA_signal_10098), .A1_f (new_AGEMA_signal_10099), .B0_t (SubBytesIns_Inst_Sbox_2_T8), .B0_f (new_AGEMA_signal_7550), .B1_t (new_AGEMA_signal_7551), .B1_f (new_AGEMA_signal_7552), .Z0_t (SubBytesIns_Inst_Sbox_2_M47), .Z0_f (new_AGEMA_signal_10484), .Z1_t (new_AGEMA_signal_10485), .Z1_f (new_AGEMA_signal_10486) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M39), .A0_f (new_AGEMA_signal_10094), .A1_t (new_AGEMA_signal_10095), .A1_f (new_AGEMA_signal_10096), .B0_t (ciphertext_s0_t[16]), .B0_f (ciphertext_s0_f[16]), .B1_t (ciphertext_s1_t[16]), .B1_f (ciphertext_s1_f[16]), .Z0_t (SubBytesIns_Inst_Sbox_2_M48), .Z0_f (new_AGEMA_signal_10487), .Z1_t (new_AGEMA_signal_10488), .Z1_f (new_AGEMA_signal_10489) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M43), .A0_f (new_AGEMA_signal_10478), .A1_t (new_AGEMA_signal_10479), .A1_f (new_AGEMA_signal_10480), .B0_t (SubBytesIns_Inst_Sbox_2_T16), .B0_f (new_AGEMA_signal_6988), .B1_t (new_AGEMA_signal_6989), .B1_f (new_AGEMA_signal_6990), .Z0_t (SubBytesIns_Inst_Sbox_2_M49), .Z0_f (new_AGEMA_signal_11198), .Z1_t (new_AGEMA_signal_11199), .Z1_f (new_AGEMA_signal_11200) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M38), .A0_f (new_AGEMA_signal_10091), .A1_t (new_AGEMA_signal_10092), .A1_f (new_AGEMA_signal_10093), .B0_t (SubBytesIns_Inst_Sbox_2_T9), .B0_f (new_AGEMA_signal_6979), .B1_t (new_AGEMA_signal_6980), .B1_f (new_AGEMA_signal_6981), .Z0_t (SubBytesIns_Inst_Sbox_2_M50), .Z0_f (new_AGEMA_signal_10490), .Z1_t (new_AGEMA_signal_10491), .Z1_f (new_AGEMA_signal_10492) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M37), .A0_f (new_AGEMA_signal_10088), .A1_t (new_AGEMA_signal_10089), .A1_f (new_AGEMA_signal_10090), .B0_t (SubBytesIns_Inst_Sbox_2_T17), .B0_f (new_AGEMA_signal_7559), .B1_t (new_AGEMA_signal_7560), .B1_f (new_AGEMA_signal_7561), .Z0_t (SubBytesIns_Inst_Sbox_2_M51), .Z0_f (new_AGEMA_signal_10493), .Z1_t (new_AGEMA_signal_10494), .Z1_f (new_AGEMA_signal_10495) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M42), .A0_f (new_AGEMA_signal_10475), .A1_t (new_AGEMA_signal_10476), .A1_f (new_AGEMA_signal_10477), .B0_t (SubBytesIns_Inst_Sbox_2_T15), .B0_f (new_AGEMA_signal_6985), .B1_t (new_AGEMA_signal_6986), .B1_f (new_AGEMA_signal_6987), .Z0_t (SubBytesIns_Inst_Sbox_2_M52), .Z0_f (new_AGEMA_signal_11201), .Z1_t (new_AGEMA_signal_11202), .Z1_f (new_AGEMA_signal_11203) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M45), .A0_f (new_AGEMA_signal_11192), .A1_t (new_AGEMA_signal_11193), .A1_f (new_AGEMA_signal_11194), .B0_t (SubBytesIns_Inst_Sbox_2_T27), .B0_f (new_AGEMA_signal_6997), .B1_t (new_AGEMA_signal_6998), .B1_f (new_AGEMA_signal_6999), .Z0_t (SubBytesIns_Inst_Sbox_2_M53), .Z0_f (new_AGEMA_signal_11876), .Z1_t (new_AGEMA_signal_11877), .Z1_f (new_AGEMA_signal_11878) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M41), .A0_f (new_AGEMA_signal_10472), .A1_t (new_AGEMA_signal_10473), .A1_f (new_AGEMA_signal_10474), .B0_t (SubBytesIns_Inst_Sbox_2_T10), .B0_f (new_AGEMA_signal_7553), .B1_t (new_AGEMA_signal_7554), .B1_f (new_AGEMA_signal_7555), .Z0_t (SubBytesIns_Inst_Sbox_2_M54), .Z0_f (new_AGEMA_signal_11204), .Z1_t (new_AGEMA_signal_11205), .Z1_f (new_AGEMA_signal_11206) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M44), .A0_f (new_AGEMA_signal_10481), .A1_t (new_AGEMA_signal_10482), .A1_f (new_AGEMA_signal_10483), .B0_t (SubBytesIns_Inst_Sbox_2_T13), .B0_f (new_AGEMA_signal_6982), .B1_t (new_AGEMA_signal_6983), .B1_f (new_AGEMA_signal_6984), .Z0_t (SubBytesIns_Inst_Sbox_2_M55), .Z0_f (new_AGEMA_signal_11207), .Z1_t (new_AGEMA_signal_11208), .Z1_f (new_AGEMA_signal_11209) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M40), .A0_f (new_AGEMA_signal_10097), .A1_t (new_AGEMA_signal_10098), .A1_f (new_AGEMA_signal_10099), .B0_t (SubBytesIns_Inst_Sbox_2_T23), .B0_f (new_AGEMA_signal_7565), .B1_t (new_AGEMA_signal_7566), .B1_f (new_AGEMA_signal_7567), .Z0_t (SubBytesIns_Inst_Sbox_2_M56), .Z0_f (new_AGEMA_signal_10496), .Z1_t (new_AGEMA_signal_10497), .Z1_f (new_AGEMA_signal_10498) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M39), .A0_f (new_AGEMA_signal_10094), .A1_t (new_AGEMA_signal_10095), .A1_f (new_AGEMA_signal_10096), .B0_t (SubBytesIns_Inst_Sbox_2_T19), .B0_f (new_AGEMA_signal_6991), .B1_t (new_AGEMA_signal_6992), .B1_f (new_AGEMA_signal_6993), .Z0_t (SubBytesIns_Inst_Sbox_2_M57), .Z0_f (new_AGEMA_signal_10499), .Z1_t (new_AGEMA_signal_10500), .Z1_f (new_AGEMA_signal_10501) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M43), .A0_f (new_AGEMA_signal_10478), .A1_t (new_AGEMA_signal_10479), .A1_f (new_AGEMA_signal_10480), .B0_t (SubBytesIns_Inst_Sbox_2_T3), .B0_f (new_AGEMA_signal_6412), .B1_t (new_AGEMA_signal_6413), .B1_f (new_AGEMA_signal_6414), .Z0_t (SubBytesIns_Inst_Sbox_2_M58), .Z0_f (new_AGEMA_signal_11210), .Z1_t (new_AGEMA_signal_11211), .Z1_f (new_AGEMA_signal_11212) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M38), .A0_f (new_AGEMA_signal_10091), .A1_t (new_AGEMA_signal_10092), .A1_f (new_AGEMA_signal_10093), .B0_t (SubBytesIns_Inst_Sbox_2_T22), .B0_f (new_AGEMA_signal_6994), .B1_t (new_AGEMA_signal_6995), .B1_f (new_AGEMA_signal_6996), .Z0_t (SubBytesIns_Inst_Sbox_2_M59), .Z0_f (new_AGEMA_signal_10502), .Z1_t (new_AGEMA_signal_10503), .Z1_f (new_AGEMA_signal_10504) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M37), .A0_f (new_AGEMA_signal_10088), .A1_t (new_AGEMA_signal_10089), .A1_f (new_AGEMA_signal_10090), .B0_t (SubBytesIns_Inst_Sbox_2_T20), .B0_f (new_AGEMA_signal_7562), .B1_t (new_AGEMA_signal_7563), .B1_f (new_AGEMA_signal_7564), .Z0_t (SubBytesIns_Inst_Sbox_2_M60), .Z0_f (new_AGEMA_signal_10505), .Z1_t (new_AGEMA_signal_10506), .Z1_f (new_AGEMA_signal_10507) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M42), .A0_f (new_AGEMA_signal_10475), .A1_t (new_AGEMA_signal_10476), .A1_f (new_AGEMA_signal_10477), .B0_t (SubBytesIns_Inst_Sbox_2_T1), .B0_f (new_AGEMA_signal_6406), .B1_t (new_AGEMA_signal_6407), .B1_f (new_AGEMA_signal_6408), .Z0_t (SubBytesIns_Inst_Sbox_2_M61), .Z0_f (new_AGEMA_signal_11213), .Z1_t (new_AGEMA_signal_11214), .Z1_f (new_AGEMA_signal_11215) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M45), .A0_f (new_AGEMA_signal_11192), .A1_t (new_AGEMA_signal_11193), .A1_f (new_AGEMA_signal_11194), .B0_t (SubBytesIns_Inst_Sbox_2_T4), .B0_f (new_AGEMA_signal_6415), .B1_t (new_AGEMA_signal_6416), .B1_f (new_AGEMA_signal_6417), .Z0_t (SubBytesIns_Inst_Sbox_2_M62), .Z0_f (new_AGEMA_signal_11879), .Z1_t (new_AGEMA_signal_11880), .Z1_f (new_AGEMA_signal_11881) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M41), .A0_f (new_AGEMA_signal_10472), .A1_t (new_AGEMA_signal_10473), .A1_f (new_AGEMA_signal_10474), .B0_t (SubBytesIns_Inst_Sbox_2_T2), .B0_f (new_AGEMA_signal_6409), .B1_t (new_AGEMA_signal_6410), .B1_f (new_AGEMA_signal_6411), .Z0_t (SubBytesIns_Inst_Sbox_2_M63), .Z0_f (new_AGEMA_signal_11216), .Z1_t (new_AGEMA_signal_11217), .Z1_f (new_AGEMA_signal_11218) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M61), .A0_f (new_AGEMA_signal_11213), .A1_t (new_AGEMA_signal_11214), .A1_f (new_AGEMA_signal_11215), .B0_t (SubBytesIns_Inst_Sbox_2_M62), .B0_f (new_AGEMA_signal_11879), .B1_t (new_AGEMA_signal_11880), .B1_f (new_AGEMA_signal_11881), .Z0_t (SubBytesIns_Inst_Sbox_2_L0), .Z0_f (new_AGEMA_signal_12458), .Z1_t (new_AGEMA_signal_12459), .Z1_f (new_AGEMA_signal_12460) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M50), .A0_f (new_AGEMA_signal_10490), .A1_t (new_AGEMA_signal_10491), .A1_f (new_AGEMA_signal_10492), .B0_t (SubBytesIns_Inst_Sbox_2_M56), .B0_f (new_AGEMA_signal_10496), .B1_t (new_AGEMA_signal_10497), .B1_f (new_AGEMA_signal_10498), .Z0_t (SubBytesIns_Inst_Sbox_2_L1), .Z0_f (new_AGEMA_signal_11219), .Z1_t (new_AGEMA_signal_11220), .Z1_f (new_AGEMA_signal_11221) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M46), .A0_f (new_AGEMA_signal_11195), .A1_t (new_AGEMA_signal_11196), .A1_f (new_AGEMA_signal_11197), .B0_t (SubBytesIns_Inst_Sbox_2_M48), .B0_f (new_AGEMA_signal_10487), .B1_t (new_AGEMA_signal_10488), .B1_f (new_AGEMA_signal_10489), .Z0_t (SubBytesIns_Inst_Sbox_2_L2), .Z0_f (new_AGEMA_signal_11882), .Z1_t (new_AGEMA_signal_11883), .Z1_f (new_AGEMA_signal_11884) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M47), .A0_f (new_AGEMA_signal_10484), .A1_t (new_AGEMA_signal_10485), .A1_f (new_AGEMA_signal_10486), .B0_t (SubBytesIns_Inst_Sbox_2_M55), .B0_f (new_AGEMA_signal_11207), .B1_t (new_AGEMA_signal_11208), .B1_f (new_AGEMA_signal_11209), .Z0_t (SubBytesIns_Inst_Sbox_2_L3), .Z0_f (new_AGEMA_signal_11885), .Z1_t (new_AGEMA_signal_11886), .Z1_f (new_AGEMA_signal_11887) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M54), .A0_f (new_AGEMA_signal_11204), .A1_t (new_AGEMA_signal_11205), .A1_f (new_AGEMA_signal_11206), .B0_t (SubBytesIns_Inst_Sbox_2_M58), .B0_f (new_AGEMA_signal_11210), .B1_t (new_AGEMA_signal_11211), .B1_f (new_AGEMA_signal_11212), .Z0_t (SubBytesIns_Inst_Sbox_2_L4), .Z0_f (new_AGEMA_signal_11888), .Z1_t (new_AGEMA_signal_11889), .Z1_f (new_AGEMA_signal_11890) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M49), .A0_f (new_AGEMA_signal_11198), .A1_t (new_AGEMA_signal_11199), .A1_f (new_AGEMA_signal_11200), .B0_t (SubBytesIns_Inst_Sbox_2_M61), .B0_f (new_AGEMA_signal_11213), .B1_t (new_AGEMA_signal_11214), .B1_f (new_AGEMA_signal_11215), .Z0_t (SubBytesIns_Inst_Sbox_2_L5), .Z0_f (new_AGEMA_signal_11891), .Z1_t (new_AGEMA_signal_11892), .Z1_f (new_AGEMA_signal_11893) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M62), .A0_f (new_AGEMA_signal_11879), .A1_t (new_AGEMA_signal_11880), .A1_f (new_AGEMA_signal_11881), .B0_t (SubBytesIns_Inst_Sbox_2_L5), .B0_f (new_AGEMA_signal_11891), .B1_t (new_AGEMA_signal_11892), .B1_f (new_AGEMA_signal_11893), .Z0_t (SubBytesIns_Inst_Sbox_2_L6), .Z0_f (new_AGEMA_signal_12461), .Z1_t (new_AGEMA_signal_12462), .Z1_f (new_AGEMA_signal_12463) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M46), .A0_f (new_AGEMA_signal_11195), .A1_t (new_AGEMA_signal_11196), .A1_f (new_AGEMA_signal_11197), .B0_t (SubBytesIns_Inst_Sbox_2_L3), .B0_f (new_AGEMA_signal_11885), .B1_t (new_AGEMA_signal_11886), .B1_f (new_AGEMA_signal_11887), .Z0_t (SubBytesIns_Inst_Sbox_2_L7), .Z0_f (new_AGEMA_signal_12464), .Z1_t (new_AGEMA_signal_12465), .Z1_f (new_AGEMA_signal_12466) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M51), .A0_f (new_AGEMA_signal_10493), .A1_t (new_AGEMA_signal_10494), .A1_f (new_AGEMA_signal_10495), .B0_t (SubBytesIns_Inst_Sbox_2_M59), .B0_f (new_AGEMA_signal_10502), .B1_t (new_AGEMA_signal_10503), .B1_f (new_AGEMA_signal_10504), .Z0_t (SubBytesIns_Inst_Sbox_2_L8), .Z0_f (new_AGEMA_signal_11222), .Z1_t (new_AGEMA_signal_11223), .Z1_f (new_AGEMA_signal_11224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M52), .A0_f (new_AGEMA_signal_11201), .A1_t (new_AGEMA_signal_11202), .A1_f (new_AGEMA_signal_11203), .B0_t (SubBytesIns_Inst_Sbox_2_M53), .B0_f (new_AGEMA_signal_11876), .B1_t (new_AGEMA_signal_11877), .B1_f (new_AGEMA_signal_11878), .Z0_t (SubBytesIns_Inst_Sbox_2_L9), .Z0_f (new_AGEMA_signal_12467), .Z1_t (new_AGEMA_signal_12468), .Z1_f (new_AGEMA_signal_12469) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M53), .A0_f (new_AGEMA_signal_11876), .A1_t (new_AGEMA_signal_11877), .A1_f (new_AGEMA_signal_11878), .B0_t (SubBytesIns_Inst_Sbox_2_L4), .B0_f (new_AGEMA_signal_11888), .B1_t (new_AGEMA_signal_11889), .B1_f (new_AGEMA_signal_11890), .Z0_t (SubBytesIns_Inst_Sbox_2_L10), .Z0_f (new_AGEMA_signal_12470), .Z1_t (new_AGEMA_signal_12471), .Z1_f (new_AGEMA_signal_12472) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M60), .A0_f (new_AGEMA_signal_10505), .A1_t (new_AGEMA_signal_10506), .A1_f (new_AGEMA_signal_10507), .B0_t (SubBytesIns_Inst_Sbox_2_L2), .B0_f (new_AGEMA_signal_11882), .B1_t (new_AGEMA_signal_11883), .B1_f (new_AGEMA_signal_11884), .Z0_t (SubBytesIns_Inst_Sbox_2_L11), .Z0_f (new_AGEMA_signal_12473), .Z1_t (new_AGEMA_signal_12474), .Z1_f (new_AGEMA_signal_12475) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M48), .A0_f (new_AGEMA_signal_10487), .A1_t (new_AGEMA_signal_10488), .A1_f (new_AGEMA_signal_10489), .B0_t (SubBytesIns_Inst_Sbox_2_M51), .B0_f (new_AGEMA_signal_10493), .B1_t (new_AGEMA_signal_10494), .B1_f (new_AGEMA_signal_10495), .Z0_t (SubBytesIns_Inst_Sbox_2_L12), .Z0_f (new_AGEMA_signal_11225), .Z1_t (new_AGEMA_signal_11226), .Z1_f (new_AGEMA_signal_11227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M50), .A0_f (new_AGEMA_signal_10490), .A1_t (new_AGEMA_signal_10491), .A1_f (new_AGEMA_signal_10492), .B0_t (SubBytesIns_Inst_Sbox_2_L0), .B0_f (new_AGEMA_signal_12458), .B1_t (new_AGEMA_signal_12459), .B1_f (new_AGEMA_signal_12460), .Z0_t (SubBytesIns_Inst_Sbox_2_L13), .Z0_f (new_AGEMA_signal_13034), .Z1_t (new_AGEMA_signal_13035), .Z1_f (new_AGEMA_signal_13036) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M52), .A0_f (new_AGEMA_signal_11201), .A1_t (new_AGEMA_signal_11202), .A1_f (new_AGEMA_signal_11203), .B0_t (SubBytesIns_Inst_Sbox_2_M61), .B0_f (new_AGEMA_signal_11213), .B1_t (new_AGEMA_signal_11214), .B1_f (new_AGEMA_signal_11215), .Z0_t (SubBytesIns_Inst_Sbox_2_L14), .Z0_f (new_AGEMA_signal_11894), .Z1_t (new_AGEMA_signal_11895), .Z1_f (new_AGEMA_signal_11896) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M55), .A0_f (new_AGEMA_signal_11207), .A1_t (new_AGEMA_signal_11208), .A1_f (new_AGEMA_signal_11209), .B0_t (SubBytesIns_Inst_Sbox_2_L1), .B0_f (new_AGEMA_signal_11219), .B1_t (new_AGEMA_signal_11220), .B1_f (new_AGEMA_signal_11221), .Z0_t (SubBytesIns_Inst_Sbox_2_L15), .Z0_f (new_AGEMA_signal_11897), .Z1_t (new_AGEMA_signal_11898), .Z1_f (new_AGEMA_signal_11899) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M56), .A0_f (new_AGEMA_signal_10496), .A1_t (new_AGEMA_signal_10497), .A1_f (new_AGEMA_signal_10498), .B0_t (SubBytesIns_Inst_Sbox_2_L0), .B0_f (new_AGEMA_signal_12458), .B1_t (new_AGEMA_signal_12459), .B1_f (new_AGEMA_signal_12460), .Z0_t (SubBytesIns_Inst_Sbox_2_L16), .Z0_f (new_AGEMA_signal_13037), .Z1_t (new_AGEMA_signal_13038), .Z1_f (new_AGEMA_signal_13039) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M57), .A0_f (new_AGEMA_signal_10499), .A1_t (new_AGEMA_signal_10500), .A1_f (new_AGEMA_signal_10501), .B0_t (SubBytesIns_Inst_Sbox_2_L1), .B0_f (new_AGEMA_signal_11219), .B1_t (new_AGEMA_signal_11220), .B1_f (new_AGEMA_signal_11221), .Z0_t (SubBytesIns_Inst_Sbox_2_L17), .Z0_f (new_AGEMA_signal_11900), .Z1_t (new_AGEMA_signal_11901), .Z1_f (new_AGEMA_signal_11902) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M58), .A0_f (new_AGEMA_signal_11210), .A1_t (new_AGEMA_signal_11211), .A1_f (new_AGEMA_signal_11212), .B0_t (SubBytesIns_Inst_Sbox_2_L8), .B0_f (new_AGEMA_signal_11222), .B1_t (new_AGEMA_signal_11223), .B1_f (new_AGEMA_signal_11224), .Z0_t (SubBytesIns_Inst_Sbox_2_L18), .Z0_f (new_AGEMA_signal_11903), .Z1_t (new_AGEMA_signal_11904), .Z1_f (new_AGEMA_signal_11905) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M63), .A0_f (new_AGEMA_signal_11216), .A1_t (new_AGEMA_signal_11217), .A1_f (new_AGEMA_signal_11218), .B0_t (SubBytesIns_Inst_Sbox_2_L4), .B0_f (new_AGEMA_signal_11888), .B1_t (new_AGEMA_signal_11889), .B1_f (new_AGEMA_signal_11890), .Z0_t (SubBytesIns_Inst_Sbox_2_L19), .Z0_f (new_AGEMA_signal_12476), .Z1_t (new_AGEMA_signal_12477), .Z1_f (new_AGEMA_signal_12478) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L0), .A0_f (new_AGEMA_signal_12458), .A1_t (new_AGEMA_signal_12459), .A1_f (new_AGEMA_signal_12460), .B0_t (SubBytesIns_Inst_Sbox_2_L1), .B0_f (new_AGEMA_signal_11219), .B1_t (new_AGEMA_signal_11220), .B1_f (new_AGEMA_signal_11221), .Z0_t (SubBytesIns_Inst_Sbox_2_L20), .Z0_f (new_AGEMA_signal_13040), .Z1_t (new_AGEMA_signal_13041), .Z1_f (new_AGEMA_signal_13042) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L1), .A0_f (new_AGEMA_signal_11219), .A1_t (new_AGEMA_signal_11220), .A1_f (new_AGEMA_signal_11221), .B0_t (SubBytesIns_Inst_Sbox_2_L7), .B0_f (new_AGEMA_signal_12464), .B1_t (new_AGEMA_signal_12465), .B1_f (new_AGEMA_signal_12466), .Z0_t (SubBytesIns_Inst_Sbox_2_L21), .Z0_f (new_AGEMA_signal_13043), .Z1_t (new_AGEMA_signal_13044), .Z1_f (new_AGEMA_signal_13045) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L3), .A0_f (new_AGEMA_signal_11885), .A1_t (new_AGEMA_signal_11886), .A1_f (new_AGEMA_signal_11887), .B0_t (SubBytesIns_Inst_Sbox_2_L12), .B0_f (new_AGEMA_signal_11225), .B1_t (new_AGEMA_signal_11226), .B1_f (new_AGEMA_signal_11227), .Z0_t (SubBytesIns_Inst_Sbox_2_L22), .Z0_f (new_AGEMA_signal_12479), .Z1_t (new_AGEMA_signal_12480), .Z1_f (new_AGEMA_signal_12481) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L18), .A0_f (new_AGEMA_signal_11903), .A1_t (new_AGEMA_signal_11904), .A1_f (new_AGEMA_signal_11905), .B0_t (SubBytesIns_Inst_Sbox_2_L2), .B0_f (new_AGEMA_signal_11882), .B1_t (new_AGEMA_signal_11883), .B1_f (new_AGEMA_signal_11884), .Z0_t (SubBytesIns_Inst_Sbox_2_L23), .Z0_f (new_AGEMA_signal_12482), .Z1_t (new_AGEMA_signal_12483), .Z1_f (new_AGEMA_signal_12484) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L15), .A0_f (new_AGEMA_signal_11897), .A1_t (new_AGEMA_signal_11898), .A1_f (new_AGEMA_signal_11899), .B0_t (SubBytesIns_Inst_Sbox_2_L9), .B0_f (new_AGEMA_signal_12467), .B1_t (new_AGEMA_signal_12468), .B1_f (new_AGEMA_signal_12469), .Z0_t (SubBytesIns_Inst_Sbox_2_L24), .Z0_f (new_AGEMA_signal_13046), .Z1_t (new_AGEMA_signal_13047), .Z1_f (new_AGEMA_signal_13048) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L6), .A0_f (new_AGEMA_signal_12461), .A1_t (new_AGEMA_signal_12462), .A1_f (new_AGEMA_signal_12463), .B0_t (SubBytesIns_Inst_Sbox_2_L10), .B0_f (new_AGEMA_signal_12470), .B1_t (new_AGEMA_signal_12471), .B1_f (new_AGEMA_signal_12472), .Z0_t (SubBytesIns_Inst_Sbox_2_L25), .Z0_f (new_AGEMA_signal_13049), .Z1_t (new_AGEMA_signal_13050), .Z1_f (new_AGEMA_signal_13051) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L7), .A0_f (new_AGEMA_signal_12464), .A1_t (new_AGEMA_signal_12465), .A1_f (new_AGEMA_signal_12466), .B0_t (SubBytesIns_Inst_Sbox_2_L9), .B0_f (new_AGEMA_signal_12467), .B1_t (new_AGEMA_signal_12468), .B1_f (new_AGEMA_signal_12469), .Z0_t (SubBytesIns_Inst_Sbox_2_L26), .Z0_f (new_AGEMA_signal_13052), .Z1_t (new_AGEMA_signal_13053), .Z1_f (new_AGEMA_signal_13054) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L8), .A0_f (new_AGEMA_signal_11222), .A1_t (new_AGEMA_signal_11223), .A1_f (new_AGEMA_signal_11224), .B0_t (SubBytesIns_Inst_Sbox_2_L10), .B0_f (new_AGEMA_signal_12470), .B1_t (new_AGEMA_signal_12471), .B1_f (new_AGEMA_signal_12472), .Z0_t (SubBytesIns_Inst_Sbox_2_L27), .Z0_f (new_AGEMA_signal_13055), .Z1_t (new_AGEMA_signal_13056), .Z1_f (new_AGEMA_signal_13057) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L11), .A0_f (new_AGEMA_signal_12473), .A1_t (new_AGEMA_signal_12474), .A1_f (new_AGEMA_signal_12475), .B0_t (SubBytesIns_Inst_Sbox_2_L14), .B0_f (new_AGEMA_signal_11894), .B1_t (new_AGEMA_signal_11895), .B1_f (new_AGEMA_signal_11896), .Z0_t (SubBytesIns_Inst_Sbox_2_L28), .Z0_f (new_AGEMA_signal_13058), .Z1_t (new_AGEMA_signal_13059), .Z1_f (new_AGEMA_signal_13060) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L11), .A0_f (new_AGEMA_signal_12473), .A1_t (new_AGEMA_signal_12474), .A1_f (new_AGEMA_signal_12475), .B0_t (SubBytesIns_Inst_Sbox_2_L17), .B0_f (new_AGEMA_signal_11900), .B1_t (new_AGEMA_signal_11901), .B1_f (new_AGEMA_signal_11902), .Z0_t (SubBytesIns_Inst_Sbox_2_L29), .Z0_f (new_AGEMA_signal_13061), .Z1_t (new_AGEMA_signal_13062), .Z1_f (new_AGEMA_signal_13063) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L6), .A0_f (new_AGEMA_signal_12461), .A1_t (new_AGEMA_signal_12462), .A1_f (new_AGEMA_signal_12463), .B0_t (SubBytesIns_Inst_Sbox_2_L24), .B0_f (new_AGEMA_signal_13046), .B1_t (new_AGEMA_signal_13047), .B1_f (new_AGEMA_signal_13048), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .Z0_f (new_AGEMA_signal_13682), .Z1_t (new_AGEMA_signal_13683), .Z1_f (new_AGEMA_signal_13684) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L16), .A0_f (new_AGEMA_signal_13037), .A1_t (new_AGEMA_signal_13038), .A1_f (new_AGEMA_signal_13039), .B0_t (SubBytesIns_Inst_Sbox_2_L26), .B0_f (new_AGEMA_signal_13052), .B1_t (new_AGEMA_signal_13053), .B1_f (new_AGEMA_signal_13054), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .Z0_f (new_AGEMA_signal_13685), .Z1_t (new_AGEMA_signal_13686), .Z1_f (new_AGEMA_signal_13687) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L19), .A0_f (new_AGEMA_signal_12476), .A1_t (new_AGEMA_signal_12477), .A1_f (new_AGEMA_signal_12478), .B0_t (SubBytesIns_Inst_Sbox_2_L28), .B0_f (new_AGEMA_signal_13058), .B1_t (new_AGEMA_signal_13059), .B1_f (new_AGEMA_signal_13060), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .Z0_f (new_AGEMA_signal_13688), .Z1_t (new_AGEMA_signal_13689), .Z1_f (new_AGEMA_signal_13690) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L6), .A0_f (new_AGEMA_signal_12461), .A1_t (new_AGEMA_signal_12462), .A1_f (new_AGEMA_signal_12463), .B0_t (SubBytesIns_Inst_Sbox_2_L21), .B0_f (new_AGEMA_signal_13043), .B1_t (new_AGEMA_signal_13044), .B1_f (new_AGEMA_signal_13045), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .Z0_f (new_AGEMA_signal_13691), .Z1_t (new_AGEMA_signal_13692), .Z1_f (new_AGEMA_signal_13693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L20), .A0_f (new_AGEMA_signal_13040), .A1_t (new_AGEMA_signal_13041), .A1_f (new_AGEMA_signal_13042), .B0_t (SubBytesIns_Inst_Sbox_2_L22), .B0_f (new_AGEMA_signal_12479), .B1_t (new_AGEMA_signal_12480), .B1_f (new_AGEMA_signal_12481), .Z0_t (MixColumnsInput[51]), .Z0_f (new_AGEMA_signal_13694), .Z1_t (new_AGEMA_signal_13695), .Z1_f (new_AGEMA_signal_13696) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L25), .A0_f (new_AGEMA_signal_13049), .A1_t (new_AGEMA_signal_13050), .A1_f (new_AGEMA_signal_13051), .B0_t (SubBytesIns_Inst_Sbox_2_L29), .B0_f (new_AGEMA_signal_13061), .B1_t (new_AGEMA_signal_13062), .B1_f (new_AGEMA_signal_13063), .Z0_t (MixColumnsInput[50]), .Z0_f (new_AGEMA_signal_13697), .Z1_t (new_AGEMA_signal_13698), .Z1_f (new_AGEMA_signal_13699) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L13), .A0_f (new_AGEMA_signal_13034), .A1_t (new_AGEMA_signal_13035), .A1_f (new_AGEMA_signal_13036), .B0_t (SubBytesIns_Inst_Sbox_2_L27), .B0_f (new_AGEMA_signal_13055), .B1_t (new_AGEMA_signal_13056), .B1_f (new_AGEMA_signal_13057), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .Z0_f (new_AGEMA_signal_13700), .Z1_t (new_AGEMA_signal_13701), .Z1_f (new_AGEMA_signal_13702) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L6), .A0_f (new_AGEMA_signal_12461), .A1_t (new_AGEMA_signal_12462), .A1_f (new_AGEMA_signal_12463), .B0_t (SubBytesIns_Inst_Sbox_2_L23), .B0_f (new_AGEMA_signal_12482), .B1_t (new_AGEMA_signal_12483), .B1_f (new_AGEMA_signal_12484), .Z0_t (MixColumnsInput[48]), .Z0_f (new_AGEMA_signal_13064), .Z1_t (new_AGEMA_signal_13065), .Z1_f (new_AGEMA_signal_13066) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[31]), .A0_f (ciphertext_s0_f[31]), .A1_t (ciphertext_s1_t[31]), .A1_f (ciphertext_s1_f[31]), .B0_t (ciphertext_s0_t[28]), .B0_f (ciphertext_s0_f[28]), .B1_t (ciphertext_s1_t[28]), .B1_f (ciphertext_s1_f[28]), .Z0_t (SubBytesIns_Inst_Sbox_3_T1), .Z0_f (new_AGEMA_signal_6436), .Z1_t (new_AGEMA_signal_6437), .Z1_f (new_AGEMA_signal_6438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[31]), .A0_f (ciphertext_s0_f[31]), .A1_t (ciphertext_s1_t[31]), .A1_f (ciphertext_s1_f[31]), .B0_t (ciphertext_s0_t[26]), .B0_f (ciphertext_s0_f[26]), .B1_t (ciphertext_s1_t[26]), .B1_f (ciphertext_s1_f[26]), .Z0_t (SubBytesIns_Inst_Sbox_3_T2), .Z0_f (new_AGEMA_signal_6439), .Z1_t (new_AGEMA_signal_6440), .Z1_f (new_AGEMA_signal_6441) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[31]), .A0_f (ciphertext_s0_f[31]), .A1_t (ciphertext_s1_t[31]), .A1_f (ciphertext_s1_f[31]), .B0_t (ciphertext_s0_t[25]), .B0_f (ciphertext_s0_f[25]), .B1_t (ciphertext_s1_t[25]), .B1_f (ciphertext_s1_f[25]), .Z0_t (SubBytesIns_Inst_Sbox_3_T3), .Z0_f (new_AGEMA_signal_6442), .Z1_t (new_AGEMA_signal_6443), .Z1_f (new_AGEMA_signal_6444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[28]), .A0_f (ciphertext_s0_f[28]), .A1_t (ciphertext_s1_t[28]), .A1_f (ciphertext_s1_f[28]), .B0_t (ciphertext_s0_t[26]), .B0_f (ciphertext_s0_f[26]), .B1_t (ciphertext_s1_t[26]), .B1_f (ciphertext_s1_f[26]), .Z0_t (SubBytesIns_Inst_Sbox_3_T4), .Z0_f (new_AGEMA_signal_6445), .Z1_t (new_AGEMA_signal_6446), .Z1_f (new_AGEMA_signal_6447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[27]), .A0_f (ciphertext_s0_f[27]), .A1_t (ciphertext_s1_t[27]), .A1_f (ciphertext_s1_f[27]), .B0_t (ciphertext_s0_t[25]), .B0_f (ciphertext_s0_f[25]), .B1_t (ciphertext_s1_t[25]), .B1_f (ciphertext_s1_f[25]), .Z0_t (SubBytesIns_Inst_Sbox_3_T5), .Z0_f (new_AGEMA_signal_6448), .Z1_t (new_AGEMA_signal_6449), .Z1_f (new_AGEMA_signal_6450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T1), .A0_f (new_AGEMA_signal_6436), .A1_t (new_AGEMA_signal_6437), .A1_f (new_AGEMA_signal_6438), .B0_t (SubBytesIns_Inst_Sbox_3_T5), .B0_f (new_AGEMA_signal_6448), .B1_t (new_AGEMA_signal_6449), .B1_f (new_AGEMA_signal_6450), .Z0_t (SubBytesIns_Inst_Sbox_3_T6), .Z0_f (new_AGEMA_signal_7000), .Z1_t (new_AGEMA_signal_7001), .Z1_f (new_AGEMA_signal_7002) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[30]), .A0_f (ciphertext_s0_f[30]), .A1_t (ciphertext_s1_t[30]), .A1_f (ciphertext_s1_f[30]), .B0_t (ciphertext_s0_t[29]), .B0_f (ciphertext_s0_f[29]), .B1_t (ciphertext_s1_t[29]), .B1_f (ciphertext_s1_f[29]), .Z0_t (SubBytesIns_Inst_Sbox_3_T7), .Z0_f (new_AGEMA_signal_6451), .Z1_t (new_AGEMA_signal_6452), .Z1_f (new_AGEMA_signal_6453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[24]), .A0_f (ciphertext_s0_f[24]), .A1_t (ciphertext_s1_t[24]), .A1_f (ciphertext_s1_f[24]), .B0_t (SubBytesIns_Inst_Sbox_3_T6), .B0_f (new_AGEMA_signal_7000), .B1_t (new_AGEMA_signal_7001), .B1_f (new_AGEMA_signal_7002), .Z0_t (SubBytesIns_Inst_Sbox_3_T8), .Z0_f (new_AGEMA_signal_7589), .Z1_t (new_AGEMA_signal_7590), .Z1_f (new_AGEMA_signal_7591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[24]), .A0_f (ciphertext_s0_f[24]), .A1_t (ciphertext_s1_t[24]), .A1_f (ciphertext_s1_f[24]), .B0_t (SubBytesIns_Inst_Sbox_3_T7), .B0_f (new_AGEMA_signal_6451), .B1_t (new_AGEMA_signal_6452), .B1_f (new_AGEMA_signal_6453), .Z0_t (SubBytesIns_Inst_Sbox_3_T9), .Z0_f (new_AGEMA_signal_7003), .Z1_t (new_AGEMA_signal_7004), .Z1_f (new_AGEMA_signal_7005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T6), .A0_f (new_AGEMA_signal_7000), .A1_t (new_AGEMA_signal_7001), .A1_f (new_AGEMA_signal_7002), .B0_t (SubBytesIns_Inst_Sbox_3_T7), .B0_f (new_AGEMA_signal_6451), .B1_t (new_AGEMA_signal_6452), .B1_f (new_AGEMA_signal_6453), .Z0_t (SubBytesIns_Inst_Sbox_3_T10), .Z0_f (new_AGEMA_signal_7592), .Z1_t (new_AGEMA_signal_7593), .Z1_f (new_AGEMA_signal_7594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[30]), .A0_f (ciphertext_s0_f[30]), .A1_t (ciphertext_s1_t[30]), .A1_f (ciphertext_s1_f[30]), .B0_t (ciphertext_s0_t[26]), .B0_f (ciphertext_s0_f[26]), .B1_t (ciphertext_s1_t[26]), .B1_f (ciphertext_s1_f[26]), .Z0_t (SubBytesIns_Inst_Sbox_3_T11), .Z0_f (new_AGEMA_signal_6454), .Z1_t (new_AGEMA_signal_6455), .Z1_f (new_AGEMA_signal_6456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[29]), .A0_f (ciphertext_s0_f[29]), .A1_t (ciphertext_s1_t[29]), .A1_f (ciphertext_s1_f[29]), .B0_t (ciphertext_s0_t[26]), .B0_f (ciphertext_s0_f[26]), .B1_t (ciphertext_s1_t[26]), .B1_f (ciphertext_s1_f[26]), .Z0_t (SubBytesIns_Inst_Sbox_3_T12), .Z0_f (new_AGEMA_signal_6457), .Z1_t (new_AGEMA_signal_6458), .Z1_f (new_AGEMA_signal_6459) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T3), .A0_f (new_AGEMA_signal_6442), .A1_t (new_AGEMA_signal_6443), .A1_f (new_AGEMA_signal_6444), .B0_t (SubBytesIns_Inst_Sbox_3_T4), .B0_f (new_AGEMA_signal_6445), .B1_t (new_AGEMA_signal_6446), .B1_f (new_AGEMA_signal_6447), .Z0_t (SubBytesIns_Inst_Sbox_3_T13), .Z0_f (new_AGEMA_signal_7006), .Z1_t (new_AGEMA_signal_7007), .Z1_f (new_AGEMA_signal_7008) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T6), .A0_f (new_AGEMA_signal_7000), .A1_t (new_AGEMA_signal_7001), .A1_f (new_AGEMA_signal_7002), .B0_t (SubBytesIns_Inst_Sbox_3_T11), .B0_f (new_AGEMA_signal_6454), .B1_t (new_AGEMA_signal_6455), .B1_f (new_AGEMA_signal_6456), .Z0_t (SubBytesIns_Inst_Sbox_3_T14), .Z0_f (new_AGEMA_signal_7595), .Z1_t (new_AGEMA_signal_7596), .Z1_f (new_AGEMA_signal_7597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T5), .A0_f (new_AGEMA_signal_6448), .A1_t (new_AGEMA_signal_6449), .A1_f (new_AGEMA_signal_6450), .B0_t (SubBytesIns_Inst_Sbox_3_T11), .B0_f (new_AGEMA_signal_6454), .B1_t (new_AGEMA_signal_6455), .B1_f (new_AGEMA_signal_6456), .Z0_t (SubBytesIns_Inst_Sbox_3_T15), .Z0_f (new_AGEMA_signal_7009), .Z1_t (new_AGEMA_signal_7010), .Z1_f (new_AGEMA_signal_7011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T5), .A0_f (new_AGEMA_signal_6448), .A1_t (new_AGEMA_signal_6449), .A1_f (new_AGEMA_signal_6450), .B0_t (SubBytesIns_Inst_Sbox_3_T12), .B0_f (new_AGEMA_signal_6457), .B1_t (new_AGEMA_signal_6458), .B1_f (new_AGEMA_signal_6459), .Z0_t (SubBytesIns_Inst_Sbox_3_T16), .Z0_f (new_AGEMA_signal_7012), .Z1_t (new_AGEMA_signal_7013), .Z1_f (new_AGEMA_signal_7014) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T9), .A0_f (new_AGEMA_signal_7003), .A1_t (new_AGEMA_signal_7004), .A1_f (new_AGEMA_signal_7005), .B0_t (SubBytesIns_Inst_Sbox_3_T16), .B0_f (new_AGEMA_signal_7012), .B1_t (new_AGEMA_signal_7013), .B1_f (new_AGEMA_signal_7014), .Z0_t (SubBytesIns_Inst_Sbox_3_T17), .Z0_f (new_AGEMA_signal_7598), .Z1_t (new_AGEMA_signal_7599), .Z1_f (new_AGEMA_signal_7600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[28]), .A0_f (ciphertext_s0_f[28]), .A1_t (ciphertext_s1_t[28]), .A1_f (ciphertext_s1_f[28]), .B0_t (ciphertext_s0_t[24]), .B0_f (ciphertext_s0_f[24]), .B1_t (ciphertext_s1_t[24]), .B1_f (ciphertext_s1_f[24]), .Z0_t (SubBytesIns_Inst_Sbox_3_T18), .Z0_f (new_AGEMA_signal_6460), .Z1_t (new_AGEMA_signal_6461), .Z1_f (new_AGEMA_signal_6462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T7), .A0_f (new_AGEMA_signal_6451), .A1_t (new_AGEMA_signal_6452), .A1_f (new_AGEMA_signal_6453), .B0_t (SubBytesIns_Inst_Sbox_3_T18), .B0_f (new_AGEMA_signal_6460), .B1_t (new_AGEMA_signal_6461), .B1_f (new_AGEMA_signal_6462), .Z0_t (SubBytesIns_Inst_Sbox_3_T19), .Z0_f (new_AGEMA_signal_7015), .Z1_t (new_AGEMA_signal_7016), .Z1_f (new_AGEMA_signal_7017) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T1), .A0_f (new_AGEMA_signal_6436), .A1_t (new_AGEMA_signal_6437), .A1_f (new_AGEMA_signal_6438), .B0_t (SubBytesIns_Inst_Sbox_3_T19), .B0_f (new_AGEMA_signal_7015), .B1_t (new_AGEMA_signal_7016), .B1_f (new_AGEMA_signal_7017), .Z0_t (SubBytesIns_Inst_Sbox_3_T20), .Z0_f (new_AGEMA_signal_7601), .Z1_t (new_AGEMA_signal_7602), .Z1_f (new_AGEMA_signal_7603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[25]), .A0_f (ciphertext_s0_f[25]), .A1_t (ciphertext_s1_t[25]), .A1_f (ciphertext_s1_f[25]), .B0_t (ciphertext_s0_t[24]), .B0_f (ciphertext_s0_f[24]), .B1_t (ciphertext_s1_t[24]), .B1_f (ciphertext_s1_f[24]), .Z0_t (SubBytesIns_Inst_Sbox_3_T21), .Z0_f (new_AGEMA_signal_6463), .Z1_t (new_AGEMA_signal_6464), .Z1_f (new_AGEMA_signal_6465) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T7), .A0_f (new_AGEMA_signal_6451), .A1_t (new_AGEMA_signal_6452), .A1_f (new_AGEMA_signal_6453), .B0_t (SubBytesIns_Inst_Sbox_3_T21), .B0_f (new_AGEMA_signal_6463), .B1_t (new_AGEMA_signal_6464), .B1_f (new_AGEMA_signal_6465), .Z0_t (SubBytesIns_Inst_Sbox_3_T22), .Z0_f (new_AGEMA_signal_7018), .Z1_t (new_AGEMA_signal_7019), .Z1_f (new_AGEMA_signal_7020) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T2), .A0_f (new_AGEMA_signal_6439), .A1_t (new_AGEMA_signal_6440), .A1_f (new_AGEMA_signal_6441), .B0_t (SubBytesIns_Inst_Sbox_3_T22), .B0_f (new_AGEMA_signal_7018), .B1_t (new_AGEMA_signal_7019), .B1_f (new_AGEMA_signal_7020), .Z0_t (SubBytesIns_Inst_Sbox_3_T23), .Z0_f (new_AGEMA_signal_7604), .Z1_t (new_AGEMA_signal_7605), .Z1_f (new_AGEMA_signal_7606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T2), .A0_f (new_AGEMA_signal_6439), .A1_t (new_AGEMA_signal_6440), .A1_f (new_AGEMA_signal_6441), .B0_t (SubBytesIns_Inst_Sbox_3_T10), .B0_f (new_AGEMA_signal_7592), .B1_t (new_AGEMA_signal_7593), .B1_f (new_AGEMA_signal_7594), .Z0_t (SubBytesIns_Inst_Sbox_3_T24), .Z0_f (new_AGEMA_signal_8285), .Z1_t (new_AGEMA_signal_8286), .Z1_f (new_AGEMA_signal_8287) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T20), .A0_f (new_AGEMA_signal_7601), .A1_t (new_AGEMA_signal_7602), .A1_f (new_AGEMA_signal_7603), .B0_t (SubBytesIns_Inst_Sbox_3_T17), .B0_f (new_AGEMA_signal_7598), .B1_t (new_AGEMA_signal_7599), .B1_f (new_AGEMA_signal_7600), .Z0_t (SubBytesIns_Inst_Sbox_3_T25), .Z0_f (new_AGEMA_signal_8288), .Z1_t (new_AGEMA_signal_8289), .Z1_f (new_AGEMA_signal_8290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T3), .A0_f (new_AGEMA_signal_6442), .A1_t (new_AGEMA_signal_6443), .A1_f (new_AGEMA_signal_6444), .B0_t (SubBytesIns_Inst_Sbox_3_T16), .B0_f (new_AGEMA_signal_7012), .B1_t (new_AGEMA_signal_7013), .B1_f (new_AGEMA_signal_7014), .Z0_t (SubBytesIns_Inst_Sbox_3_T26), .Z0_f (new_AGEMA_signal_7607), .Z1_t (new_AGEMA_signal_7608), .Z1_f (new_AGEMA_signal_7609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T1), .A0_f (new_AGEMA_signal_6436), .A1_t (new_AGEMA_signal_6437), .A1_f (new_AGEMA_signal_6438), .B0_t (SubBytesIns_Inst_Sbox_3_T12), .B0_f (new_AGEMA_signal_6457), .B1_t (new_AGEMA_signal_6458), .B1_f (new_AGEMA_signal_6459), .Z0_t (SubBytesIns_Inst_Sbox_3_T27), .Z0_f (new_AGEMA_signal_7021), .Z1_t (new_AGEMA_signal_7022), .Z1_f (new_AGEMA_signal_7023) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T13), .A0_f (new_AGEMA_signal_7006), .A1_t (new_AGEMA_signal_7007), .A1_f (new_AGEMA_signal_7008), .B0_t (SubBytesIns_Inst_Sbox_3_T6), .B0_f (new_AGEMA_signal_7000), .B1_t (new_AGEMA_signal_7001), .B1_f (new_AGEMA_signal_7002), .Z0_t (SubBytesIns_Inst_Sbox_3_M1), .Z0_f (new_AGEMA_signal_7610), .Z1_t (new_AGEMA_signal_7611), .Z1_f (new_AGEMA_signal_7612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T23), .A0_f (new_AGEMA_signal_7604), .A1_t (new_AGEMA_signal_7605), .A1_f (new_AGEMA_signal_7606), .B0_t (SubBytesIns_Inst_Sbox_3_T8), .B0_f (new_AGEMA_signal_7589), .B1_t (new_AGEMA_signal_7590), .B1_f (new_AGEMA_signal_7591), .Z0_t (SubBytesIns_Inst_Sbox_3_M2), .Z0_f (new_AGEMA_signal_8291), .Z1_t (new_AGEMA_signal_8292), .Z1_f (new_AGEMA_signal_8293) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T14), .A0_f (new_AGEMA_signal_7595), .A1_t (new_AGEMA_signal_7596), .A1_f (new_AGEMA_signal_7597), .B0_t (SubBytesIns_Inst_Sbox_3_M1), .B0_f (new_AGEMA_signal_7610), .B1_t (new_AGEMA_signal_7611), .B1_f (new_AGEMA_signal_7612), .Z0_t (SubBytesIns_Inst_Sbox_3_M3), .Z0_f (new_AGEMA_signal_8294), .Z1_t (new_AGEMA_signal_8295), .Z1_f (new_AGEMA_signal_8296) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T19), .A0_f (new_AGEMA_signal_7015), .A1_t (new_AGEMA_signal_7016), .A1_f (new_AGEMA_signal_7017), .B0_t (ciphertext_s0_t[24]), .B0_f (ciphertext_s0_f[24]), .B1_t (ciphertext_s1_t[24]), .B1_f (ciphertext_s1_f[24]), .Z0_t (SubBytesIns_Inst_Sbox_3_M4), .Z0_f (new_AGEMA_signal_7613), .Z1_t (new_AGEMA_signal_7614), .Z1_f (new_AGEMA_signal_7615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M4), .A0_f (new_AGEMA_signal_7613), .A1_t (new_AGEMA_signal_7614), .A1_f (new_AGEMA_signal_7615), .B0_t (SubBytesIns_Inst_Sbox_3_M1), .B0_f (new_AGEMA_signal_7610), .B1_t (new_AGEMA_signal_7611), .B1_f (new_AGEMA_signal_7612), .Z0_t (SubBytesIns_Inst_Sbox_3_M5), .Z0_f (new_AGEMA_signal_8297), .Z1_t (new_AGEMA_signal_8298), .Z1_f (new_AGEMA_signal_8299) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T3), .A0_f (new_AGEMA_signal_6442), .A1_t (new_AGEMA_signal_6443), .A1_f (new_AGEMA_signal_6444), .B0_t (SubBytesIns_Inst_Sbox_3_T16), .B0_f (new_AGEMA_signal_7012), .B1_t (new_AGEMA_signal_7013), .B1_f (new_AGEMA_signal_7014), .Z0_t (SubBytesIns_Inst_Sbox_3_M6), .Z0_f (new_AGEMA_signal_7616), .Z1_t (new_AGEMA_signal_7617), .Z1_f (new_AGEMA_signal_7618) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T22), .A0_f (new_AGEMA_signal_7018), .A1_t (new_AGEMA_signal_7019), .A1_f (new_AGEMA_signal_7020), .B0_t (SubBytesIns_Inst_Sbox_3_T9), .B0_f (new_AGEMA_signal_7003), .B1_t (new_AGEMA_signal_7004), .B1_f (new_AGEMA_signal_7005), .Z0_t (SubBytesIns_Inst_Sbox_3_M7), .Z0_f (new_AGEMA_signal_7619), .Z1_t (new_AGEMA_signal_7620), .Z1_f (new_AGEMA_signal_7621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T26), .A0_f (new_AGEMA_signal_7607), .A1_t (new_AGEMA_signal_7608), .A1_f (new_AGEMA_signal_7609), .B0_t (SubBytesIns_Inst_Sbox_3_M6), .B0_f (new_AGEMA_signal_7616), .B1_t (new_AGEMA_signal_7617), .B1_f (new_AGEMA_signal_7618), .Z0_t (SubBytesIns_Inst_Sbox_3_M8), .Z0_f (new_AGEMA_signal_8300), .Z1_t (new_AGEMA_signal_8301), .Z1_f (new_AGEMA_signal_8302) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T20), .A0_f (new_AGEMA_signal_7601), .A1_t (new_AGEMA_signal_7602), .A1_f (new_AGEMA_signal_7603), .B0_t (SubBytesIns_Inst_Sbox_3_T17), .B0_f (new_AGEMA_signal_7598), .B1_t (new_AGEMA_signal_7599), .B1_f (new_AGEMA_signal_7600), .Z0_t (SubBytesIns_Inst_Sbox_3_M9), .Z0_f (new_AGEMA_signal_8303), .Z1_t (new_AGEMA_signal_8304), .Z1_f (new_AGEMA_signal_8305) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M9), .A0_f (new_AGEMA_signal_8303), .A1_t (new_AGEMA_signal_8304), .A1_f (new_AGEMA_signal_8305), .B0_t (SubBytesIns_Inst_Sbox_3_M6), .B0_f (new_AGEMA_signal_7616), .B1_t (new_AGEMA_signal_7617), .B1_f (new_AGEMA_signal_7618), .Z0_t (SubBytesIns_Inst_Sbox_3_M10), .Z0_f (new_AGEMA_signal_8741), .Z1_t (new_AGEMA_signal_8742), .Z1_f (new_AGEMA_signal_8743) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T1), .A0_f (new_AGEMA_signal_6436), .A1_t (new_AGEMA_signal_6437), .A1_f (new_AGEMA_signal_6438), .B0_t (SubBytesIns_Inst_Sbox_3_T15), .B0_f (new_AGEMA_signal_7009), .B1_t (new_AGEMA_signal_7010), .B1_f (new_AGEMA_signal_7011), .Z0_t (SubBytesIns_Inst_Sbox_3_M11), .Z0_f (new_AGEMA_signal_7622), .Z1_t (new_AGEMA_signal_7623), .Z1_f (new_AGEMA_signal_7624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T4), .A0_f (new_AGEMA_signal_6445), .A1_t (new_AGEMA_signal_6446), .A1_f (new_AGEMA_signal_6447), .B0_t (SubBytesIns_Inst_Sbox_3_T27), .B0_f (new_AGEMA_signal_7021), .B1_t (new_AGEMA_signal_7022), .B1_f (new_AGEMA_signal_7023), .Z0_t (SubBytesIns_Inst_Sbox_3_M12), .Z0_f (new_AGEMA_signal_7625), .Z1_t (new_AGEMA_signal_7626), .Z1_f (new_AGEMA_signal_7627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M12), .A0_f (new_AGEMA_signal_7625), .A1_t (new_AGEMA_signal_7626), .A1_f (new_AGEMA_signal_7627), .B0_t (SubBytesIns_Inst_Sbox_3_M11), .B0_f (new_AGEMA_signal_7622), .B1_t (new_AGEMA_signal_7623), .B1_f (new_AGEMA_signal_7624), .Z0_t (SubBytesIns_Inst_Sbox_3_M13), .Z0_f (new_AGEMA_signal_8306), .Z1_t (new_AGEMA_signal_8307), .Z1_f (new_AGEMA_signal_8308) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T2), .A0_f (new_AGEMA_signal_6439), .A1_t (new_AGEMA_signal_6440), .A1_f (new_AGEMA_signal_6441), .B0_t (SubBytesIns_Inst_Sbox_3_T10), .B0_f (new_AGEMA_signal_7592), .B1_t (new_AGEMA_signal_7593), .B1_f (new_AGEMA_signal_7594), .Z0_t (SubBytesIns_Inst_Sbox_3_M14), .Z0_f (new_AGEMA_signal_8309), .Z1_t (new_AGEMA_signal_8310), .Z1_f (new_AGEMA_signal_8311) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M14), .A0_f (new_AGEMA_signal_8309), .A1_t (new_AGEMA_signal_8310), .A1_f (new_AGEMA_signal_8311), .B0_t (SubBytesIns_Inst_Sbox_3_M11), .B0_f (new_AGEMA_signal_7622), .B1_t (new_AGEMA_signal_7623), .B1_f (new_AGEMA_signal_7624), .Z0_t (SubBytesIns_Inst_Sbox_3_M15), .Z0_f (new_AGEMA_signal_8744), .Z1_t (new_AGEMA_signal_8745), .Z1_f (new_AGEMA_signal_8746) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M3), .A0_f (new_AGEMA_signal_8294), .A1_t (new_AGEMA_signal_8295), .A1_f (new_AGEMA_signal_8296), .B0_t (SubBytesIns_Inst_Sbox_3_M2), .B0_f (new_AGEMA_signal_8291), .B1_t (new_AGEMA_signal_8292), .B1_f (new_AGEMA_signal_8293), .Z0_t (SubBytesIns_Inst_Sbox_3_M16), .Z0_f (new_AGEMA_signal_8747), .Z1_t (new_AGEMA_signal_8748), .Z1_f (new_AGEMA_signal_8749) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M5), .A0_f (new_AGEMA_signal_8297), .A1_t (new_AGEMA_signal_8298), .A1_f (new_AGEMA_signal_8299), .B0_t (SubBytesIns_Inst_Sbox_3_T24), .B0_f (new_AGEMA_signal_8285), .B1_t (new_AGEMA_signal_8286), .B1_f (new_AGEMA_signal_8287), .Z0_t (SubBytesIns_Inst_Sbox_3_M17), .Z0_f (new_AGEMA_signal_8750), .Z1_t (new_AGEMA_signal_8751), .Z1_f (new_AGEMA_signal_8752) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M8), .A0_f (new_AGEMA_signal_8300), .A1_t (new_AGEMA_signal_8301), .A1_f (new_AGEMA_signal_8302), .B0_t (SubBytesIns_Inst_Sbox_3_M7), .B0_f (new_AGEMA_signal_7619), .B1_t (new_AGEMA_signal_7620), .B1_f (new_AGEMA_signal_7621), .Z0_t (SubBytesIns_Inst_Sbox_3_M18), .Z0_f (new_AGEMA_signal_8753), .Z1_t (new_AGEMA_signal_8754), .Z1_f (new_AGEMA_signal_8755) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M10), .A0_f (new_AGEMA_signal_8741), .A1_t (new_AGEMA_signal_8742), .A1_f (new_AGEMA_signal_8743), .B0_t (SubBytesIns_Inst_Sbox_3_M15), .B0_f (new_AGEMA_signal_8744), .B1_t (new_AGEMA_signal_8745), .B1_f (new_AGEMA_signal_8746), .Z0_t (SubBytesIns_Inst_Sbox_3_M19), .Z0_f (new_AGEMA_signal_9020), .Z1_t (new_AGEMA_signal_9021), .Z1_f (new_AGEMA_signal_9022) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M16), .A0_f (new_AGEMA_signal_8747), .A1_t (new_AGEMA_signal_8748), .A1_f (new_AGEMA_signal_8749), .B0_t (SubBytesIns_Inst_Sbox_3_M13), .B0_f (new_AGEMA_signal_8306), .B1_t (new_AGEMA_signal_8307), .B1_f (new_AGEMA_signal_8308), .Z0_t (SubBytesIns_Inst_Sbox_3_M20), .Z0_f (new_AGEMA_signal_9023), .Z1_t (new_AGEMA_signal_9024), .Z1_f (new_AGEMA_signal_9025) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M17), .A0_f (new_AGEMA_signal_8750), .A1_t (new_AGEMA_signal_8751), .A1_f (new_AGEMA_signal_8752), .B0_t (SubBytesIns_Inst_Sbox_3_M15), .B0_f (new_AGEMA_signal_8744), .B1_t (new_AGEMA_signal_8745), .B1_f (new_AGEMA_signal_8746), .Z0_t (SubBytesIns_Inst_Sbox_3_M21), .Z0_f (new_AGEMA_signal_9026), .Z1_t (new_AGEMA_signal_9027), .Z1_f (new_AGEMA_signal_9028) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M18), .A0_f (new_AGEMA_signal_8753), .A1_t (new_AGEMA_signal_8754), .A1_f (new_AGEMA_signal_8755), .B0_t (SubBytesIns_Inst_Sbox_3_M13), .B0_f (new_AGEMA_signal_8306), .B1_t (new_AGEMA_signal_8307), .B1_f (new_AGEMA_signal_8308), .Z0_t (SubBytesIns_Inst_Sbox_3_M22), .Z0_f (new_AGEMA_signal_9029), .Z1_t (new_AGEMA_signal_9030), .Z1_f (new_AGEMA_signal_9031) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M19), .A0_f (new_AGEMA_signal_9020), .A1_t (new_AGEMA_signal_9021), .A1_f (new_AGEMA_signal_9022), .B0_t (SubBytesIns_Inst_Sbox_3_T25), .B0_f (new_AGEMA_signal_8288), .B1_t (new_AGEMA_signal_8289), .B1_f (new_AGEMA_signal_8290), .Z0_t (SubBytesIns_Inst_Sbox_3_M23), .Z0_f (new_AGEMA_signal_9260), .Z1_t (new_AGEMA_signal_9261), .Z1_f (new_AGEMA_signal_9262) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M22), .A0_f (new_AGEMA_signal_9029), .A1_t (new_AGEMA_signal_9030), .A1_f (new_AGEMA_signal_9031), .B0_t (SubBytesIns_Inst_Sbox_3_M23), .B0_f (new_AGEMA_signal_9260), .B1_t (new_AGEMA_signal_9261), .B1_f (new_AGEMA_signal_9262), .Z0_t (SubBytesIns_Inst_Sbox_3_M24), .Z0_f (new_AGEMA_signal_9521), .Z1_t (new_AGEMA_signal_9522), .Z1_f (new_AGEMA_signal_9523) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M22), .A0_f (new_AGEMA_signal_9029), .A1_t (new_AGEMA_signal_9030), .A1_f (new_AGEMA_signal_9031), .B0_t (SubBytesIns_Inst_Sbox_3_M20), .B0_f (new_AGEMA_signal_9023), .B1_t (new_AGEMA_signal_9024), .B1_f (new_AGEMA_signal_9025), .Z0_t (SubBytesIns_Inst_Sbox_3_M25), .Z0_f (new_AGEMA_signal_9263), .Z1_t (new_AGEMA_signal_9264), .Z1_f (new_AGEMA_signal_9265) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M21), .A0_f (new_AGEMA_signal_9026), .A1_t (new_AGEMA_signal_9027), .A1_f (new_AGEMA_signal_9028), .B0_t (SubBytesIns_Inst_Sbox_3_M25), .B0_f (new_AGEMA_signal_9263), .B1_t (new_AGEMA_signal_9264), .B1_f (new_AGEMA_signal_9265), .Z0_t (SubBytesIns_Inst_Sbox_3_M26), .Z0_f (new_AGEMA_signal_9524), .Z1_t (new_AGEMA_signal_9525), .Z1_f (new_AGEMA_signal_9526) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M20), .A0_f (new_AGEMA_signal_9023), .A1_t (new_AGEMA_signal_9024), .A1_f (new_AGEMA_signal_9025), .B0_t (SubBytesIns_Inst_Sbox_3_M21), .B0_f (new_AGEMA_signal_9026), .B1_t (new_AGEMA_signal_9027), .B1_f (new_AGEMA_signal_9028), .Z0_t (SubBytesIns_Inst_Sbox_3_M27), .Z0_f (new_AGEMA_signal_9266), .Z1_t (new_AGEMA_signal_9267), .Z1_f (new_AGEMA_signal_9268) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M23), .A0_f (new_AGEMA_signal_9260), .A1_t (new_AGEMA_signal_9261), .A1_f (new_AGEMA_signal_9262), .B0_t (SubBytesIns_Inst_Sbox_3_M25), .B0_f (new_AGEMA_signal_9263), .B1_t (new_AGEMA_signal_9264), .B1_f (new_AGEMA_signal_9265), .Z0_t (SubBytesIns_Inst_Sbox_3_M28), .Z0_f (new_AGEMA_signal_9527), .Z1_t (new_AGEMA_signal_9528), .Z1_f (new_AGEMA_signal_9529) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M28), .A0_f (new_AGEMA_signal_9527), .A1_t (new_AGEMA_signal_9528), .A1_f (new_AGEMA_signal_9529), .B0_t (SubBytesIns_Inst_Sbox_3_M27), .B0_f (new_AGEMA_signal_9266), .B1_t (new_AGEMA_signal_9267), .B1_f (new_AGEMA_signal_9268), .Z0_t (SubBytesIns_Inst_Sbox_3_M29), .Z0_f (new_AGEMA_signal_9821), .Z1_t (new_AGEMA_signal_9822), .Z1_f (new_AGEMA_signal_9823) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M26), .A0_f (new_AGEMA_signal_9524), .A1_t (new_AGEMA_signal_9525), .A1_f (new_AGEMA_signal_9526), .B0_t (SubBytesIns_Inst_Sbox_3_M24), .B0_f (new_AGEMA_signal_9521), .B1_t (new_AGEMA_signal_9522), .B1_f (new_AGEMA_signal_9523), .Z0_t (SubBytesIns_Inst_Sbox_3_M30), .Z0_f (new_AGEMA_signal_9824), .Z1_t (new_AGEMA_signal_9825), .Z1_f (new_AGEMA_signal_9826) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M20), .A0_f (new_AGEMA_signal_9023), .A1_t (new_AGEMA_signal_9024), .A1_f (new_AGEMA_signal_9025), .B0_t (SubBytesIns_Inst_Sbox_3_M23), .B0_f (new_AGEMA_signal_9260), .B1_t (new_AGEMA_signal_9261), .B1_f (new_AGEMA_signal_9262), .Z0_t (SubBytesIns_Inst_Sbox_3_M31), .Z0_f (new_AGEMA_signal_9530), .Z1_t (new_AGEMA_signal_9531), .Z1_f (new_AGEMA_signal_9532) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M27), .A0_f (new_AGEMA_signal_9266), .A1_t (new_AGEMA_signal_9267), .A1_f (new_AGEMA_signal_9268), .B0_t (SubBytesIns_Inst_Sbox_3_M31), .B0_f (new_AGEMA_signal_9530), .B1_t (new_AGEMA_signal_9531), .B1_f (new_AGEMA_signal_9532), .Z0_t (SubBytesIns_Inst_Sbox_3_M32), .Z0_f (new_AGEMA_signal_9827), .Z1_t (new_AGEMA_signal_9828), .Z1_f (new_AGEMA_signal_9829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M27), .A0_f (new_AGEMA_signal_9266), .A1_t (new_AGEMA_signal_9267), .A1_f (new_AGEMA_signal_9268), .B0_t (SubBytesIns_Inst_Sbox_3_M25), .B0_f (new_AGEMA_signal_9263), .B1_t (new_AGEMA_signal_9264), .B1_f (new_AGEMA_signal_9265), .Z0_t (SubBytesIns_Inst_Sbox_3_M33), .Z0_f (new_AGEMA_signal_9533), .Z1_t (new_AGEMA_signal_9534), .Z1_f (new_AGEMA_signal_9535) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M21), .A0_f (new_AGEMA_signal_9026), .A1_t (new_AGEMA_signal_9027), .A1_f (new_AGEMA_signal_9028), .B0_t (SubBytesIns_Inst_Sbox_3_M22), .B0_f (new_AGEMA_signal_9029), .B1_t (new_AGEMA_signal_9030), .B1_f (new_AGEMA_signal_9031), .Z0_t (SubBytesIns_Inst_Sbox_3_M34), .Z0_f (new_AGEMA_signal_9269), .Z1_t (new_AGEMA_signal_9270), .Z1_f (new_AGEMA_signal_9271) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M24), .A0_f (new_AGEMA_signal_9521), .A1_t (new_AGEMA_signal_9522), .A1_f (new_AGEMA_signal_9523), .B0_t (SubBytesIns_Inst_Sbox_3_M34), .B0_f (new_AGEMA_signal_9269), .B1_t (new_AGEMA_signal_9270), .B1_f (new_AGEMA_signal_9271), .Z0_t (SubBytesIns_Inst_Sbox_3_M35), .Z0_f (new_AGEMA_signal_9830), .Z1_t (new_AGEMA_signal_9831), .Z1_f (new_AGEMA_signal_9832) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M24), .A0_f (new_AGEMA_signal_9521), .A1_t (new_AGEMA_signal_9522), .A1_f (new_AGEMA_signal_9523), .B0_t (SubBytesIns_Inst_Sbox_3_M25), .B0_f (new_AGEMA_signal_9263), .B1_t (new_AGEMA_signal_9264), .B1_f (new_AGEMA_signal_9265), .Z0_t (SubBytesIns_Inst_Sbox_3_M36), .Z0_f (new_AGEMA_signal_9833), .Z1_t (new_AGEMA_signal_9834), .Z1_f (new_AGEMA_signal_9835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M21), .A0_f (new_AGEMA_signal_9026), .A1_t (new_AGEMA_signal_9027), .A1_f (new_AGEMA_signal_9028), .B0_t (SubBytesIns_Inst_Sbox_3_M29), .B0_f (new_AGEMA_signal_9821), .B1_t (new_AGEMA_signal_9822), .B1_f (new_AGEMA_signal_9823), .Z0_t (SubBytesIns_Inst_Sbox_3_M37), .Z0_f (new_AGEMA_signal_10100), .Z1_t (new_AGEMA_signal_10101), .Z1_f (new_AGEMA_signal_10102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M32), .A0_f (new_AGEMA_signal_9827), .A1_t (new_AGEMA_signal_9828), .A1_f (new_AGEMA_signal_9829), .B0_t (SubBytesIns_Inst_Sbox_3_M33), .B0_f (new_AGEMA_signal_9533), .B1_t (new_AGEMA_signal_9534), .B1_f (new_AGEMA_signal_9535), .Z0_t (SubBytesIns_Inst_Sbox_3_M38), .Z0_f (new_AGEMA_signal_10103), .Z1_t (new_AGEMA_signal_10104), .Z1_f (new_AGEMA_signal_10105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M23), .A0_f (new_AGEMA_signal_9260), .A1_t (new_AGEMA_signal_9261), .A1_f (new_AGEMA_signal_9262), .B0_t (SubBytesIns_Inst_Sbox_3_M30), .B0_f (new_AGEMA_signal_9824), .B1_t (new_AGEMA_signal_9825), .B1_f (new_AGEMA_signal_9826), .Z0_t (SubBytesIns_Inst_Sbox_3_M39), .Z0_f (new_AGEMA_signal_10106), .Z1_t (new_AGEMA_signal_10107), .Z1_f (new_AGEMA_signal_10108) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M35), .A0_f (new_AGEMA_signal_9830), .A1_t (new_AGEMA_signal_9831), .A1_f (new_AGEMA_signal_9832), .B0_t (SubBytesIns_Inst_Sbox_3_M36), .B0_f (new_AGEMA_signal_9833), .B1_t (new_AGEMA_signal_9834), .B1_f (new_AGEMA_signal_9835), .Z0_t (SubBytesIns_Inst_Sbox_3_M40), .Z0_f (new_AGEMA_signal_10109), .Z1_t (new_AGEMA_signal_10110), .Z1_f (new_AGEMA_signal_10111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M38), .A0_f (new_AGEMA_signal_10103), .A1_t (new_AGEMA_signal_10104), .A1_f (new_AGEMA_signal_10105), .B0_t (SubBytesIns_Inst_Sbox_3_M40), .B0_f (new_AGEMA_signal_10109), .B1_t (new_AGEMA_signal_10110), .B1_f (new_AGEMA_signal_10111), .Z0_t (SubBytesIns_Inst_Sbox_3_M41), .Z0_f (new_AGEMA_signal_10508), .Z1_t (new_AGEMA_signal_10509), .Z1_f (new_AGEMA_signal_10510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M37), .A0_f (new_AGEMA_signal_10100), .A1_t (new_AGEMA_signal_10101), .A1_f (new_AGEMA_signal_10102), .B0_t (SubBytesIns_Inst_Sbox_3_M39), .B0_f (new_AGEMA_signal_10106), .B1_t (new_AGEMA_signal_10107), .B1_f (new_AGEMA_signal_10108), .Z0_t (SubBytesIns_Inst_Sbox_3_M42), .Z0_f (new_AGEMA_signal_10511), .Z1_t (new_AGEMA_signal_10512), .Z1_f (new_AGEMA_signal_10513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M37), .A0_f (new_AGEMA_signal_10100), .A1_t (new_AGEMA_signal_10101), .A1_f (new_AGEMA_signal_10102), .B0_t (SubBytesIns_Inst_Sbox_3_M38), .B0_f (new_AGEMA_signal_10103), .B1_t (new_AGEMA_signal_10104), .B1_f (new_AGEMA_signal_10105), .Z0_t (SubBytesIns_Inst_Sbox_3_M43), .Z0_f (new_AGEMA_signal_10514), .Z1_t (new_AGEMA_signal_10515), .Z1_f (new_AGEMA_signal_10516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M39), .A0_f (new_AGEMA_signal_10106), .A1_t (new_AGEMA_signal_10107), .A1_f (new_AGEMA_signal_10108), .B0_t (SubBytesIns_Inst_Sbox_3_M40), .B0_f (new_AGEMA_signal_10109), .B1_t (new_AGEMA_signal_10110), .B1_f (new_AGEMA_signal_10111), .Z0_t (SubBytesIns_Inst_Sbox_3_M44), .Z0_f (new_AGEMA_signal_10517), .Z1_t (new_AGEMA_signal_10518), .Z1_f (new_AGEMA_signal_10519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M42), .A0_f (new_AGEMA_signal_10511), .A1_t (new_AGEMA_signal_10512), .A1_f (new_AGEMA_signal_10513), .B0_t (SubBytesIns_Inst_Sbox_3_M41), .B0_f (new_AGEMA_signal_10508), .B1_t (new_AGEMA_signal_10509), .B1_f (new_AGEMA_signal_10510), .Z0_t (SubBytesIns_Inst_Sbox_3_M45), .Z0_f (new_AGEMA_signal_11228), .Z1_t (new_AGEMA_signal_11229), .Z1_f (new_AGEMA_signal_11230) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M44), .A0_f (new_AGEMA_signal_10517), .A1_t (new_AGEMA_signal_10518), .A1_f (new_AGEMA_signal_10519), .B0_t (SubBytesIns_Inst_Sbox_3_T6), .B0_f (new_AGEMA_signal_7000), .B1_t (new_AGEMA_signal_7001), .B1_f (new_AGEMA_signal_7002), .Z0_t (SubBytesIns_Inst_Sbox_3_M46), .Z0_f (new_AGEMA_signal_11231), .Z1_t (new_AGEMA_signal_11232), .Z1_f (new_AGEMA_signal_11233) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M40), .A0_f (new_AGEMA_signal_10109), .A1_t (new_AGEMA_signal_10110), .A1_f (new_AGEMA_signal_10111), .B0_t (SubBytesIns_Inst_Sbox_3_T8), .B0_f (new_AGEMA_signal_7589), .B1_t (new_AGEMA_signal_7590), .B1_f (new_AGEMA_signal_7591), .Z0_t (SubBytesIns_Inst_Sbox_3_M47), .Z0_f (new_AGEMA_signal_10520), .Z1_t (new_AGEMA_signal_10521), .Z1_f (new_AGEMA_signal_10522) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M39), .A0_f (new_AGEMA_signal_10106), .A1_t (new_AGEMA_signal_10107), .A1_f (new_AGEMA_signal_10108), .B0_t (ciphertext_s0_t[24]), .B0_f (ciphertext_s0_f[24]), .B1_t (ciphertext_s1_t[24]), .B1_f (ciphertext_s1_f[24]), .Z0_t (SubBytesIns_Inst_Sbox_3_M48), .Z0_f (new_AGEMA_signal_10523), .Z1_t (new_AGEMA_signal_10524), .Z1_f (new_AGEMA_signal_10525) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M43), .A0_f (new_AGEMA_signal_10514), .A1_t (new_AGEMA_signal_10515), .A1_f (new_AGEMA_signal_10516), .B0_t (SubBytesIns_Inst_Sbox_3_T16), .B0_f (new_AGEMA_signal_7012), .B1_t (new_AGEMA_signal_7013), .B1_f (new_AGEMA_signal_7014), .Z0_t (SubBytesIns_Inst_Sbox_3_M49), .Z0_f (new_AGEMA_signal_11234), .Z1_t (new_AGEMA_signal_11235), .Z1_f (new_AGEMA_signal_11236) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M38), .A0_f (new_AGEMA_signal_10103), .A1_t (new_AGEMA_signal_10104), .A1_f (new_AGEMA_signal_10105), .B0_t (SubBytesIns_Inst_Sbox_3_T9), .B0_f (new_AGEMA_signal_7003), .B1_t (new_AGEMA_signal_7004), .B1_f (new_AGEMA_signal_7005), .Z0_t (SubBytesIns_Inst_Sbox_3_M50), .Z0_f (new_AGEMA_signal_10526), .Z1_t (new_AGEMA_signal_10527), .Z1_f (new_AGEMA_signal_10528) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M37), .A0_f (new_AGEMA_signal_10100), .A1_t (new_AGEMA_signal_10101), .A1_f (new_AGEMA_signal_10102), .B0_t (SubBytesIns_Inst_Sbox_3_T17), .B0_f (new_AGEMA_signal_7598), .B1_t (new_AGEMA_signal_7599), .B1_f (new_AGEMA_signal_7600), .Z0_t (SubBytesIns_Inst_Sbox_3_M51), .Z0_f (new_AGEMA_signal_10529), .Z1_t (new_AGEMA_signal_10530), .Z1_f (new_AGEMA_signal_10531) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M42), .A0_f (new_AGEMA_signal_10511), .A1_t (new_AGEMA_signal_10512), .A1_f (new_AGEMA_signal_10513), .B0_t (SubBytesIns_Inst_Sbox_3_T15), .B0_f (new_AGEMA_signal_7009), .B1_t (new_AGEMA_signal_7010), .B1_f (new_AGEMA_signal_7011), .Z0_t (SubBytesIns_Inst_Sbox_3_M52), .Z0_f (new_AGEMA_signal_11237), .Z1_t (new_AGEMA_signal_11238), .Z1_f (new_AGEMA_signal_11239) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M45), .A0_f (new_AGEMA_signal_11228), .A1_t (new_AGEMA_signal_11229), .A1_f (new_AGEMA_signal_11230), .B0_t (SubBytesIns_Inst_Sbox_3_T27), .B0_f (new_AGEMA_signal_7021), .B1_t (new_AGEMA_signal_7022), .B1_f (new_AGEMA_signal_7023), .Z0_t (SubBytesIns_Inst_Sbox_3_M53), .Z0_f (new_AGEMA_signal_11906), .Z1_t (new_AGEMA_signal_11907), .Z1_f (new_AGEMA_signal_11908) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M41), .A0_f (new_AGEMA_signal_10508), .A1_t (new_AGEMA_signal_10509), .A1_f (new_AGEMA_signal_10510), .B0_t (SubBytesIns_Inst_Sbox_3_T10), .B0_f (new_AGEMA_signal_7592), .B1_t (new_AGEMA_signal_7593), .B1_f (new_AGEMA_signal_7594), .Z0_t (SubBytesIns_Inst_Sbox_3_M54), .Z0_f (new_AGEMA_signal_11240), .Z1_t (new_AGEMA_signal_11241), .Z1_f (new_AGEMA_signal_11242) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M44), .A0_f (new_AGEMA_signal_10517), .A1_t (new_AGEMA_signal_10518), .A1_f (new_AGEMA_signal_10519), .B0_t (SubBytesIns_Inst_Sbox_3_T13), .B0_f (new_AGEMA_signal_7006), .B1_t (new_AGEMA_signal_7007), .B1_f (new_AGEMA_signal_7008), .Z0_t (SubBytesIns_Inst_Sbox_3_M55), .Z0_f (new_AGEMA_signal_11243), .Z1_t (new_AGEMA_signal_11244), .Z1_f (new_AGEMA_signal_11245) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M40), .A0_f (new_AGEMA_signal_10109), .A1_t (new_AGEMA_signal_10110), .A1_f (new_AGEMA_signal_10111), .B0_t (SubBytesIns_Inst_Sbox_3_T23), .B0_f (new_AGEMA_signal_7604), .B1_t (new_AGEMA_signal_7605), .B1_f (new_AGEMA_signal_7606), .Z0_t (SubBytesIns_Inst_Sbox_3_M56), .Z0_f (new_AGEMA_signal_10532), .Z1_t (new_AGEMA_signal_10533), .Z1_f (new_AGEMA_signal_10534) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M39), .A0_f (new_AGEMA_signal_10106), .A1_t (new_AGEMA_signal_10107), .A1_f (new_AGEMA_signal_10108), .B0_t (SubBytesIns_Inst_Sbox_3_T19), .B0_f (new_AGEMA_signal_7015), .B1_t (new_AGEMA_signal_7016), .B1_f (new_AGEMA_signal_7017), .Z0_t (SubBytesIns_Inst_Sbox_3_M57), .Z0_f (new_AGEMA_signal_10535), .Z1_t (new_AGEMA_signal_10536), .Z1_f (new_AGEMA_signal_10537) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M43), .A0_f (new_AGEMA_signal_10514), .A1_t (new_AGEMA_signal_10515), .A1_f (new_AGEMA_signal_10516), .B0_t (SubBytesIns_Inst_Sbox_3_T3), .B0_f (new_AGEMA_signal_6442), .B1_t (new_AGEMA_signal_6443), .B1_f (new_AGEMA_signal_6444), .Z0_t (SubBytesIns_Inst_Sbox_3_M58), .Z0_f (new_AGEMA_signal_11246), .Z1_t (new_AGEMA_signal_11247), .Z1_f (new_AGEMA_signal_11248) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M38), .A0_f (new_AGEMA_signal_10103), .A1_t (new_AGEMA_signal_10104), .A1_f (new_AGEMA_signal_10105), .B0_t (SubBytesIns_Inst_Sbox_3_T22), .B0_f (new_AGEMA_signal_7018), .B1_t (new_AGEMA_signal_7019), .B1_f (new_AGEMA_signal_7020), .Z0_t (SubBytesIns_Inst_Sbox_3_M59), .Z0_f (new_AGEMA_signal_10538), .Z1_t (new_AGEMA_signal_10539), .Z1_f (new_AGEMA_signal_10540) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M37), .A0_f (new_AGEMA_signal_10100), .A1_t (new_AGEMA_signal_10101), .A1_f (new_AGEMA_signal_10102), .B0_t (SubBytesIns_Inst_Sbox_3_T20), .B0_f (new_AGEMA_signal_7601), .B1_t (new_AGEMA_signal_7602), .B1_f (new_AGEMA_signal_7603), .Z0_t (SubBytesIns_Inst_Sbox_3_M60), .Z0_f (new_AGEMA_signal_10541), .Z1_t (new_AGEMA_signal_10542), .Z1_f (new_AGEMA_signal_10543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M42), .A0_f (new_AGEMA_signal_10511), .A1_t (new_AGEMA_signal_10512), .A1_f (new_AGEMA_signal_10513), .B0_t (SubBytesIns_Inst_Sbox_3_T1), .B0_f (new_AGEMA_signal_6436), .B1_t (new_AGEMA_signal_6437), .B1_f (new_AGEMA_signal_6438), .Z0_t (SubBytesIns_Inst_Sbox_3_M61), .Z0_f (new_AGEMA_signal_11249), .Z1_t (new_AGEMA_signal_11250), .Z1_f (new_AGEMA_signal_11251) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M45), .A0_f (new_AGEMA_signal_11228), .A1_t (new_AGEMA_signal_11229), .A1_f (new_AGEMA_signal_11230), .B0_t (SubBytesIns_Inst_Sbox_3_T4), .B0_f (new_AGEMA_signal_6445), .B1_t (new_AGEMA_signal_6446), .B1_f (new_AGEMA_signal_6447), .Z0_t (SubBytesIns_Inst_Sbox_3_M62), .Z0_f (new_AGEMA_signal_11909), .Z1_t (new_AGEMA_signal_11910), .Z1_f (new_AGEMA_signal_11911) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M41), .A0_f (new_AGEMA_signal_10508), .A1_t (new_AGEMA_signal_10509), .A1_f (new_AGEMA_signal_10510), .B0_t (SubBytesIns_Inst_Sbox_3_T2), .B0_f (new_AGEMA_signal_6439), .B1_t (new_AGEMA_signal_6440), .B1_f (new_AGEMA_signal_6441), .Z0_t (SubBytesIns_Inst_Sbox_3_M63), .Z0_f (new_AGEMA_signal_11252), .Z1_t (new_AGEMA_signal_11253), .Z1_f (new_AGEMA_signal_11254) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M61), .A0_f (new_AGEMA_signal_11249), .A1_t (new_AGEMA_signal_11250), .A1_f (new_AGEMA_signal_11251), .B0_t (SubBytesIns_Inst_Sbox_3_M62), .B0_f (new_AGEMA_signal_11909), .B1_t (new_AGEMA_signal_11910), .B1_f (new_AGEMA_signal_11911), .Z0_t (SubBytesIns_Inst_Sbox_3_L0), .Z0_f (new_AGEMA_signal_12485), .Z1_t (new_AGEMA_signal_12486), .Z1_f (new_AGEMA_signal_12487) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M50), .A0_f (new_AGEMA_signal_10526), .A1_t (new_AGEMA_signal_10527), .A1_f (new_AGEMA_signal_10528), .B0_t (SubBytesIns_Inst_Sbox_3_M56), .B0_f (new_AGEMA_signal_10532), .B1_t (new_AGEMA_signal_10533), .B1_f (new_AGEMA_signal_10534), .Z0_t (SubBytesIns_Inst_Sbox_3_L1), .Z0_f (new_AGEMA_signal_11255), .Z1_t (new_AGEMA_signal_11256), .Z1_f (new_AGEMA_signal_11257) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M46), .A0_f (new_AGEMA_signal_11231), .A1_t (new_AGEMA_signal_11232), .A1_f (new_AGEMA_signal_11233), .B0_t (SubBytesIns_Inst_Sbox_3_M48), .B0_f (new_AGEMA_signal_10523), .B1_t (new_AGEMA_signal_10524), .B1_f (new_AGEMA_signal_10525), .Z0_t (SubBytesIns_Inst_Sbox_3_L2), .Z0_f (new_AGEMA_signal_11912), .Z1_t (new_AGEMA_signal_11913), .Z1_f (new_AGEMA_signal_11914) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M47), .A0_f (new_AGEMA_signal_10520), .A1_t (new_AGEMA_signal_10521), .A1_f (new_AGEMA_signal_10522), .B0_t (SubBytesIns_Inst_Sbox_3_M55), .B0_f (new_AGEMA_signal_11243), .B1_t (new_AGEMA_signal_11244), .B1_f (new_AGEMA_signal_11245), .Z0_t (SubBytesIns_Inst_Sbox_3_L3), .Z0_f (new_AGEMA_signal_11915), .Z1_t (new_AGEMA_signal_11916), .Z1_f (new_AGEMA_signal_11917) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M54), .A0_f (new_AGEMA_signal_11240), .A1_t (new_AGEMA_signal_11241), .A1_f (new_AGEMA_signal_11242), .B0_t (SubBytesIns_Inst_Sbox_3_M58), .B0_f (new_AGEMA_signal_11246), .B1_t (new_AGEMA_signal_11247), .B1_f (new_AGEMA_signal_11248), .Z0_t (SubBytesIns_Inst_Sbox_3_L4), .Z0_f (new_AGEMA_signal_11918), .Z1_t (new_AGEMA_signal_11919), .Z1_f (new_AGEMA_signal_11920) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M49), .A0_f (new_AGEMA_signal_11234), .A1_t (new_AGEMA_signal_11235), .A1_f (new_AGEMA_signal_11236), .B0_t (SubBytesIns_Inst_Sbox_3_M61), .B0_f (new_AGEMA_signal_11249), .B1_t (new_AGEMA_signal_11250), .B1_f (new_AGEMA_signal_11251), .Z0_t (SubBytesIns_Inst_Sbox_3_L5), .Z0_f (new_AGEMA_signal_11921), .Z1_t (new_AGEMA_signal_11922), .Z1_f (new_AGEMA_signal_11923) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M62), .A0_f (new_AGEMA_signal_11909), .A1_t (new_AGEMA_signal_11910), .A1_f (new_AGEMA_signal_11911), .B0_t (SubBytesIns_Inst_Sbox_3_L5), .B0_f (new_AGEMA_signal_11921), .B1_t (new_AGEMA_signal_11922), .B1_f (new_AGEMA_signal_11923), .Z0_t (SubBytesIns_Inst_Sbox_3_L6), .Z0_f (new_AGEMA_signal_12488), .Z1_t (new_AGEMA_signal_12489), .Z1_f (new_AGEMA_signal_12490) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M46), .A0_f (new_AGEMA_signal_11231), .A1_t (new_AGEMA_signal_11232), .A1_f (new_AGEMA_signal_11233), .B0_t (SubBytesIns_Inst_Sbox_3_L3), .B0_f (new_AGEMA_signal_11915), .B1_t (new_AGEMA_signal_11916), .B1_f (new_AGEMA_signal_11917), .Z0_t (SubBytesIns_Inst_Sbox_3_L7), .Z0_f (new_AGEMA_signal_12491), .Z1_t (new_AGEMA_signal_12492), .Z1_f (new_AGEMA_signal_12493) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M51), .A0_f (new_AGEMA_signal_10529), .A1_t (new_AGEMA_signal_10530), .A1_f (new_AGEMA_signal_10531), .B0_t (SubBytesIns_Inst_Sbox_3_M59), .B0_f (new_AGEMA_signal_10538), .B1_t (new_AGEMA_signal_10539), .B1_f (new_AGEMA_signal_10540), .Z0_t (SubBytesIns_Inst_Sbox_3_L8), .Z0_f (new_AGEMA_signal_11258), .Z1_t (new_AGEMA_signal_11259), .Z1_f (new_AGEMA_signal_11260) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M52), .A0_f (new_AGEMA_signal_11237), .A1_t (new_AGEMA_signal_11238), .A1_f (new_AGEMA_signal_11239), .B0_t (SubBytesIns_Inst_Sbox_3_M53), .B0_f (new_AGEMA_signal_11906), .B1_t (new_AGEMA_signal_11907), .B1_f (new_AGEMA_signal_11908), .Z0_t (SubBytesIns_Inst_Sbox_3_L9), .Z0_f (new_AGEMA_signal_12494), .Z1_t (new_AGEMA_signal_12495), .Z1_f (new_AGEMA_signal_12496) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M53), .A0_f (new_AGEMA_signal_11906), .A1_t (new_AGEMA_signal_11907), .A1_f (new_AGEMA_signal_11908), .B0_t (SubBytesIns_Inst_Sbox_3_L4), .B0_f (new_AGEMA_signal_11918), .B1_t (new_AGEMA_signal_11919), .B1_f (new_AGEMA_signal_11920), .Z0_t (SubBytesIns_Inst_Sbox_3_L10), .Z0_f (new_AGEMA_signal_12497), .Z1_t (new_AGEMA_signal_12498), .Z1_f (new_AGEMA_signal_12499) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M60), .A0_f (new_AGEMA_signal_10541), .A1_t (new_AGEMA_signal_10542), .A1_f (new_AGEMA_signal_10543), .B0_t (SubBytesIns_Inst_Sbox_3_L2), .B0_f (new_AGEMA_signal_11912), .B1_t (new_AGEMA_signal_11913), .B1_f (new_AGEMA_signal_11914), .Z0_t (SubBytesIns_Inst_Sbox_3_L11), .Z0_f (new_AGEMA_signal_12500), .Z1_t (new_AGEMA_signal_12501), .Z1_f (new_AGEMA_signal_12502) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M48), .A0_f (new_AGEMA_signal_10523), .A1_t (new_AGEMA_signal_10524), .A1_f (new_AGEMA_signal_10525), .B0_t (SubBytesIns_Inst_Sbox_3_M51), .B0_f (new_AGEMA_signal_10529), .B1_t (new_AGEMA_signal_10530), .B1_f (new_AGEMA_signal_10531), .Z0_t (SubBytesIns_Inst_Sbox_3_L12), .Z0_f (new_AGEMA_signal_11261), .Z1_t (new_AGEMA_signal_11262), .Z1_f (new_AGEMA_signal_11263) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M50), .A0_f (new_AGEMA_signal_10526), .A1_t (new_AGEMA_signal_10527), .A1_f (new_AGEMA_signal_10528), .B0_t (SubBytesIns_Inst_Sbox_3_L0), .B0_f (new_AGEMA_signal_12485), .B1_t (new_AGEMA_signal_12486), .B1_f (new_AGEMA_signal_12487), .Z0_t (SubBytesIns_Inst_Sbox_3_L13), .Z0_f (new_AGEMA_signal_13067), .Z1_t (new_AGEMA_signal_13068), .Z1_f (new_AGEMA_signal_13069) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M52), .A0_f (new_AGEMA_signal_11237), .A1_t (new_AGEMA_signal_11238), .A1_f (new_AGEMA_signal_11239), .B0_t (SubBytesIns_Inst_Sbox_3_M61), .B0_f (new_AGEMA_signal_11249), .B1_t (new_AGEMA_signal_11250), .B1_f (new_AGEMA_signal_11251), .Z0_t (SubBytesIns_Inst_Sbox_3_L14), .Z0_f (new_AGEMA_signal_11924), .Z1_t (new_AGEMA_signal_11925), .Z1_f (new_AGEMA_signal_11926) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M55), .A0_f (new_AGEMA_signal_11243), .A1_t (new_AGEMA_signal_11244), .A1_f (new_AGEMA_signal_11245), .B0_t (SubBytesIns_Inst_Sbox_3_L1), .B0_f (new_AGEMA_signal_11255), .B1_t (new_AGEMA_signal_11256), .B1_f (new_AGEMA_signal_11257), .Z0_t (SubBytesIns_Inst_Sbox_3_L15), .Z0_f (new_AGEMA_signal_11927), .Z1_t (new_AGEMA_signal_11928), .Z1_f (new_AGEMA_signal_11929) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M56), .A0_f (new_AGEMA_signal_10532), .A1_t (new_AGEMA_signal_10533), .A1_f (new_AGEMA_signal_10534), .B0_t (SubBytesIns_Inst_Sbox_3_L0), .B0_f (new_AGEMA_signal_12485), .B1_t (new_AGEMA_signal_12486), .B1_f (new_AGEMA_signal_12487), .Z0_t (SubBytesIns_Inst_Sbox_3_L16), .Z0_f (new_AGEMA_signal_13070), .Z1_t (new_AGEMA_signal_13071), .Z1_f (new_AGEMA_signal_13072) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M57), .A0_f (new_AGEMA_signal_10535), .A1_t (new_AGEMA_signal_10536), .A1_f (new_AGEMA_signal_10537), .B0_t (SubBytesIns_Inst_Sbox_3_L1), .B0_f (new_AGEMA_signal_11255), .B1_t (new_AGEMA_signal_11256), .B1_f (new_AGEMA_signal_11257), .Z0_t (SubBytesIns_Inst_Sbox_3_L17), .Z0_f (new_AGEMA_signal_11930), .Z1_t (new_AGEMA_signal_11931), .Z1_f (new_AGEMA_signal_11932) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M58), .A0_f (new_AGEMA_signal_11246), .A1_t (new_AGEMA_signal_11247), .A1_f (new_AGEMA_signal_11248), .B0_t (SubBytesIns_Inst_Sbox_3_L8), .B0_f (new_AGEMA_signal_11258), .B1_t (new_AGEMA_signal_11259), .B1_f (new_AGEMA_signal_11260), .Z0_t (SubBytesIns_Inst_Sbox_3_L18), .Z0_f (new_AGEMA_signal_11933), .Z1_t (new_AGEMA_signal_11934), .Z1_f (new_AGEMA_signal_11935) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M63), .A0_f (new_AGEMA_signal_11252), .A1_t (new_AGEMA_signal_11253), .A1_f (new_AGEMA_signal_11254), .B0_t (SubBytesIns_Inst_Sbox_3_L4), .B0_f (new_AGEMA_signal_11918), .B1_t (new_AGEMA_signal_11919), .B1_f (new_AGEMA_signal_11920), .Z0_t (SubBytesIns_Inst_Sbox_3_L19), .Z0_f (new_AGEMA_signal_12503), .Z1_t (new_AGEMA_signal_12504), .Z1_f (new_AGEMA_signal_12505) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L0), .A0_f (new_AGEMA_signal_12485), .A1_t (new_AGEMA_signal_12486), .A1_f (new_AGEMA_signal_12487), .B0_t (SubBytesIns_Inst_Sbox_3_L1), .B0_f (new_AGEMA_signal_11255), .B1_t (new_AGEMA_signal_11256), .B1_f (new_AGEMA_signal_11257), .Z0_t (SubBytesIns_Inst_Sbox_3_L20), .Z0_f (new_AGEMA_signal_13073), .Z1_t (new_AGEMA_signal_13074), .Z1_f (new_AGEMA_signal_13075) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L1), .A0_f (new_AGEMA_signal_11255), .A1_t (new_AGEMA_signal_11256), .A1_f (new_AGEMA_signal_11257), .B0_t (SubBytesIns_Inst_Sbox_3_L7), .B0_f (new_AGEMA_signal_12491), .B1_t (new_AGEMA_signal_12492), .B1_f (new_AGEMA_signal_12493), .Z0_t (SubBytesIns_Inst_Sbox_3_L21), .Z0_f (new_AGEMA_signal_13076), .Z1_t (new_AGEMA_signal_13077), .Z1_f (new_AGEMA_signal_13078) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L3), .A0_f (new_AGEMA_signal_11915), .A1_t (new_AGEMA_signal_11916), .A1_f (new_AGEMA_signal_11917), .B0_t (SubBytesIns_Inst_Sbox_3_L12), .B0_f (new_AGEMA_signal_11261), .B1_t (new_AGEMA_signal_11262), .B1_f (new_AGEMA_signal_11263), .Z0_t (SubBytesIns_Inst_Sbox_3_L22), .Z0_f (new_AGEMA_signal_12506), .Z1_t (new_AGEMA_signal_12507), .Z1_f (new_AGEMA_signal_12508) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L18), .A0_f (new_AGEMA_signal_11933), .A1_t (new_AGEMA_signal_11934), .A1_f (new_AGEMA_signal_11935), .B0_t (SubBytesIns_Inst_Sbox_3_L2), .B0_f (new_AGEMA_signal_11912), .B1_t (new_AGEMA_signal_11913), .B1_f (new_AGEMA_signal_11914), .Z0_t (SubBytesIns_Inst_Sbox_3_L23), .Z0_f (new_AGEMA_signal_12509), .Z1_t (new_AGEMA_signal_12510), .Z1_f (new_AGEMA_signal_12511) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L15), .A0_f (new_AGEMA_signal_11927), .A1_t (new_AGEMA_signal_11928), .A1_f (new_AGEMA_signal_11929), .B0_t (SubBytesIns_Inst_Sbox_3_L9), .B0_f (new_AGEMA_signal_12494), .B1_t (new_AGEMA_signal_12495), .B1_f (new_AGEMA_signal_12496), .Z0_t (SubBytesIns_Inst_Sbox_3_L24), .Z0_f (new_AGEMA_signal_13079), .Z1_t (new_AGEMA_signal_13080), .Z1_f (new_AGEMA_signal_13081) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L6), .A0_f (new_AGEMA_signal_12488), .A1_t (new_AGEMA_signal_12489), .A1_f (new_AGEMA_signal_12490), .B0_t (SubBytesIns_Inst_Sbox_3_L10), .B0_f (new_AGEMA_signal_12497), .B1_t (new_AGEMA_signal_12498), .B1_f (new_AGEMA_signal_12499), .Z0_t (SubBytesIns_Inst_Sbox_3_L25), .Z0_f (new_AGEMA_signal_13082), .Z1_t (new_AGEMA_signal_13083), .Z1_f (new_AGEMA_signal_13084) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L7), .A0_f (new_AGEMA_signal_12491), .A1_t (new_AGEMA_signal_12492), .A1_f (new_AGEMA_signal_12493), .B0_t (SubBytesIns_Inst_Sbox_3_L9), .B0_f (new_AGEMA_signal_12494), .B1_t (new_AGEMA_signal_12495), .B1_f (new_AGEMA_signal_12496), .Z0_t (SubBytesIns_Inst_Sbox_3_L26), .Z0_f (new_AGEMA_signal_13085), .Z1_t (new_AGEMA_signal_13086), .Z1_f (new_AGEMA_signal_13087) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L8), .A0_f (new_AGEMA_signal_11258), .A1_t (new_AGEMA_signal_11259), .A1_f (new_AGEMA_signal_11260), .B0_t (SubBytesIns_Inst_Sbox_3_L10), .B0_f (new_AGEMA_signal_12497), .B1_t (new_AGEMA_signal_12498), .B1_f (new_AGEMA_signal_12499), .Z0_t (SubBytesIns_Inst_Sbox_3_L27), .Z0_f (new_AGEMA_signal_13088), .Z1_t (new_AGEMA_signal_13089), .Z1_f (new_AGEMA_signal_13090) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L11), .A0_f (new_AGEMA_signal_12500), .A1_t (new_AGEMA_signal_12501), .A1_f (new_AGEMA_signal_12502), .B0_t (SubBytesIns_Inst_Sbox_3_L14), .B0_f (new_AGEMA_signal_11924), .B1_t (new_AGEMA_signal_11925), .B1_f (new_AGEMA_signal_11926), .Z0_t (SubBytesIns_Inst_Sbox_3_L28), .Z0_f (new_AGEMA_signal_13091), .Z1_t (new_AGEMA_signal_13092), .Z1_f (new_AGEMA_signal_13093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L11), .A0_f (new_AGEMA_signal_12500), .A1_t (new_AGEMA_signal_12501), .A1_f (new_AGEMA_signal_12502), .B0_t (SubBytesIns_Inst_Sbox_3_L17), .B0_f (new_AGEMA_signal_11930), .B1_t (new_AGEMA_signal_11931), .B1_f (new_AGEMA_signal_11932), .Z0_t (SubBytesIns_Inst_Sbox_3_L29), .Z0_f (new_AGEMA_signal_13094), .Z1_t (new_AGEMA_signal_13095), .Z1_f (new_AGEMA_signal_13096) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L6), .A0_f (new_AGEMA_signal_12488), .A1_t (new_AGEMA_signal_12489), .A1_f (new_AGEMA_signal_12490), .B0_t (SubBytesIns_Inst_Sbox_3_L24), .B0_f (new_AGEMA_signal_13079), .B1_t (new_AGEMA_signal_13080), .B1_f (new_AGEMA_signal_13081), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .Z0_f (new_AGEMA_signal_13703), .Z1_t (new_AGEMA_signal_13704), .Z1_f (new_AGEMA_signal_13705) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L16), .A0_f (new_AGEMA_signal_13070), .A1_t (new_AGEMA_signal_13071), .A1_f (new_AGEMA_signal_13072), .B0_t (SubBytesIns_Inst_Sbox_3_L26), .B0_f (new_AGEMA_signal_13085), .B1_t (new_AGEMA_signal_13086), .B1_f (new_AGEMA_signal_13087), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .Z0_f (new_AGEMA_signal_13706), .Z1_t (new_AGEMA_signal_13707), .Z1_f (new_AGEMA_signal_13708) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L19), .A0_f (new_AGEMA_signal_12503), .A1_t (new_AGEMA_signal_12504), .A1_f (new_AGEMA_signal_12505), .B0_t (SubBytesIns_Inst_Sbox_3_L28), .B0_f (new_AGEMA_signal_13091), .B1_t (new_AGEMA_signal_13092), .B1_f (new_AGEMA_signal_13093), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .Z0_f (new_AGEMA_signal_13709), .Z1_t (new_AGEMA_signal_13710), .Z1_f (new_AGEMA_signal_13711) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L6), .A0_f (new_AGEMA_signal_12488), .A1_t (new_AGEMA_signal_12489), .A1_f (new_AGEMA_signal_12490), .B0_t (SubBytesIns_Inst_Sbox_3_L21), .B0_f (new_AGEMA_signal_13076), .B1_t (new_AGEMA_signal_13077), .B1_f (new_AGEMA_signal_13078), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .Z0_f (new_AGEMA_signal_13712), .Z1_t (new_AGEMA_signal_13713), .Z1_f (new_AGEMA_signal_13714) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L20), .A0_f (new_AGEMA_signal_13073), .A1_t (new_AGEMA_signal_13074), .A1_f (new_AGEMA_signal_13075), .B0_t (SubBytesIns_Inst_Sbox_3_L22), .B0_f (new_AGEMA_signal_12506), .B1_t (new_AGEMA_signal_12507), .B1_f (new_AGEMA_signal_12508), .Z0_t (MixColumnsInput[27]), .Z0_f (new_AGEMA_signal_13715), .Z1_t (new_AGEMA_signal_13716), .Z1_f (new_AGEMA_signal_13717) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L25), .A0_f (new_AGEMA_signal_13082), .A1_t (new_AGEMA_signal_13083), .A1_f (new_AGEMA_signal_13084), .B0_t (SubBytesIns_Inst_Sbox_3_L29), .B0_f (new_AGEMA_signal_13094), .B1_t (new_AGEMA_signal_13095), .B1_f (new_AGEMA_signal_13096), .Z0_t (MixColumnsInput[26]), .Z0_f (new_AGEMA_signal_13718), .Z1_t (new_AGEMA_signal_13719), .Z1_f (new_AGEMA_signal_13720) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L13), .A0_f (new_AGEMA_signal_13067), .A1_t (new_AGEMA_signal_13068), .A1_f (new_AGEMA_signal_13069), .B0_t (SubBytesIns_Inst_Sbox_3_L27), .B0_f (new_AGEMA_signal_13088), .B1_t (new_AGEMA_signal_13089), .B1_f (new_AGEMA_signal_13090), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .Z0_f (new_AGEMA_signal_13721), .Z1_t (new_AGEMA_signal_13722), .Z1_f (new_AGEMA_signal_13723) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L6), .A0_f (new_AGEMA_signal_12488), .A1_t (new_AGEMA_signal_12489), .A1_f (new_AGEMA_signal_12490), .B0_t (SubBytesIns_Inst_Sbox_3_L23), .B0_f (new_AGEMA_signal_12509), .B1_t (new_AGEMA_signal_12510), .B1_f (new_AGEMA_signal_12511), .Z0_t (MixColumnsInput[24]), .Z0_f (new_AGEMA_signal_13097), .Z1_t (new_AGEMA_signal_13098), .Z1_f (new_AGEMA_signal_13099) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[39]), .A0_f (ciphertext_s0_f[39]), .A1_t (ciphertext_s1_t[39]), .A1_f (ciphertext_s1_f[39]), .B0_t (ciphertext_s0_t[36]), .B0_f (ciphertext_s0_f[36]), .B1_t (ciphertext_s1_t[36]), .B1_f (ciphertext_s1_f[36]), .Z0_t (SubBytesIns_Inst_Sbox_4_T1), .Z0_f (new_AGEMA_signal_6466), .Z1_t (new_AGEMA_signal_6467), .Z1_f (new_AGEMA_signal_6468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[39]), .A0_f (ciphertext_s0_f[39]), .A1_t (ciphertext_s1_t[39]), .A1_f (ciphertext_s1_f[39]), .B0_t (ciphertext_s0_t[34]), .B0_f (ciphertext_s0_f[34]), .B1_t (ciphertext_s1_t[34]), .B1_f (ciphertext_s1_f[34]), .Z0_t (SubBytesIns_Inst_Sbox_4_T2), .Z0_f (new_AGEMA_signal_6469), .Z1_t (new_AGEMA_signal_6470), .Z1_f (new_AGEMA_signal_6471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[39]), .A0_f (ciphertext_s0_f[39]), .A1_t (ciphertext_s1_t[39]), .A1_f (ciphertext_s1_f[39]), .B0_t (ciphertext_s0_t[33]), .B0_f (ciphertext_s0_f[33]), .B1_t (ciphertext_s1_t[33]), .B1_f (ciphertext_s1_f[33]), .Z0_t (SubBytesIns_Inst_Sbox_4_T3), .Z0_f (new_AGEMA_signal_6472), .Z1_t (new_AGEMA_signal_6473), .Z1_f (new_AGEMA_signal_6474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[36]), .A0_f (ciphertext_s0_f[36]), .A1_t (ciphertext_s1_t[36]), .A1_f (ciphertext_s1_f[36]), .B0_t (ciphertext_s0_t[34]), .B0_f (ciphertext_s0_f[34]), .B1_t (ciphertext_s1_t[34]), .B1_f (ciphertext_s1_f[34]), .Z0_t (SubBytesIns_Inst_Sbox_4_T4), .Z0_f (new_AGEMA_signal_6475), .Z1_t (new_AGEMA_signal_6476), .Z1_f (new_AGEMA_signal_6477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[35]), .A0_f (ciphertext_s0_f[35]), .A1_t (ciphertext_s1_t[35]), .A1_f (ciphertext_s1_f[35]), .B0_t (ciphertext_s0_t[33]), .B0_f (ciphertext_s0_f[33]), .B1_t (ciphertext_s1_t[33]), .B1_f (ciphertext_s1_f[33]), .Z0_t (SubBytesIns_Inst_Sbox_4_T5), .Z0_f (new_AGEMA_signal_6478), .Z1_t (new_AGEMA_signal_6479), .Z1_f (new_AGEMA_signal_6480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T1), .A0_f (new_AGEMA_signal_6466), .A1_t (new_AGEMA_signal_6467), .A1_f (new_AGEMA_signal_6468), .B0_t (SubBytesIns_Inst_Sbox_4_T5), .B0_f (new_AGEMA_signal_6478), .B1_t (new_AGEMA_signal_6479), .B1_f (new_AGEMA_signal_6480), .Z0_t (SubBytesIns_Inst_Sbox_4_T6), .Z0_f (new_AGEMA_signal_7024), .Z1_t (new_AGEMA_signal_7025), .Z1_f (new_AGEMA_signal_7026) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[38]), .A0_f (ciphertext_s0_f[38]), .A1_t (ciphertext_s1_t[38]), .A1_f (ciphertext_s1_f[38]), .B0_t (ciphertext_s0_t[37]), .B0_f (ciphertext_s0_f[37]), .B1_t (ciphertext_s1_t[37]), .B1_f (ciphertext_s1_f[37]), .Z0_t (SubBytesIns_Inst_Sbox_4_T7), .Z0_f (new_AGEMA_signal_6481), .Z1_t (new_AGEMA_signal_6482), .Z1_f (new_AGEMA_signal_6483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[32]), .A0_f (ciphertext_s0_f[32]), .A1_t (ciphertext_s1_t[32]), .A1_f (ciphertext_s1_f[32]), .B0_t (SubBytesIns_Inst_Sbox_4_T6), .B0_f (new_AGEMA_signal_7024), .B1_t (new_AGEMA_signal_7025), .B1_f (new_AGEMA_signal_7026), .Z0_t (SubBytesIns_Inst_Sbox_4_T8), .Z0_f (new_AGEMA_signal_7628), .Z1_t (new_AGEMA_signal_7629), .Z1_f (new_AGEMA_signal_7630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[32]), .A0_f (ciphertext_s0_f[32]), .A1_t (ciphertext_s1_t[32]), .A1_f (ciphertext_s1_f[32]), .B0_t (SubBytesIns_Inst_Sbox_4_T7), .B0_f (new_AGEMA_signal_6481), .B1_t (new_AGEMA_signal_6482), .B1_f (new_AGEMA_signal_6483), .Z0_t (SubBytesIns_Inst_Sbox_4_T9), .Z0_f (new_AGEMA_signal_7027), .Z1_t (new_AGEMA_signal_7028), .Z1_f (new_AGEMA_signal_7029) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T6), .A0_f (new_AGEMA_signal_7024), .A1_t (new_AGEMA_signal_7025), .A1_f (new_AGEMA_signal_7026), .B0_t (SubBytesIns_Inst_Sbox_4_T7), .B0_f (new_AGEMA_signal_6481), .B1_t (new_AGEMA_signal_6482), .B1_f (new_AGEMA_signal_6483), .Z0_t (SubBytesIns_Inst_Sbox_4_T10), .Z0_f (new_AGEMA_signal_7631), .Z1_t (new_AGEMA_signal_7632), .Z1_f (new_AGEMA_signal_7633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[38]), .A0_f (ciphertext_s0_f[38]), .A1_t (ciphertext_s1_t[38]), .A1_f (ciphertext_s1_f[38]), .B0_t (ciphertext_s0_t[34]), .B0_f (ciphertext_s0_f[34]), .B1_t (ciphertext_s1_t[34]), .B1_f (ciphertext_s1_f[34]), .Z0_t (SubBytesIns_Inst_Sbox_4_T11), .Z0_f (new_AGEMA_signal_6484), .Z1_t (new_AGEMA_signal_6485), .Z1_f (new_AGEMA_signal_6486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[37]), .A0_f (ciphertext_s0_f[37]), .A1_t (ciphertext_s1_t[37]), .A1_f (ciphertext_s1_f[37]), .B0_t (ciphertext_s0_t[34]), .B0_f (ciphertext_s0_f[34]), .B1_t (ciphertext_s1_t[34]), .B1_f (ciphertext_s1_f[34]), .Z0_t (SubBytesIns_Inst_Sbox_4_T12), .Z0_f (new_AGEMA_signal_6487), .Z1_t (new_AGEMA_signal_6488), .Z1_f (new_AGEMA_signal_6489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T3), .A0_f (new_AGEMA_signal_6472), .A1_t (new_AGEMA_signal_6473), .A1_f (new_AGEMA_signal_6474), .B0_t (SubBytesIns_Inst_Sbox_4_T4), .B0_f (new_AGEMA_signal_6475), .B1_t (new_AGEMA_signal_6476), .B1_f (new_AGEMA_signal_6477), .Z0_t (SubBytesIns_Inst_Sbox_4_T13), .Z0_f (new_AGEMA_signal_7030), .Z1_t (new_AGEMA_signal_7031), .Z1_f (new_AGEMA_signal_7032) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T6), .A0_f (new_AGEMA_signal_7024), .A1_t (new_AGEMA_signal_7025), .A1_f (new_AGEMA_signal_7026), .B0_t (SubBytesIns_Inst_Sbox_4_T11), .B0_f (new_AGEMA_signal_6484), .B1_t (new_AGEMA_signal_6485), .B1_f (new_AGEMA_signal_6486), .Z0_t (SubBytesIns_Inst_Sbox_4_T14), .Z0_f (new_AGEMA_signal_7634), .Z1_t (new_AGEMA_signal_7635), .Z1_f (new_AGEMA_signal_7636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T5), .A0_f (new_AGEMA_signal_6478), .A1_t (new_AGEMA_signal_6479), .A1_f (new_AGEMA_signal_6480), .B0_t (SubBytesIns_Inst_Sbox_4_T11), .B0_f (new_AGEMA_signal_6484), .B1_t (new_AGEMA_signal_6485), .B1_f (new_AGEMA_signal_6486), .Z0_t (SubBytesIns_Inst_Sbox_4_T15), .Z0_f (new_AGEMA_signal_7033), .Z1_t (new_AGEMA_signal_7034), .Z1_f (new_AGEMA_signal_7035) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T5), .A0_f (new_AGEMA_signal_6478), .A1_t (new_AGEMA_signal_6479), .A1_f (new_AGEMA_signal_6480), .B0_t (SubBytesIns_Inst_Sbox_4_T12), .B0_f (new_AGEMA_signal_6487), .B1_t (new_AGEMA_signal_6488), .B1_f (new_AGEMA_signal_6489), .Z0_t (SubBytesIns_Inst_Sbox_4_T16), .Z0_f (new_AGEMA_signal_7036), .Z1_t (new_AGEMA_signal_7037), .Z1_f (new_AGEMA_signal_7038) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T9), .A0_f (new_AGEMA_signal_7027), .A1_t (new_AGEMA_signal_7028), .A1_f (new_AGEMA_signal_7029), .B0_t (SubBytesIns_Inst_Sbox_4_T16), .B0_f (new_AGEMA_signal_7036), .B1_t (new_AGEMA_signal_7037), .B1_f (new_AGEMA_signal_7038), .Z0_t (SubBytesIns_Inst_Sbox_4_T17), .Z0_f (new_AGEMA_signal_7637), .Z1_t (new_AGEMA_signal_7638), .Z1_f (new_AGEMA_signal_7639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[36]), .A0_f (ciphertext_s0_f[36]), .A1_t (ciphertext_s1_t[36]), .A1_f (ciphertext_s1_f[36]), .B0_t (ciphertext_s0_t[32]), .B0_f (ciphertext_s0_f[32]), .B1_t (ciphertext_s1_t[32]), .B1_f (ciphertext_s1_f[32]), .Z0_t (SubBytesIns_Inst_Sbox_4_T18), .Z0_f (new_AGEMA_signal_6490), .Z1_t (new_AGEMA_signal_6491), .Z1_f (new_AGEMA_signal_6492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T7), .A0_f (new_AGEMA_signal_6481), .A1_t (new_AGEMA_signal_6482), .A1_f (new_AGEMA_signal_6483), .B0_t (SubBytesIns_Inst_Sbox_4_T18), .B0_f (new_AGEMA_signal_6490), .B1_t (new_AGEMA_signal_6491), .B1_f (new_AGEMA_signal_6492), .Z0_t (SubBytesIns_Inst_Sbox_4_T19), .Z0_f (new_AGEMA_signal_7039), .Z1_t (new_AGEMA_signal_7040), .Z1_f (new_AGEMA_signal_7041) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T1), .A0_f (new_AGEMA_signal_6466), .A1_t (new_AGEMA_signal_6467), .A1_f (new_AGEMA_signal_6468), .B0_t (SubBytesIns_Inst_Sbox_4_T19), .B0_f (new_AGEMA_signal_7039), .B1_t (new_AGEMA_signal_7040), .B1_f (new_AGEMA_signal_7041), .Z0_t (SubBytesIns_Inst_Sbox_4_T20), .Z0_f (new_AGEMA_signal_7640), .Z1_t (new_AGEMA_signal_7641), .Z1_f (new_AGEMA_signal_7642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[33]), .A0_f (ciphertext_s0_f[33]), .A1_t (ciphertext_s1_t[33]), .A1_f (ciphertext_s1_f[33]), .B0_t (ciphertext_s0_t[32]), .B0_f (ciphertext_s0_f[32]), .B1_t (ciphertext_s1_t[32]), .B1_f (ciphertext_s1_f[32]), .Z0_t (SubBytesIns_Inst_Sbox_4_T21), .Z0_f (new_AGEMA_signal_6493), .Z1_t (new_AGEMA_signal_6494), .Z1_f (new_AGEMA_signal_6495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T7), .A0_f (new_AGEMA_signal_6481), .A1_t (new_AGEMA_signal_6482), .A1_f (new_AGEMA_signal_6483), .B0_t (SubBytesIns_Inst_Sbox_4_T21), .B0_f (new_AGEMA_signal_6493), .B1_t (new_AGEMA_signal_6494), .B1_f (new_AGEMA_signal_6495), .Z0_t (SubBytesIns_Inst_Sbox_4_T22), .Z0_f (new_AGEMA_signal_7042), .Z1_t (new_AGEMA_signal_7043), .Z1_f (new_AGEMA_signal_7044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T2), .A0_f (new_AGEMA_signal_6469), .A1_t (new_AGEMA_signal_6470), .A1_f (new_AGEMA_signal_6471), .B0_t (SubBytesIns_Inst_Sbox_4_T22), .B0_f (new_AGEMA_signal_7042), .B1_t (new_AGEMA_signal_7043), .B1_f (new_AGEMA_signal_7044), .Z0_t (SubBytesIns_Inst_Sbox_4_T23), .Z0_f (new_AGEMA_signal_7643), .Z1_t (new_AGEMA_signal_7644), .Z1_f (new_AGEMA_signal_7645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T2), .A0_f (new_AGEMA_signal_6469), .A1_t (new_AGEMA_signal_6470), .A1_f (new_AGEMA_signal_6471), .B0_t (SubBytesIns_Inst_Sbox_4_T10), .B0_f (new_AGEMA_signal_7631), .B1_t (new_AGEMA_signal_7632), .B1_f (new_AGEMA_signal_7633), .Z0_t (SubBytesIns_Inst_Sbox_4_T24), .Z0_f (new_AGEMA_signal_8312), .Z1_t (new_AGEMA_signal_8313), .Z1_f (new_AGEMA_signal_8314) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T20), .A0_f (new_AGEMA_signal_7640), .A1_t (new_AGEMA_signal_7641), .A1_f (new_AGEMA_signal_7642), .B0_t (SubBytesIns_Inst_Sbox_4_T17), .B0_f (new_AGEMA_signal_7637), .B1_t (new_AGEMA_signal_7638), .B1_f (new_AGEMA_signal_7639), .Z0_t (SubBytesIns_Inst_Sbox_4_T25), .Z0_f (new_AGEMA_signal_8315), .Z1_t (new_AGEMA_signal_8316), .Z1_f (new_AGEMA_signal_8317) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T3), .A0_f (new_AGEMA_signal_6472), .A1_t (new_AGEMA_signal_6473), .A1_f (new_AGEMA_signal_6474), .B0_t (SubBytesIns_Inst_Sbox_4_T16), .B0_f (new_AGEMA_signal_7036), .B1_t (new_AGEMA_signal_7037), .B1_f (new_AGEMA_signal_7038), .Z0_t (SubBytesIns_Inst_Sbox_4_T26), .Z0_f (new_AGEMA_signal_7646), .Z1_t (new_AGEMA_signal_7647), .Z1_f (new_AGEMA_signal_7648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T1), .A0_f (new_AGEMA_signal_6466), .A1_t (new_AGEMA_signal_6467), .A1_f (new_AGEMA_signal_6468), .B0_t (SubBytesIns_Inst_Sbox_4_T12), .B0_f (new_AGEMA_signal_6487), .B1_t (new_AGEMA_signal_6488), .B1_f (new_AGEMA_signal_6489), .Z0_t (SubBytesIns_Inst_Sbox_4_T27), .Z0_f (new_AGEMA_signal_7045), .Z1_t (new_AGEMA_signal_7046), .Z1_f (new_AGEMA_signal_7047) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T13), .A0_f (new_AGEMA_signal_7030), .A1_t (new_AGEMA_signal_7031), .A1_f (new_AGEMA_signal_7032), .B0_t (SubBytesIns_Inst_Sbox_4_T6), .B0_f (new_AGEMA_signal_7024), .B1_t (new_AGEMA_signal_7025), .B1_f (new_AGEMA_signal_7026), .Z0_t (SubBytesIns_Inst_Sbox_4_M1), .Z0_f (new_AGEMA_signal_7649), .Z1_t (new_AGEMA_signal_7650), .Z1_f (new_AGEMA_signal_7651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T23), .A0_f (new_AGEMA_signal_7643), .A1_t (new_AGEMA_signal_7644), .A1_f (new_AGEMA_signal_7645), .B0_t (SubBytesIns_Inst_Sbox_4_T8), .B0_f (new_AGEMA_signal_7628), .B1_t (new_AGEMA_signal_7629), .B1_f (new_AGEMA_signal_7630), .Z0_t (SubBytesIns_Inst_Sbox_4_M2), .Z0_f (new_AGEMA_signal_8318), .Z1_t (new_AGEMA_signal_8319), .Z1_f (new_AGEMA_signal_8320) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T14), .A0_f (new_AGEMA_signal_7634), .A1_t (new_AGEMA_signal_7635), .A1_f (new_AGEMA_signal_7636), .B0_t (SubBytesIns_Inst_Sbox_4_M1), .B0_f (new_AGEMA_signal_7649), .B1_t (new_AGEMA_signal_7650), .B1_f (new_AGEMA_signal_7651), .Z0_t (SubBytesIns_Inst_Sbox_4_M3), .Z0_f (new_AGEMA_signal_8321), .Z1_t (new_AGEMA_signal_8322), .Z1_f (new_AGEMA_signal_8323) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T19), .A0_f (new_AGEMA_signal_7039), .A1_t (new_AGEMA_signal_7040), .A1_f (new_AGEMA_signal_7041), .B0_t (ciphertext_s0_t[32]), .B0_f (ciphertext_s0_f[32]), .B1_t (ciphertext_s1_t[32]), .B1_f (ciphertext_s1_f[32]), .Z0_t (SubBytesIns_Inst_Sbox_4_M4), .Z0_f (new_AGEMA_signal_7652), .Z1_t (new_AGEMA_signal_7653), .Z1_f (new_AGEMA_signal_7654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M4), .A0_f (new_AGEMA_signal_7652), .A1_t (new_AGEMA_signal_7653), .A1_f (new_AGEMA_signal_7654), .B0_t (SubBytesIns_Inst_Sbox_4_M1), .B0_f (new_AGEMA_signal_7649), .B1_t (new_AGEMA_signal_7650), .B1_f (new_AGEMA_signal_7651), .Z0_t (SubBytesIns_Inst_Sbox_4_M5), .Z0_f (new_AGEMA_signal_8324), .Z1_t (new_AGEMA_signal_8325), .Z1_f (new_AGEMA_signal_8326) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T3), .A0_f (new_AGEMA_signal_6472), .A1_t (new_AGEMA_signal_6473), .A1_f (new_AGEMA_signal_6474), .B0_t (SubBytesIns_Inst_Sbox_4_T16), .B0_f (new_AGEMA_signal_7036), .B1_t (new_AGEMA_signal_7037), .B1_f (new_AGEMA_signal_7038), .Z0_t (SubBytesIns_Inst_Sbox_4_M6), .Z0_f (new_AGEMA_signal_7655), .Z1_t (new_AGEMA_signal_7656), .Z1_f (new_AGEMA_signal_7657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T22), .A0_f (new_AGEMA_signal_7042), .A1_t (new_AGEMA_signal_7043), .A1_f (new_AGEMA_signal_7044), .B0_t (SubBytesIns_Inst_Sbox_4_T9), .B0_f (new_AGEMA_signal_7027), .B1_t (new_AGEMA_signal_7028), .B1_f (new_AGEMA_signal_7029), .Z0_t (SubBytesIns_Inst_Sbox_4_M7), .Z0_f (new_AGEMA_signal_7658), .Z1_t (new_AGEMA_signal_7659), .Z1_f (new_AGEMA_signal_7660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T26), .A0_f (new_AGEMA_signal_7646), .A1_t (new_AGEMA_signal_7647), .A1_f (new_AGEMA_signal_7648), .B0_t (SubBytesIns_Inst_Sbox_4_M6), .B0_f (new_AGEMA_signal_7655), .B1_t (new_AGEMA_signal_7656), .B1_f (new_AGEMA_signal_7657), .Z0_t (SubBytesIns_Inst_Sbox_4_M8), .Z0_f (new_AGEMA_signal_8327), .Z1_t (new_AGEMA_signal_8328), .Z1_f (new_AGEMA_signal_8329) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T20), .A0_f (new_AGEMA_signal_7640), .A1_t (new_AGEMA_signal_7641), .A1_f (new_AGEMA_signal_7642), .B0_t (SubBytesIns_Inst_Sbox_4_T17), .B0_f (new_AGEMA_signal_7637), .B1_t (new_AGEMA_signal_7638), .B1_f (new_AGEMA_signal_7639), .Z0_t (SubBytesIns_Inst_Sbox_4_M9), .Z0_f (new_AGEMA_signal_8330), .Z1_t (new_AGEMA_signal_8331), .Z1_f (new_AGEMA_signal_8332) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M9), .A0_f (new_AGEMA_signal_8330), .A1_t (new_AGEMA_signal_8331), .A1_f (new_AGEMA_signal_8332), .B0_t (SubBytesIns_Inst_Sbox_4_M6), .B0_f (new_AGEMA_signal_7655), .B1_t (new_AGEMA_signal_7656), .B1_f (new_AGEMA_signal_7657), .Z0_t (SubBytesIns_Inst_Sbox_4_M10), .Z0_f (new_AGEMA_signal_8756), .Z1_t (new_AGEMA_signal_8757), .Z1_f (new_AGEMA_signal_8758) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T1), .A0_f (new_AGEMA_signal_6466), .A1_t (new_AGEMA_signal_6467), .A1_f (new_AGEMA_signal_6468), .B0_t (SubBytesIns_Inst_Sbox_4_T15), .B0_f (new_AGEMA_signal_7033), .B1_t (new_AGEMA_signal_7034), .B1_f (new_AGEMA_signal_7035), .Z0_t (SubBytesIns_Inst_Sbox_4_M11), .Z0_f (new_AGEMA_signal_7661), .Z1_t (new_AGEMA_signal_7662), .Z1_f (new_AGEMA_signal_7663) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T4), .A0_f (new_AGEMA_signal_6475), .A1_t (new_AGEMA_signal_6476), .A1_f (new_AGEMA_signal_6477), .B0_t (SubBytesIns_Inst_Sbox_4_T27), .B0_f (new_AGEMA_signal_7045), .B1_t (new_AGEMA_signal_7046), .B1_f (new_AGEMA_signal_7047), .Z0_t (SubBytesIns_Inst_Sbox_4_M12), .Z0_f (new_AGEMA_signal_7664), .Z1_t (new_AGEMA_signal_7665), .Z1_f (new_AGEMA_signal_7666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M12), .A0_f (new_AGEMA_signal_7664), .A1_t (new_AGEMA_signal_7665), .A1_f (new_AGEMA_signal_7666), .B0_t (SubBytesIns_Inst_Sbox_4_M11), .B0_f (new_AGEMA_signal_7661), .B1_t (new_AGEMA_signal_7662), .B1_f (new_AGEMA_signal_7663), .Z0_t (SubBytesIns_Inst_Sbox_4_M13), .Z0_f (new_AGEMA_signal_8333), .Z1_t (new_AGEMA_signal_8334), .Z1_f (new_AGEMA_signal_8335) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T2), .A0_f (new_AGEMA_signal_6469), .A1_t (new_AGEMA_signal_6470), .A1_f (new_AGEMA_signal_6471), .B0_t (SubBytesIns_Inst_Sbox_4_T10), .B0_f (new_AGEMA_signal_7631), .B1_t (new_AGEMA_signal_7632), .B1_f (new_AGEMA_signal_7633), .Z0_t (SubBytesIns_Inst_Sbox_4_M14), .Z0_f (new_AGEMA_signal_8336), .Z1_t (new_AGEMA_signal_8337), .Z1_f (new_AGEMA_signal_8338) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M14), .A0_f (new_AGEMA_signal_8336), .A1_t (new_AGEMA_signal_8337), .A1_f (new_AGEMA_signal_8338), .B0_t (SubBytesIns_Inst_Sbox_4_M11), .B0_f (new_AGEMA_signal_7661), .B1_t (new_AGEMA_signal_7662), .B1_f (new_AGEMA_signal_7663), .Z0_t (SubBytesIns_Inst_Sbox_4_M15), .Z0_f (new_AGEMA_signal_8759), .Z1_t (new_AGEMA_signal_8760), .Z1_f (new_AGEMA_signal_8761) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M3), .A0_f (new_AGEMA_signal_8321), .A1_t (new_AGEMA_signal_8322), .A1_f (new_AGEMA_signal_8323), .B0_t (SubBytesIns_Inst_Sbox_4_M2), .B0_f (new_AGEMA_signal_8318), .B1_t (new_AGEMA_signal_8319), .B1_f (new_AGEMA_signal_8320), .Z0_t (SubBytesIns_Inst_Sbox_4_M16), .Z0_f (new_AGEMA_signal_8762), .Z1_t (new_AGEMA_signal_8763), .Z1_f (new_AGEMA_signal_8764) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M5), .A0_f (new_AGEMA_signal_8324), .A1_t (new_AGEMA_signal_8325), .A1_f (new_AGEMA_signal_8326), .B0_t (SubBytesIns_Inst_Sbox_4_T24), .B0_f (new_AGEMA_signal_8312), .B1_t (new_AGEMA_signal_8313), .B1_f (new_AGEMA_signal_8314), .Z0_t (SubBytesIns_Inst_Sbox_4_M17), .Z0_f (new_AGEMA_signal_8765), .Z1_t (new_AGEMA_signal_8766), .Z1_f (new_AGEMA_signal_8767) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M8), .A0_f (new_AGEMA_signal_8327), .A1_t (new_AGEMA_signal_8328), .A1_f (new_AGEMA_signal_8329), .B0_t (SubBytesIns_Inst_Sbox_4_M7), .B0_f (new_AGEMA_signal_7658), .B1_t (new_AGEMA_signal_7659), .B1_f (new_AGEMA_signal_7660), .Z0_t (SubBytesIns_Inst_Sbox_4_M18), .Z0_f (new_AGEMA_signal_8768), .Z1_t (new_AGEMA_signal_8769), .Z1_f (new_AGEMA_signal_8770) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M10), .A0_f (new_AGEMA_signal_8756), .A1_t (new_AGEMA_signal_8757), .A1_f (new_AGEMA_signal_8758), .B0_t (SubBytesIns_Inst_Sbox_4_M15), .B0_f (new_AGEMA_signal_8759), .B1_t (new_AGEMA_signal_8760), .B1_f (new_AGEMA_signal_8761), .Z0_t (SubBytesIns_Inst_Sbox_4_M19), .Z0_f (new_AGEMA_signal_9032), .Z1_t (new_AGEMA_signal_9033), .Z1_f (new_AGEMA_signal_9034) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M16), .A0_f (new_AGEMA_signal_8762), .A1_t (new_AGEMA_signal_8763), .A1_f (new_AGEMA_signal_8764), .B0_t (SubBytesIns_Inst_Sbox_4_M13), .B0_f (new_AGEMA_signal_8333), .B1_t (new_AGEMA_signal_8334), .B1_f (new_AGEMA_signal_8335), .Z0_t (SubBytesIns_Inst_Sbox_4_M20), .Z0_f (new_AGEMA_signal_9035), .Z1_t (new_AGEMA_signal_9036), .Z1_f (new_AGEMA_signal_9037) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M17), .A0_f (new_AGEMA_signal_8765), .A1_t (new_AGEMA_signal_8766), .A1_f (new_AGEMA_signal_8767), .B0_t (SubBytesIns_Inst_Sbox_4_M15), .B0_f (new_AGEMA_signal_8759), .B1_t (new_AGEMA_signal_8760), .B1_f (new_AGEMA_signal_8761), .Z0_t (SubBytesIns_Inst_Sbox_4_M21), .Z0_f (new_AGEMA_signal_9038), .Z1_t (new_AGEMA_signal_9039), .Z1_f (new_AGEMA_signal_9040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M18), .A0_f (new_AGEMA_signal_8768), .A1_t (new_AGEMA_signal_8769), .A1_f (new_AGEMA_signal_8770), .B0_t (SubBytesIns_Inst_Sbox_4_M13), .B0_f (new_AGEMA_signal_8333), .B1_t (new_AGEMA_signal_8334), .B1_f (new_AGEMA_signal_8335), .Z0_t (SubBytesIns_Inst_Sbox_4_M22), .Z0_f (new_AGEMA_signal_9041), .Z1_t (new_AGEMA_signal_9042), .Z1_f (new_AGEMA_signal_9043) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M19), .A0_f (new_AGEMA_signal_9032), .A1_t (new_AGEMA_signal_9033), .A1_f (new_AGEMA_signal_9034), .B0_t (SubBytesIns_Inst_Sbox_4_T25), .B0_f (new_AGEMA_signal_8315), .B1_t (new_AGEMA_signal_8316), .B1_f (new_AGEMA_signal_8317), .Z0_t (SubBytesIns_Inst_Sbox_4_M23), .Z0_f (new_AGEMA_signal_9272), .Z1_t (new_AGEMA_signal_9273), .Z1_f (new_AGEMA_signal_9274) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M22), .A0_f (new_AGEMA_signal_9041), .A1_t (new_AGEMA_signal_9042), .A1_f (new_AGEMA_signal_9043), .B0_t (SubBytesIns_Inst_Sbox_4_M23), .B0_f (new_AGEMA_signal_9272), .B1_t (new_AGEMA_signal_9273), .B1_f (new_AGEMA_signal_9274), .Z0_t (SubBytesIns_Inst_Sbox_4_M24), .Z0_f (new_AGEMA_signal_9536), .Z1_t (new_AGEMA_signal_9537), .Z1_f (new_AGEMA_signal_9538) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M22), .A0_f (new_AGEMA_signal_9041), .A1_t (new_AGEMA_signal_9042), .A1_f (new_AGEMA_signal_9043), .B0_t (SubBytesIns_Inst_Sbox_4_M20), .B0_f (new_AGEMA_signal_9035), .B1_t (new_AGEMA_signal_9036), .B1_f (new_AGEMA_signal_9037), .Z0_t (SubBytesIns_Inst_Sbox_4_M25), .Z0_f (new_AGEMA_signal_9275), .Z1_t (new_AGEMA_signal_9276), .Z1_f (new_AGEMA_signal_9277) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M21), .A0_f (new_AGEMA_signal_9038), .A1_t (new_AGEMA_signal_9039), .A1_f (new_AGEMA_signal_9040), .B0_t (SubBytesIns_Inst_Sbox_4_M25), .B0_f (new_AGEMA_signal_9275), .B1_t (new_AGEMA_signal_9276), .B1_f (new_AGEMA_signal_9277), .Z0_t (SubBytesIns_Inst_Sbox_4_M26), .Z0_f (new_AGEMA_signal_9539), .Z1_t (new_AGEMA_signal_9540), .Z1_f (new_AGEMA_signal_9541) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M20), .A0_f (new_AGEMA_signal_9035), .A1_t (new_AGEMA_signal_9036), .A1_f (new_AGEMA_signal_9037), .B0_t (SubBytesIns_Inst_Sbox_4_M21), .B0_f (new_AGEMA_signal_9038), .B1_t (new_AGEMA_signal_9039), .B1_f (new_AGEMA_signal_9040), .Z0_t (SubBytesIns_Inst_Sbox_4_M27), .Z0_f (new_AGEMA_signal_9278), .Z1_t (new_AGEMA_signal_9279), .Z1_f (new_AGEMA_signal_9280) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M23), .A0_f (new_AGEMA_signal_9272), .A1_t (new_AGEMA_signal_9273), .A1_f (new_AGEMA_signal_9274), .B0_t (SubBytesIns_Inst_Sbox_4_M25), .B0_f (new_AGEMA_signal_9275), .B1_t (new_AGEMA_signal_9276), .B1_f (new_AGEMA_signal_9277), .Z0_t (SubBytesIns_Inst_Sbox_4_M28), .Z0_f (new_AGEMA_signal_9542), .Z1_t (new_AGEMA_signal_9543), .Z1_f (new_AGEMA_signal_9544) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M28), .A0_f (new_AGEMA_signal_9542), .A1_t (new_AGEMA_signal_9543), .A1_f (new_AGEMA_signal_9544), .B0_t (SubBytesIns_Inst_Sbox_4_M27), .B0_f (new_AGEMA_signal_9278), .B1_t (new_AGEMA_signal_9279), .B1_f (new_AGEMA_signal_9280), .Z0_t (SubBytesIns_Inst_Sbox_4_M29), .Z0_f (new_AGEMA_signal_9836), .Z1_t (new_AGEMA_signal_9837), .Z1_f (new_AGEMA_signal_9838) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M26), .A0_f (new_AGEMA_signal_9539), .A1_t (new_AGEMA_signal_9540), .A1_f (new_AGEMA_signal_9541), .B0_t (SubBytesIns_Inst_Sbox_4_M24), .B0_f (new_AGEMA_signal_9536), .B1_t (new_AGEMA_signal_9537), .B1_f (new_AGEMA_signal_9538), .Z0_t (SubBytesIns_Inst_Sbox_4_M30), .Z0_f (new_AGEMA_signal_9839), .Z1_t (new_AGEMA_signal_9840), .Z1_f (new_AGEMA_signal_9841) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M20), .A0_f (new_AGEMA_signal_9035), .A1_t (new_AGEMA_signal_9036), .A1_f (new_AGEMA_signal_9037), .B0_t (SubBytesIns_Inst_Sbox_4_M23), .B0_f (new_AGEMA_signal_9272), .B1_t (new_AGEMA_signal_9273), .B1_f (new_AGEMA_signal_9274), .Z0_t (SubBytesIns_Inst_Sbox_4_M31), .Z0_f (new_AGEMA_signal_9545), .Z1_t (new_AGEMA_signal_9546), .Z1_f (new_AGEMA_signal_9547) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M27), .A0_f (new_AGEMA_signal_9278), .A1_t (new_AGEMA_signal_9279), .A1_f (new_AGEMA_signal_9280), .B0_t (SubBytesIns_Inst_Sbox_4_M31), .B0_f (new_AGEMA_signal_9545), .B1_t (new_AGEMA_signal_9546), .B1_f (new_AGEMA_signal_9547), .Z0_t (SubBytesIns_Inst_Sbox_4_M32), .Z0_f (new_AGEMA_signal_9842), .Z1_t (new_AGEMA_signal_9843), .Z1_f (new_AGEMA_signal_9844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M27), .A0_f (new_AGEMA_signal_9278), .A1_t (new_AGEMA_signal_9279), .A1_f (new_AGEMA_signal_9280), .B0_t (SubBytesIns_Inst_Sbox_4_M25), .B0_f (new_AGEMA_signal_9275), .B1_t (new_AGEMA_signal_9276), .B1_f (new_AGEMA_signal_9277), .Z0_t (SubBytesIns_Inst_Sbox_4_M33), .Z0_f (new_AGEMA_signal_9548), .Z1_t (new_AGEMA_signal_9549), .Z1_f (new_AGEMA_signal_9550) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M21), .A0_f (new_AGEMA_signal_9038), .A1_t (new_AGEMA_signal_9039), .A1_f (new_AGEMA_signal_9040), .B0_t (SubBytesIns_Inst_Sbox_4_M22), .B0_f (new_AGEMA_signal_9041), .B1_t (new_AGEMA_signal_9042), .B1_f (new_AGEMA_signal_9043), .Z0_t (SubBytesIns_Inst_Sbox_4_M34), .Z0_f (new_AGEMA_signal_9281), .Z1_t (new_AGEMA_signal_9282), .Z1_f (new_AGEMA_signal_9283) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M24), .A0_f (new_AGEMA_signal_9536), .A1_t (new_AGEMA_signal_9537), .A1_f (new_AGEMA_signal_9538), .B0_t (SubBytesIns_Inst_Sbox_4_M34), .B0_f (new_AGEMA_signal_9281), .B1_t (new_AGEMA_signal_9282), .B1_f (new_AGEMA_signal_9283), .Z0_t (SubBytesIns_Inst_Sbox_4_M35), .Z0_f (new_AGEMA_signal_9845), .Z1_t (new_AGEMA_signal_9846), .Z1_f (new_AGEMA_signal_9847) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M24), .A0_f (new_AGEMA_signal_9536), .A1_t (new_AGEMA_signal_9537), .A1_f (new_AGEMA_signal_9538), .B0_t (SubBytesIns_Inst_Sbox_4_M25), .B0_f (new_AGEMA_signal_9275), .B1_t (new_AGEMA_signal_9276), .B1_f (new_AGEMA_signal_9277), .Z0_t (SubBytesIns_Inst_Sbox_4_M36), .Z0_f (new_AGEMA_signal_9848), .Z1_t (new_AGEMA_signal_9849), .Z1_f (new_AGEMA_signal_9850) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M21), .A0_f (new_AGEMA_signal_9038), .A1_t (new_AGEMA_signal_9039), .A1_f (new_AGEMA_signal_9040), .B0_t (SubBytesIns_Inst_Sbox_4_M29), .B0_f (new_AGEMA_signal_9836), .B1_t (new_AGEMA_signal_9837), .B1_f (new_AGEMA_signal_9838), .Z0_t (SubBytesIns_Inst_Sbox_4_M37), .Z0_f (new_AGEMA_signal_10112), .Z1_t (new_AGEMA_signal_10113), .Z1_f (new_AGEMA_signal_10114) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M32), .A0_f (new_AGEMA_signal_9842), .A1_t (new_AGEMA_signal_9843), .A1_f (new_AGEMA_signal_9844), .B0_t (SubBytesIns_Inst_Sbox_4_M33), .B0_f (new_AGEMA_signal_9548), .B1_t (new_AGEMA_signal_9549), .B1_f (new_AGEMA_signal_9550), .Z0_t (SubBytesIns_Inst_Sbox_4_M38), .Z0_f (new_AGEMA_signal_10115), .Z1_t (new_AGEMA_signal_10116), .Z1_f (new_AGEMA_signal_10117) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M23), .A0_f (new_AGEMA_signal_9272), .A1_t (new_AGEMA_signal_9273), .A1_f (new_AGEMA_signal_9274), .B0_t (SubBytesIns_Inst_Sbox_4_M30), .B0_f (new_AGEMA_signal_9839), .B1_t (new_AGEMA_signal_9840), .B1_f (new_AGEMA_signal_9841), .Z0_t (SubBytesIns_Inst_Sbox_4_M39), .Z0_f (new_AGEMA_signal_10118), .Z1_t (new_AGEMA_signal_10119), .Z1_f (new_AGEMA_signal_10120) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M35), .A0_f (new_AGEMA_signal_9845), .A1_t (new_AGEMA_signal_9846), .A1_f (new_AGEMA_signal_9847), .B0_t (SubBytesIns_Inst_Sbox_4_M36), .B0_f (new_AGEMA_signal_9848), .B1_t (new_AGEMA_signal_9849), .B1_f (new_AGEMA_signal_9850), .Z0_t (SubBytesIns_Inst_Sbox_4_M40), .Z0_f (new_AGEMA_signal_10121), .Z1_t (new_AGEMA_signal_10122), .Z1_f (new_AGEMA_signal_10123) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M38), .A0_f (new_AGEMA_signal_10115), .A1_t (new_AGEMA_signal_10116), .A1_f (new_AGEMA_signal_10117), .B0_t (SubBytesIns_Inst_Sbox_4_M40), .B0_f (new_AGEMA_signal_10121), .B1_t (new_AGEMA_signal_10122), .B1_f (new_AGEMA_signal_10123), .Z0_t (SubBytesIns_Inst_Sbox_4_M41), .Z0_f (new_AGEMA_signal_10544), .Z1_t (new_AGEMA_signal_10545), .Z1_f (new_AGEMA_signal_10546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M37), .A0_f (new_AGEMA_signal_10112), .A1_t (new_AGEMA_signal_10113), .A1_f (new_AGEMA_signal_10114), .B0_t (SubBytesIns_Inst_Sbox_4_M39), .B0_f (new_AGEMA_signal_10118), .B1_t (new_AGEMA_signal_10119), .B1_f (new_AGEMA_signal_10120), .Z0_t (SubBytesIns_Inst_Sbox_4_M42), .Z0_f (new_AGEMA_signal_10547), .Z1_t (new_AGEMA_signal_10548), .Z1_f (new_AGEMA_signal_10549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M37), .A0_f (new_AGEMA_signal_10112), .A1_t (new_AGEMA_signal_10113), .A1_f (new_AGEMA_signal_10114), .B0_t (SubBytesIns_Inst_Sbox_4_M38), .B0_f (new_AGEMA_signal_10115), .B1_t (new_AGEMA_signal_10116), .B1_f (new_AGEMA_signal_10117), .Z0_t (SubBytesIns_Inst_Sbox_4_M43), .Z0_f (new_AGEMA_signal_10550), .Z1_t (new_AGEMA_signal_10551), .Z1_f (new_AGEMA_signal_10552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M39), .A0_f (new_AGEMA_signal_10118), .A1_t (new_AGEMA_signal_10119), .A1_f (new_AGEMA_signal_10120), .B0_t (SubBytesIns_Inst_Sbox_4_M40), .B0_f (new_AGEMA_signal_10121), .B1_t (new_AGEMA_signal_10122), .B1_f (new_AGEMA_signal_10123), .Z0_t (SubBytesIns_Inst_Sbox_4_M44), .Z0_f (new_AGEMA_signal_10553), .Z1_t (new_AGEMA_signal_10554), .Z1_f (new_AGEMA_signal_10555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M42), .A0_f (new_AGEMA_signal_10547), .A1_t (new_AGEMA_signal_10548), .A1_f (new_AGEMA_signal_10549), .B0_t (SubBytesIns_Inst_Sbox_4_M41), .B0_f (new_AGEMA_signal_10544), .B1_t (new_AGEMA_signal_10545), .B1_f (new_AGEMA_signal_10546), .Z0_t (SubBytesIns_Inst_Sbox_4_M45), .Z0_f (new_AGEMA_signal_11264), .Z1_t (new_AGEMA_signal_11265), .Z1_f (new_AGEMA_signal_11266) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M44), .A0_f (new_AGEMA_signal_10553), .A1_t (new_AGEMA_signal_10554), .A1_f (new_AGEMA_signal_10555), .B0_t (SubBytesIns_Inst_Sbox_4_T6), .B0_f (new_AGEMA_signal_7024), .B1_t (new_AGEMA_signal_7025), .B1_f (new_AGEMA_signal_7026), .Z0_t (SubBytesIns_Inst_Sbox_4_M46), .Z0_f (new_AGEMA_signal_11267), .Z1_t (new_AGEMA_signal_11268), .Z1_f (new_AGEMA_signal_11269) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M40), .A0_f (new_AGEMA_signal_10121), .A1_t (new_AGEMA_signal_10122), .A1_f (new_AGEMA_signal_10123), .B0_t (SubBytesIns_Inst_Sbox_4_T8), .B0_f (new_AGEMA_signal_7628), .B1_t (new_AGEMA_signal_7629), .B1_f (new_AGEMA_signal_7630), .Z0_t (SubBytesIns_Inst_Sbox_4_M47), .Z0_f (new_AGEMA_signal_10556), .Z1_t (new_AGEMA_signal_10557), .Z1_f (new_AGEMA_signal_10558) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M39), .A0_f (new_AGEMA_signal_10118), .A1_t (new_AGEMA_signal_10119), .A1_f (new_AGEMA_signal_10120), .B0_t (ciphertext_s0_t[32]), .B0_f (ciphertext_s0_f[32]), .B1_t (ciphertext_s1_t[32]), .B1_f (ciphertext_s1_f[32]), .Z0_t (SubBytesIns_Inst_Sbox_4_M48), .Z0_f (new_AGEMA_signal_10559), .Z1_t (new_AGEMA_signal_10560), .Z1_f (new_AGEMA_signal_10561) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M43), .A0_f (new_AGEMA_signal_10550), .A1_t (new_AGEMA_signal_10551), .A1_f (new_AGEMA_signal_10552), .B0_t (SubBytesIns_Inst_Sbox_4_T16), .B0_f (new_AGEMA_signal_7036), .B1_t (new_AGEMA_signal_7037), .B1_f (new_AGEMA_signal_7038), .Z0_t (SubBytesIns_Inst_Sbox_4_M49), .Z0_f (new_AGEMA_signal_11270), .Z1_t (new_AGEMA_signal_11271), .Z1_f (new_AGEMA_signal_11272) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M38), .A0_f (new_AGEMA_signal_10115), .A1_t (new_AGEMA_signal_10116), .A1_f (new_AGEMA_signal_10117), .B0_t (SubBytesIns_Inst_Sbox_4_T9), .B0_f (new_AGEMA_signal_7027), .B1_t (new_AGEMA_signal_7028), .B1_f (new_AGEMA_signal_7029), .Z0_t (SubBytesIns_Inst_Sbox_4_M50), .Z0_f (new_AGEMA_signal_10562), .Z1_t (new_AGEMA_signal_10563), .Z1_f (new_AGEMA_signal_10564) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M37), .A0_f (new_AGEMA_signal_10112), .A1_t (new_AGEMA_signal_10113), .A1_f (new_AGEMA_signal_10114), .B0_t (SubBytesIns_Inst_Sbox_4_T17), .B0_f (new_AGEMA_signal_7637), .B1_t (new_AGEMA_signal_7638), .B1_f (new_AGEMA_signal_7639), .Z0_t (SubBytesIns_Inst_Sbox_4_M51), .Z0_f (new_AGEMA_signal_10565), .Z1_t (new_AGEMA_signal_10566), .Z1_f (new_AGEMA_signal_10567) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M42), .A0_f (new_AGEMA_signal_10547), .A1_t (new_AGEMA_signal_10548), .A1_f (new_AGEMA_signal_10549), .B0_t (SubBytesIns_Inst_Sbox_4_T15), .B0_f (new_AGEMA_signal_7033), .B1_t (new_AGEMA_signal_7034), .B1_f (new_AGEMA_signal_7035), .Z0_t (SubBytesIns_Inst_Sbox_4_M52), .Z0_f (new_AGEMA_signal_11273), .Z1_t (new_AGEMA_signal_11274), .Z1_f (new_AGEMA_signal_11275) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M45), .A0_f (new_AGEMA_signal_11264), .A1_t (new_AGEMA_signal_11265), .A1_f (new_AGEMA_signal_11266), .B0_t (SubBytesIns_Inst_Sbox_4_T27), .B0_f (new_AGEMA_signal_7045), .B1_t (new_AGEMA_signal_7046), .B1_f (new_AGEMA_signal_7047), .Z0_t (SubBytesIns_Inst_Sbox_4_M53), .Z0_f (new_AGEMA_signal_11936), .Z1_t (new_AGEMA_signal_11937), .Z1_f (new_AGEMA_signal_11938) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M41), .A0_f (new_AGEMA_signal_10544), .A1_t (new_AGEMA_signal_10545), .A1_f (new_AGEMA_signal_10546), .B0_t (SubBytesIns_Inst_Sbox_4_T10), .B0_f (new_AGEMA_signal_7631), .B1_t (new_AGEMA_signal_7632), .B1_f (new_AGEMA_signal_7633), .Z0_t (SubBytesIns_Inst_Sbox_4_M54), .Z0_f (new_AGEMA_signal_11276), .Z1_t (new_AGEMA_signal_11277), .Z1_f (new_AGEMA_signal_11278) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M44), .A0_f (new_AGEMA_signal_10553), .A1_t (new_AGEMA_signal_10554), .A1_f (new_AGEMA_signal_10555), .B0_t (SubBytesIns_Inst_Sbox_4_T13), .B0_f (new_AGEMA_signal_7030), .B1_t (new_AGEMA_signal_7031), .B1_f (new_AGEMA_signal_7032), .Z0_t (SubBytesIns_Inst_Sbox_4_M55), .Z0_f (new_AGEMA_signal_11279), .Z1_t (new_AGEMA_signal_11280), .Z1_f (new_AGEMA_signal_11281) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M40), .A0_f (new_AGEMA_signal_10121), .A1_t (new_AGEMA_signal_10122), .A1_f (new_AGEMA_signal_10123), .B0_t (SubBytesIns_Inst_Sbox_4_T23), .B0_f (new_AGEMA_signal_7643), .B1_t (new_AGEMA_signal_7644), .B1_f (new_AGEMA_signal_7645), .Z0_t (SubBytesIns_Inst_Sbox_4_M56), .Z0_f (new_AGEMA_signal_10568), .Z1_t (new_AGEMA_signal_10569), .Z1_f (new_AGEMA_signal_10570) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M39), .A0_f (new_AGEMA_signal_10118), .A1_t (new_AGEMA_signal_10119), .A1_f (new_AGEMA_signal_10120), .B0_t (SubBytesIns_Inst_Sbox_4_T19), .B0_f (new_AGEMA_signal_7039), .B1_t (new_AGEMA_signal_7040), .B1_f (new_AGEMA_signal_7041), .Z0_t (SubBytesIns_Inst_Sbox_4_M57), .Z0_f (new_AGEMA_signal_10571), .Z1_t (new_AGEMA_signal_10572), .Z1_f (new_AGEMA_signal_10573) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M43), .A0_f (new_AGEMA_signal_10550), .A1_t (new_AGEMA_signal_10551), .A1_f (new_AGEMA_signal_10552), .B0_t (SubBytesIns_Inst_Sbox_4_T3), .B0_f (new_AGEMA_signal_6472), .B1_t (new_AGEMA_signal_6473), .B1_f (new_AGEMA_signal_6474), .Z0_t (SubBytesIns_Inst_Sbox_4_M58), .Z0_f (new_AGEMA_signal_11282), .Z1_t (new_AGEMA_signal_11283), .Z1_f (new_AGEMA_signal_11284) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M38), .A0_f (new_AGEMA_signal_10115), .A1_t (new_AGEMA_signal_10116), .A1_f (new_AGEMA_signal_10117), .B0_t (SubBytesIns_Inst_Sbox_4_T22), .B0_f (new_AGEMA_signal_7042), .B1_t (new_AGEMA_signal_7043), .B1_f (new_AGEMA_signal_7044), .Z0_t (SubBytesIns_Inst_Sbox_4_M59), .Z0_f (new_AGEMA_signal_10574), .Z1_t (new_AGEMA_signal_10575), .Z1_f (new_AGEMA_signal_10576) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M37), .A0_f (new_AGEMA_signal_10112), .A1_t (new_AGEMA_signal_10113), .A1_f (new_AGEMA_signal_10114), .B0_t (SubBytesIns_Inst_Sbox_4_T20), .B0_f (new_AGEMA_signal_7640), .B1_t (new_AGEMA_signal_7641), .B1_f (new_AGEMA_signal_7642), .Z0_t (SubBytesIns_Inst_Sbox_4_M60), .Z0_f (new_AGEMA_signal_10577), .Z1_t (new_AGEMA_signal_10578), .Z1_f (new_AGEMA_signal_10579) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M42), .A0_f (new_AGEMA_signal_10547), .A1_t (new_AGEMA_signal_10548), .A1_f (new_AGEMA_signal_10549), .B0_t (SubBytesIns_Inst_Sbox_4_T1), .B0_f (new_AGEMA_signal_6466), .B1_t (new_AGEMA_signal_6467), .B1_f (new_AGEMA_signal_6468), .Z0_t (SubBytesIns_Inst_Sbox_4_M61), .Z0_f (new_AGEMA_signal_11285), .Z1_t (new_AGEMA_signal_11286), .Z1_f (new_AGEMA_signal_11287) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M45), .A0_f (new_AGEMA_signal_11264), .A1_t (new_AGEMA_signal_11265), .A1_f (new_AGEMA_signal_11266), .B0_t (SubBytesIns_Inst_Sbox_4_T4), .B0_f (new_AGEMA_signal_6475), .B1_t (new_AGEMA_signal_6476), .B1_f (new_AGEMA_signal_6477), .Z0_t (SubBytesIns_Inst_Sbox_4_M62), .Z0_f (new_AGEMA_signal_11939), .Z1_t (new_AGEMA_signal_11940), .Z1_f (new_AGEMA_signal_11941) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M41), .A0_f (new_AGEMA_signal_10544), .A1_t (new_AGEMA_signal_10545), .A1_f (new_AGEMA_signal_10546), .B0_t (SubBytesIns_Inst_Sbox_4_T2), .B0_f (new_AGEMA_signal_6469), .B1_t (new_AGEMA_signal_6470), .B1_f (new_AGEMA_signal_6471), .Z0_t (SubBytesIns_Inst_Sbox_4_M63), .Z0_f (new_AGEMA_signal_11288), .Z1_t (new_AGEMA_signal_11289), .Z1_f (new_AGEMA_signal_11290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M61), .A0_f (new_AGEMA_signal_11285), .A1_t (new_AGEMA_signal_11286), .A1_f (new_AGEMA_signal_11287), .B0_t (SubBytesIns_Inst_Sbox_4_M62), .B0_f (new_AGEMA_signal_11939), .B1_t (new_AGEMA_signal_11940), .B1_f (new_AGEMA_signal_11941), .Z0_t (SubBytesIns_Inst_Sbox_4_L0), .Z0_f (new_AGEMA_signal_12512), .Z1_t (new_AGEMA_signal_12513), .Z1_f (new_AGEMA_signal_12514) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M50), .A0_f (new_AGEMA_signal_10562), .A1_t (new_AGEMA_signal_10563), .A1_f (new_AGEMA_signal_10564), .B0_t (SubBytesIns_Inst_Sbox_4_M56), .B0_f (new_AGEMA_signal_10568), .B1_t (new_AGEMA_signal_10569), .B1_f (new_AGEMA_signal_10570), .Z0_t (SubBytesIns_Inst_Sbox_4_L1), .Z0_f (new_AGEMA_signal_11291), .Z1_t (new_AGEMA_signal_11292), .Z1_f (new_AGEMA_signal_11293) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M46), .A0_f (new_AGEMA_signal_11267), .A1_t (new_AGEMA_signal_11268), .A1_f (new_AGEMA_signal_11269), .B0_t (SubBytesIns_Inst_Sbox_4_M48), .B0_f (new_AGEMA_signal_10559), .B1_t (new_AGEMA_signal_10560), .B1_f (new_AGEMA_signal_10561), .Z0_t (SubBytesIns_Inst_Sbox_4_L2), .Z0_f (new_AGEMA_signal_11942), .Z1_t (new_AGEMA_signal_11943), .Z1_f (new_AGEMA_signal_11944) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M47), .A0_f (new_AGEMA_signal_10556), .A1_t (new_AGEMA_signal_10557), .A1_f (new_AGEMA_signal_10558), .B0_t (SubBytesIns_Inst_Sbox_4_M55), .B0_f (new_AGEMA_signal_11279), .B1_t (new_AGEMA_signal_11280), .B1_f (new_AGEMA_signal_11281), .Z0_t (SubBytesIns_Inst_Sbox_4_L3), .Z0_f (new_AGEMA_signal_11945), .Z1_t (new_AGEMA_signal_11946), .Z1_f (new_AGEMA_signal_11947) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M54), .A0_f (new_AGEMA_signal_11276), .A1_t (new_AGEMA_signal_11277), .A1_f (new_AGEMA_signal_11278), .B0_t (SubBytesIns_Inst_Sbox_4_M58), .B0_f (new_AGEMA_signal_11282), .B1_t (new_AGEMA_signal_11283), .B1_f (new_AGEMA_signal_11284), .Z0_t (SubBytesIns_Inst_Sbox_4_L4), .Z0_f (new_AGEMA_signal_11948), .Z1_t (new_AGEMA_signal_11949), .Z1_f (new_AGEMA_signal_11950) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M49), .A0_f (new_AGEMA_signal_11270), .A1_t (new_AGEMA_signal_11271), .A1_f (new_AGEMA_signal_11272), .B0_t (SubBytesIns_Inst_Sbox_4_M61), .B0_f (new_AGEMA_signal_11285), .B1_t (new_AGEMA_signal_11286), .B1_f (new_AGEMA_signal_11287), .Z0_t (SubBytesIns_Inst_Sbox_4_L5), .Z0_f (new_AGEMA_signal_11951), .Z1_t (new_AGEMA_signal_11952), .Z1_f (new_AGEMA_signal_11953) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M62), .A0_f (new_AGEMA_signal_11939), .A1_t (new_AGEMA_signal_11940), .A1_f (new_AGEMA_signal_11941), .B0_t (SubBytesIns_Inst_Sbox_4_L5), .B0_f (new_AGEMA_signal_11951), .B1_t (new_AGEMA_signal_11952), .B1_f (new_AGEMA_signal_11953), .Z0_t (SubBytesIns_Inst_Sbox_4_L6), .Z0_f (new_AGEMA_signal_12515), .Z1_t (new_AGEMA_signal_12516), .Z1_f (new_AGEMA_signal_12517) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M46), .A0_f (new_AGEMA_signal_11267), .A1_t (new_AGEMA_signal_11268), .A1_f (new_AGEMA_signal_11269), .B0_t (SubBytesIns_Inst_Sbox_4_L3), .B0_f (new_AGEMA_signal_11945), .B1_t (new_AGEMA_signal_11946), .B1_f (new_AGEMA_signal_11947), .Z0_t (SubBytesIns_Inst_Sbox_4_L7), .Z0_f (new_AGEMA_signal_12518), .Z1_t (new_AGEMA_signal_12519), .Z1_f (new_AGEMA_signal_12520) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M51), .A0_f (new_AGEMA_signal_10565), .A1_t (new_AGEMA_signal_10566), .A1_f (new_AGEMA_signal_10567), .B0_t (SubBytesIns_Inst_Sbox_4_M59), .B0_f (new_AGEMA_signal_10574), .B1_t (new_AGEMA_signal_10575), .B1_f (new_AGEMA_signal_10576), .Z0_t (SubBytesIns_Inst_Sbox_4_L8), .Z0_f (new_AGEMA_signal_11294), .Z1_t (new_AGEMA_signal_11295), .Z1_f (new_AGEMA_signal_11296) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M52), .A0_f (new_AGEMA_signal_11273), .A1_t (new_AGEMA_signal_11274), .A1_f (new_AGEMA_signal_11275), .B0_t (SubBytesIns_Inst_Sbox_4_M53), .B0_f (new_AGEMA_signal_11936), .B1_t (new_AGEMA_signal_11937), .B1_f (new_AGEMA_signal_11938), .Z0_t (SubBytesIns_Inst_Sbox_4_L9), .Z0_f (new_AGEMA_signal_12521), .Z1_t (new_AGEMA_signal_12522), .Z1_f (new_AGEMA_signal_12523) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M53), .A0_f (new_AGEMA_signal_11936), .A1_t (new_AGEMA_signal_11937), .A1_f (new_AGEMA_signal_11938), .B0_t (SubBytesIns_Inst_Sbox_4_L4), .B0_f (new_AGEMA_signal_11948), .B1_t (new_AGEMA_signal_11949), .B1_f (new_AGEMA_signal_11950), .Z0_t (SubBytesIns_Inst_Sbox_4_L10), .Z0_f (new_AGEMA_signal_12524), .Z1_t (new_AGEMA_signal_12525), .Z1_f (new_AGEMA_signal_12526) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M60), .A0_f (new_AGEMA_signal_10577), .A1_t (new_AGEMA_signal_10578), .A1_f (new_AGEMA_signal_10579), .B0_t (SubBytesIns_Inst_Sbox_4_L2), .B0_f (new_AGEMA_signal_11942), .B1_t (new_AGEMA_signal_11943), .B1_f (new_AGEMA_signal_11944), .Z0_t (SubBytesIns_Inst_Sbox_4_L11), .Z0_f (new_AGEMA_signal_12527), .Z1_t (new_AGEMA_signal_12528), .Z1_f (new_AGEMA_signal_12529) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M48), .A0_f (new_AGEMA_signal_10559), .A1_t (new_AGEMA_signal_10560), .A1_f (new_AGEMA_signal_10561), .B0_t (SubBytesIns_Inst_Sbox_4_M51), .B0_f (new_AGEMA_signal_10565), .B1_t (new_AGEMA_signal_10566), .B1_f (new_AGEMA_signal_10567), .Z0_t (SubBytesIns_Inst_Sbox_4_L12), .Z0_f (new_AGEMA_signal_11297), .Z1_t (new_AGEMA_signal_11298), .Z1_f (new_AGEMA_signal_11299) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M50), .A0_f (new_AGEMA_signal_10562), .A1_t (new_AGEMA_signal_10563), .A1_f (new_AGEMA_signal_10564), .B0_t (SubBytesIns_Inst_Sbox_4_L0), .B0_f (new_AGEMA_signal_12512), .B1_t (new_AGEMA_signal_12513), .B1_f (new_AGEMA_signal_12514), .Z0_t (SubBytesIns_Inst_Sbox_4_L13), .Z0_f (new_AGEMA_signal_13100), .Z1_t (new_AGEMA_signal_13101), .Z1_f (new_AGEMA_signal_13102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M52), .A0_f (new_AGEMA_signal_11273), .A1_t (new_AGEMA_signal_11274), .A1_f (new_AGEMA_signal_11275), .B0_t (SubBytesIns_Inst_Sbox_4_M61), .B0_f (new_AGEMA_signal_11285), .B1_t (new_AGEMA_signal_11286), .B1_f (new_AGEMA_signal_11287), .Z0_t (SubBytesIns_Inst_Sbox_4_L14), .Z0_f (new_AGEMA_signal_11954), .Z1_t (new_AGEMA_signal_11955), .Z1_f (new_AGEMA_signal_11956) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M55), .A0_f (new_AGEMA_signal_11279), .A1_t (new_AGEMA_signal_11280), .A1_f (new_AGEMA_signal_11281), .B0_t (SubBytesIns_Inst_Sbox_4_L1), .B0_f (new_AGEMA_signal_11291), .B1_t (new_AGEMA_signal_11292), .B1_f (new_AGEMA_signal_11293), .Z0_t (SubBytesIns_Inst_Sbox_4_L15), .Z0_f (new_AGEMA_signal_11957), .Z1_t (new_AGEMA_signal_11958), .Z1_f (new_AGEMA_signal_11959) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M56), .A0_f (new_AGEMA_signal_10568), .A1_t (new_AGEMA_signal_10569), .A1_f (new_AGEMA_signal_10570), .B0_t (SubBytesIns_Inst_Sbox_4_L0), .B0_f (new_AGEMA_signal_12512), .B1_t (new_AGEMA_signal_12513), .B1_f (new_AGEMA_signal_12514), .Z0_t (SubBytesIns_Inst_Sbox_4_L16), .Z0_f (new_AGEMA_signal_13103), .Z1_t (new_AGEMA_signal_13104), .Z1_f (new_AGEMA_signal_13105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M57), .A0_f (new_AGEMA_signal_10571), .A1_t (new_AGEMA_signal_10572), .A1_f (new_AGEMA_signal_10573), .B0_t (SubBytesIns_Inst_Sbox_4_L1), .B0_f (new_AGEMA_signal_11291), .B1_t (new_AGEMA_signal_11292), .B1_f (new_AGEMA_signal_11293), .Z0_t (SubBytesIns_Inst_Sbox_4_L17), .Z0_f (new_AGEMA_signal_11960), .Z1_t (new_AGEMA_signal_11961), .Z1_f (new_AGEMA_signal_11962) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M58), .A0_f (new_AGEMA_signal_11282), .A1_t (new_AGEMA_signal_11283), .A1_f (new_AGEMA_signal_11284), .B0_t (SubBytesIns_Inst_Sbox_4_L8), .B0_f (new_AGEMA_signal_11294), .B1_t (new_AGEMA_signal_11295), .B1_f (new_AGEMA_signal_11296), .Z0_t (SubBytesIns_Inst_Sbox_4_L18), .Z0_f (new_AGEMA_signal_11963), .Z1_t (new_AGEMA_signal_11964), .Z1_f (new_AGEMA_signal_11965) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M63), .A0_f (new_AGEMA_signal_11288), .A1_t (new_AGEMA_signal_11289), .A1_f (new_AGEMA_signal_11290), .B0_t (SubBytesIns_Inst_Sbox_4_L4), .B0_f (new_AGEMA_signal_11948), .B1_t (new_AGEMA_signal_11949), .B1_f (new_AGEMA_signal_11950), .Z0_t (SubBytesIns_Inst_Sbox_4_L19), .Z0_f (new_AGEMA_signal_12530), .Z1_t (new_AGEMA_signal_12531), .Z1_f (new_AGEMA_signal_12532) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L0), .A0_f (new_AGEMA_signal_12512), .A1_t (new_AGEMA_signal_12513), .A1_f (new_AGEMA_signal_12514), .B0_t (SubBytesIns_Inst_Sbox_4_L1), .B0_f (new_AGEMA_signal_11291), .B1_t (new_AGEMA_signal_11292), .B1_f (new_AGEMA_signal_11293), .Z0_t (SubBytesIns_Inst_Sbox_4_L20), .Z0_f (new_AGEMA_signal_13106), .Z1_t (new_AGEMA_signal_13107), .Z1_f (new_AGEMA_signal_13108) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L1), .A0_f (new_AGEMA_signal_11291), .A1_t (new_AGEMA_signal_11292), .A1_f (new_AGEMA_signal_11293), .B0_t (SubBytesIns_Inst_Sbox_4_L7), .B0_f (new_AGEMA_signal_12518), .B1_t (new_AGEMA_signal_12519), .B1_f (new_AGEMA_signal_12520), .Z0_t (SubBytesIns_Inst_Sbox_4_L21), .Z0_f (new_AGEMA_signal_13109), .Z1_t (new_AGEMA_signal_13110), .Z1_f (new_AGEMA_signal_13111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L3), .A0_f (new_AGEMA_signal_11945), .A1_t (new_AGEMA_signal_11946), .A1_f (new_AGEMA_signal_11947), .B0_t (SubBytesIns_Inst_Sbox_4_L12), .B0_f (new_AGEMA_signal_11297), .B1_t (new_AGEMA_signal_11298), .B1_f (new_AGEMA_signal_11299), .Z0_t (SubBytesIns_Inst_Sbox_4_L22), .Z0_f (new_AGEMA_signal_12533), .Z1_t (new_AGEMA_signal_12534), .Z1_f (new_AGEMA_signal_12535) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L18), .A0_f (new_AGEMA_signal_11963), .A1_t (new_AGEMA_signal_11964), .A1_f (new_AGEMA_signal_11965), .B0_t (SubBytesIns_Inst_Sbox_4_L2), .B0_f (new_AGEMA_signal_11942), .B1_t (new_AGEMA_signal_11943), .B1_f (new_AGEMA_signal_11944), .Z0_t (SubBytesIns_Inst_Sbox_4_L23), .Z0_f (new_AGEMA_signal_12536), .Z1_t (new_AGEMA_signal_12537), .Z1_f (new_AGEMA_signal_12538) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L15), .A0_f (new_AGEMA_signal_11957), .A1_t (new_AGEMA_signal_11958), .A1_f (new_AGEMA_signal_11959), .B0_t (SubBytesIns_Inst_Sbox_4_L9), .B0_f (new_AGEMA_signal_12521), .B1_t (new_AGEMA_signal_12522), .B1_f (new_AGEMA_signal_12523), .Z0_t (SubBytesIns_Inst_Sbox_4_L24), .Z0_f (new_AGEMA_signal_13112), .Z1_t (new_AGEMA_signal_13113), .Z1_f (new_AGEMA_signal_13114) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L6), .A0_f (new_AGEMA_signal_12515), .A1_t (new_AGEMA_signal_12516), .A1_f (new_AGEMA_signal_12517), .B0_t (SubBytesIns_Inst_Sbox_4_L10), .B0_f (new_AGEMA_signal_12524), .B1_t (new_AGEMA_signal_12525), .B1_f (new_AGEMA_signal_12526), .Z0_t (SubBytesIns_Inst_Sbox_4_L25), .Z0_f (new_AGEMA_signal_13115), .Z1_t (new_AGEMA_signal_13116), .Z1_f (new_AGEMA_signal_13117) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L7), .A0_f (new_AGEMA_signal_12518), .A1_t (new_AGEMA_signal_12519), .A1_f (new_AGEMA_signal_12520), .B0_t (SubBytesIns_Inst_Sbox_4_L9), .B0_f (new_AGEMA_signal_12521), .B1_t (new_AGEMA_signal_12522), .B1_f (new_AGEMA_signal_12523), .Z0_t (SubBytesIns_Inst_Sbox_4_L26), .Z0_f (new_AGEMA_signal_13118), .Z1_t (new_AGEMA_signal_13119), .Z1_f (new_AGEMA_signal_13120) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L8), .A0_f (new_AGEMA_signal_11294), .A1_t (new_AGEMA_signal_11295), .A1_f (new_AGEMA_signal_11296), .B0_t (SubBytesIns_Inst_Sbox_4_L10), .B0_f (new_AGEMA_signal_12524), .B1_t (new_AGEMA_signal_12525), .B1_f (new_AGEMA_signal_12526), .Z0_t (SubBytesIns_Inst_Sbox_4_L27), .Z0_f (new_AGEMA_signal_13121), .Z1_t (new_AGEMA_signal_13122), .Z1_f (new_AGEMA_signal_13123) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L11), .A0_f (new_AGEMA_signal_12527), .A1_t (new_AGEMA_signal_12528), .A1_f (new_AGEMA_signal_12529), .B0_t (SubBytesIns_Inst_Sbox_4_L14), .B0_f (new_AGEMA_signal_11954), .B1_t (new_AGEMA_signal_11955), .B1_f (new_AGEMA_signal_11956), .Z0_t (SubBytesIns_Inst_Sbox_4_L28), .Z0_f (new_AGEMA_signal_13124), .Z1_t (new_AGEMA_signal_13125), .Z1_f (new_AGEMA_signal_13126) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L11), .A0_f (new_AGEMA_signal_12527), .A1_t (new_AGEMA_signal_12528), .A1_f (new_AGEMA_signal_12529), .B0_t (SubBytesIns_Inst_Sbox_4_L17), .B0_f (new_AGEMA_signal_11960), .B1_t (new_AGEMA_signal_11961), .B1_f (new_AGEMA_signal_11962), .Z0_t (SubBytesIns_Inst_Sbox_4_L29), .Z0_f (new_AGEMA_signal_13127), .Z1_t (new_AGEMA_signal_13128), .Z1_f (new_AGEMA_signal_13129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L6), .A0_f (new_AGEMA_signal_12515), .A1_t (new_AGEMA_signal_12516), .A1_f (new_AGEMA_signal_12517), .B0_t (SubBytesIns_Inst_Sbox_4_L24), .B0_f (new_AGEMA_signal_13112), .B1_t (new_AGEMA_signal_13113), .B1_f (new_AGEMA_signal_13114), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .Z0_f (new_AGEMA_signal_13724), .Z1_t (new_AGEMA_signal_13725), .Z1_f (new_AGEMA_signal_13726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L16), .A0_f (new_AGEMA_signal_13103), .A1_t (new_AGEMA_signal_13104), .A1_f (new_AGEMA_signal_13105), .B0_t (SubBytesIns_Inst_Sbox_4_L26), .B0_f (new_AGEMA_signal_13118), .B1_t (new_AGEMA_signal_13119), .B1_f (new_AGEMA_signal_13120), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .Z0_f (new_AGEMA_signal_13727), .Z1_t (new_AGEMA_signal_13728), .Z1_f (new_AGEMA_signal_13729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L19), .A0_f (new_AGEMA_signal_12530), .A1_t (new_AGEMA_signal_12531), .A1_f (new_AGEMA_signal_12532), .B0_t (SubBytesIns_Inst_Sbox_4_L28), .B0_f (new_AGEMA_signal_13124), .B1_t (new_AGEMA_signal_13125), .B1_f (new_AGEMA_signal_13126), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .Z0_f (new_AGEMA_signal_13730), .Z1_t (new_AGEMA_signal_13731), .Z1_f (new_AGEMA_signal_13732) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L6), .A0_f (new_AGEMA_signal_12515), .A1_t (new_AGEMA_signal_12516), .A1_f (new_AGEMA_signal_12517), .B0_t (SubBytesIns_Inst_Sbox_4_L21), .B0_f (new_AGEMA_signal_13109), .B1_t (new_AGEMA_signal_13110), .B1_f (new_AGEMA_signal_13111), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .Z0_f (new_AGEMA_signal_13733), .Z1_t (new_AGEMA_signal_13734), .Z1_f (new_AGEMA_signal_13735) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L20), .A0_f (new_AGEMA_signal_13106), .A1_t (new_AGEMA_signal_13107), .A1_f (new_AGEMA_signal_13108), .B0_t (SubBytesIns_Inst_Sbox_4_L22), .B0_f (new_AGEMA_signal_12533), .B1_t (new_AGEMA_signal_12534), .B1_f (new_AGEMA_signal_12535), .Z0_t (MixColumnsInput[3]), .Z0_f (new_AGEMA_signal_13736), .Z1_t (new_AGEMA_signal_13737), .Z1_f (new_AGEMA_signal_13738) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L25), .A0_f (new_AGEMA_signal_13115), .A1_t (new_AGEMA_signal_13116), .A1_f (new_AGEMA_signal_13117), .B0_t (SubBytesIns_Inst_Sbox_4_L29), .B0_f (new_AGEMA_signal_13127), .B1_t (new_AGEMA_signal_13128), .B1_f (new_AGEMA_signal_13129), .Z0_t (MixColumnsInput[2]), .Z0_f (new_AGEMA_signal_13739), .Z1_t (new_AGEMA_signal_13740), .Z1_f (new_AGEMA_signal_13741) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L13), .A0_f (new_AGEMA_signal_13100), .A1_t (new_AGEMA_signal_13101), .A1_f (new_AGEMA_signal_13102), .B0_t (SubBytesIns_Inst_Sbox_4_L27), .B0_f (new_AGEMA_signal_13121), .B1_t (new_AGEMA_signal_13122), .B1_f (new_AGEMA_signal_13123), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .Z0_f (new_AGEMA_signal_13742), .Z1_t (new_AGEMA_signal_13743), .Z1_f (new_AGEMA_signal_13744) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L6), .A0_f (new_AGEMA_signal_12515), .A1_t (new_AGEMA_signal_12516), .A1_f (new_AGEMA_signal_12517), .B0_t (SubBytesIns_Inst_Sbox_4_L23), .B0_f (new_AGEMA_signal_12536), .B1_t (new_AGEMA_signal_12537), .B1_f (new_AGEMA_signal_12538), .Z0_t (MixColumnsInput[0]), .Z0_f (new_AGEMA_signal_13130), .Z1_t (new_AGEMA_signal_13131), .Z1_f (new_AGEMA_signal_13132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[47]), .A0_f (ciphertext_s0_f[47]), .A1_t (ciphertext_s1_t[47]), .A1_f (ciphertext_s1_f[47]), .B0_t (ciphertext_s0_t[44]), .B0_f (ciphertext_s0_f[44]), .B1_t (ciphertext_s1_t[44]), .B1_f (ciphertext_s1_f[44]), .Z0_t (SubBytesIns_Inst_Sbox_5_T1), .Z0_f (new_AGEMA_signal_6496), .Z1_t (new_AGEMA_signal_6497), .Z1_f (new_AGEMA_signal_6498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[47]), .A0_f (ciphertext_s0_f[47]), .A1_t (ciphertext_s1_t[47]), .A1_f (ciphertext_s1_f[47]), .B0_t (ciphertext_s0_t[42]), .B0_f (ciphertext_s0_f[42]), .B1_t (ciphertext_s1_t[42]), .B1_f (ciphertext_s1_f[42]), .Z0_t (SubBytesIns_Inst_Sbox_5_T2), .Z0_f (new_AGEMA_signal_6499), .Z1_t (new_AGEMA_signal_6500), .Z1_f (new_AGEMA_signal_6501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[47]), .A0_f (ciphertext_s0_f[47]), .A1_t (ciphertext_s1_t[47]), .A1_f (ciphertext_s1_f[47]), .B0_t (ciphertext_s0_t[41]), .B0_f (ciphertext_s0_f[41]), .B1_t (ciphertext_s1_t[41]), .B1_f (ciphertext_s1_f[41]), .Z0_t (SubBytesIns_Inst_Sbox_5_T3), .Z0_f (new_AGEMA_signal_6502), .Z1_t (new_AGEMA_signal_6503), .Z1_f (new_AGEMA_signal_6504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[44]), .A0_f (ciphertext_s0_f[44]), .A1_t (ciphertext_s1_t[44]), .A1_f (ciphertext_s1_f[44]), .B0_t (ciphertext_s0_t[42]), .B0_f (ciphertext_s0_f[42]), .B1_t (ciphertext_s1_t[42]), .B1_f (ciphertext_s1_f[42]), .Z0_t (SubBytesIns_Inst_Sbox_5_T4), .Z0_f (new_AGEMA_signal_6505), .Z1_t (new_AGEMA_signal_6506), .Z1_f (new_AGEMA_signal_6507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[43]), .A0_f (ciphertext_s0_f[43]), .A1_t (ciphertext_s1_t[43]), .A1_f (ciphertext_s1_f[43]), .B0_t (ciphertext_s0_t[41]), .B0_f (ciphertext_s0_f[41]), .B1_t (ciphertext_s1_t[41]), .B1_f (ciphertext_s1_f[41]), .Z0_t (SubBytesIns_Inst_Sbox_5_T5), .Z0_f (new_AGEMA_signal_6508), .Z1_t (new_AGEMA_signal_6509), .Z1_f (new_AGEMA_signal_6510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T1), .A0_f (new_AGEMA_signal_6496), .A1_t (new_AGEMA_signal_6497), .A1_f (new_AGEMA_signal_6498), .B0_t (SubBytesIns_Inst_Sbox_5_T5), .B0_f (new_AGEMA_signal_6508), .B1_t (new_AGEMA_signal_6509), .B1_f (new_AGEMA_signal_6510), .Z0_t (SubBytesIns_Inst_Sbox_5_T6), .Z0_f (new_AGEMA_signal_7048), .Z1_t (new_AGEMA_signal_7049), .Z1_f (new_AGEMA_signal_7050) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[46]), .A0_f (ciphertext_s0_f[46]), .A1_t (ciphertext_s1_t[46]), .A1_f (ciphertext_s1_f[46]), .B0_t (ciphertext_s0_t[45]), .B0_f (ciphertext_s0_f[45]), .B1_t (ciphertext_s1_t[45]), .B1_f (ciphertext_s1_f[45]), .Z0_t (SubBytesIns_Inst_Sbox_5_T7), .Z0_f (new_AGEMA_signal_6511), .Z1_t (new_AGEMA_signal_6512), .Z1_f (new_AGEMA_signal_6513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[40]), .A0_f (ciphertext_s0_f[40]), .A1_t (ciphertext_s1_t[40]), .A1_f (ciphertext_s1_f[40]), .B0_t (SubBytesIns_Inst_Sbox_5_T6), .B0_f (new_AGEMA_signal_7048), .B1_t (new_AGEMA_signal_7049), .B1_f (new_AGEMA_signal_7050), .Z0_t (SubBytesIns_Inst_Sbox_5_T8), .Z0_f (new_AGEMA_signal_7667), .Z1_t (new_AGEMA_signal_7668), .Z1_f (new_AGEMA_signal_7669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[40]), .A0_f (ciphertext_s0_f[40]), .A1_t (ciphertext_s1_t[40]), .A1_f (ciphertext_s1_f[40]), .B0_t (SubBytesIns_Inst_Sbox_5_T7), .B0_f (new_AGEMA_signal_6511), .B1_t (new_AGEMA_signal_6512), .B1_f (new_AGEMA_signal_6513), .Z0_t (SubBytesIns_Inst_Sbox_5_T9), .Z0_f (new_AGEMA_signal_7051), .Z1_t (new_AGEMA_signal_7052), .Z1_f (new_AGEMA_signal_7053) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T6), .A0_f (new_AGEMA_signal_7048), .A1_t (new_AGEMA_signal_7049), .A1_f (new_AGEMA_signal_7050), .B0_t (SubBytesIns_Inst_Sbox_5_T7), .B0_f (new_AGEMA_signal_6511), .B1_t (new_AGEMA_signal_6512), .B1_f (new_AGEMA_signal_6513), .Z0_t (SubBytesIns_Inst_Sbox_5_T10), .Z0_f (new_AGEMA_signal_7670), .Z1_t (new_AGEMA_signal_7671), .Z1_f (new_AGEMA_signal_7672) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[46]), .A0_f (ciphertext_s0_f[46]), .A1_t (ciphertext_s1_t[46]), .A1_f (ciphertext_s1_f[46]), .B0_t (ciphertext_s0_t[42]), .B0_f (ciphertext_s0_f[42]), .B1_t (ciphertext_s1_t[42]), .B1_f (ciphertext_s1_f[42]), .Z0_t (SubBytesIns_Inst_Sbox_5_T11), .Z0_f (new_AGEMA_signal_6514), .Z1_t (new_AGEMA_signal_6515), .Z1_f (new_AGEMA_signal_6516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[45]), .A0_f (ciphertext_s0_f[45]), .A1_t (ciphertext_s1_t[45]), .A1_f (ciphertext_s1_f[45]), .B0_t (ciphertext_s0_t[42]), .B0_f (ciphertext_s0_f[42]), .B1_t (ciphertext_s1_t[42]), .B1_f (ciphertext_s1_f[42]), .Z0_t (SubBytesIns_Inst_Sbox_5_T12), .Z0_f (new_AGEMA_signal_6517), .Z1_t (new_AGEMA_signal_6518), .Z1_f (new_AGEMA_signal_6519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T3), .A0_f (new_AGEMA_signal_6502), .A1_t (new_AGEMA_signal_6503), .A1_f (new_AGEMA_signal_6504), .B0_t (SubBytesIns_Inst_Sbox_5_T4), .B0_f (new_AGEMA_signal_6505), .B1_t (new_AGEMA_signal_6506), .B1_f (new_AGEMA_signal_6507), .Z0_t (SubBytesIns_Inst_Sbox_5_T13), .Z0_f (new_AGEMA_signal_7054), .Z1_t (new_AGEMA_signal_7055), .Z1_f (new_AGEMA_signal_7056) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T6), .A0_f (new_AGEMA_signal_7048), .A1_t (new_AGEMA_signal_7049), .A1_f (new_AGEMA_signal_7050), .B0_t (SubBytesIns_Inst_Sbox_5_T11), .B0_f (new_AGEMA_signal_6514), .B1_t (new_AGEMA_signal_6515), .B1_f (new_AGEMA_signal_6516), .Z0_t (SubBytesIns_Inst_Sbox_5_T14), .Z0_f (new_AGEMA_signal_7673), .Z1_t (new_AGEMA_signal_7674), .Z1_f (new_AGEMA_signal_7675) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T5), .A0_f (new_AGEMA_signal_6508), .A1_t (new_AGEMA_signal_6509), .A1_f (new_AGEMA_signal_6510), .B0_t (SubBytesIns_Inst_Sbox_5_T11), .B0_f (new_AGEMA_signal_6514), .B1_t (new_AGEMA_signal_6515), .B1_f (new_AGEMA_signal_6516), .Z0_t (SubBytesIns_Inst_Sbox_5_T15), .Z0_f (new_AGEMA_signal_7057), .Z1_t (new_AGEMA_signal_7058), .Z1_f (new_AGEMA_signal_7059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T5), .A0_f (new_AGEMA_signal_6508), .A1_t (new_AGEMA_signal_6509), .A1_f (new_AGEMA_signal_6510), .B0_t (SubBytesIns_Inst_Sbox_5_T12), .B0_f (new_AGEMA_signal_6517), .B1_t (new_AGEMA_signal_6518), .B1_f (new_AGEMA_signal_6519), .Z0_t (SubBytesIns_Inst_Sbox_5_T16), .Z0_f (new_AGEMA_signal_7060), .Z1_t (new_AGEMA_signal_7061), .Z1_f (new_AGEMA_signal_7062) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T9), .A0_f (new_AGEMA_signal_7051), .A1_t (new_AGEMA_signal_7052), .A1_f (new_AGEMA_signal_7053), .B0_t (SubBytesIns_Inst_Sbox_5_T16), .B0_f (new_AGEMA_signal_7060), .B1_t (new_AGEMA_signal_7061), .B1_f (new_AGEMA_signal_7062), .Z0_t (SubBytesIns_Inst_Sbox_5_T17), .Z0_f (new_AGEMA_signal_7676), .Z1_t (new_AGEMA_signal_7677), .Z1_f (new_AGEMA_signal_7678) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[44]), .A0_f (ciphertext_s0_f[44]), .A1_t (ciphertext_s1_t[44]), .A1_f (ciphertext_s1_f[44]), .B0_t (ciphertext_s0_t[40]), .B0_f (ciphertext_s0_f[40]), .B1_t (ciphertext_s1_t[40]), .B1_f (ciphertext_s1_f[40]), .Z0_t (SubBytesIns_Inst_Sbox_5_T18), .Z0_f (new_AGEMA_signal_6520), .Z1_t (new_AGEMA_signal_6521), .Z1_f (new_AGEMA_signal_6522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T7), .A0_f (new_AGEMA_signal_6511), .A1_t (new_AGEMA_signal_6512), .A1_f (new_AGEMA_signal_6513), .B0_t (SubBytesIns_Inst_Sbox_5_T18), .B0_f (new_AGEMA_signal_6520), .B1_t (new_AGEMA_signal_6521), .B1_f (new_AGEMA_signal_6522), .Z0_t (SubBytesIns_Inst_Sbox_5_T19), .Z0_f (new_AGEMA_signal_7063), .Z1_t (new_AGEMA_signal_7064), .Z1_f (new_AGEMA_signal_7065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T1), .A0_f (new_AGEMA_signal_6496), .A1_t (new_AGEMA_signal_6497), .A1_f (new_AGEMA_signal_6498), .B0_t (SubBytesIns_Inst_Sbox_5_T19), .B0_f (new_AGEMA_signal_7063), .B1_t (new_AGEMA_signal_7064), .B1_f (new_AGEMA_signal_7065), .Z0_t (SubBytesIns_Inst_Sbox_5_T20), .Z0_f (new_AGEMA_signal_7679), .Z1_t (new_AGEMA_signal_7680), .Z1_f (new_AGEMA_signal_7681) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[41]), .A0_f (ciphertext_s0_f[41]), .A1_t (ciphertext_s1_t[41]), .A1_f (ciphertext_s1_f[41]), .B0_t (ciphertext_s0_t[40]), .B0_f (ciphertext_s0_f[40]), .B1_t (ciphertext_s1_t[40]), .B1_f (ciphertext_s1_f[40]), .Z0_t (SubBytesIns_Inst_Sbox_5_T21), .Z0_f (new_AGEMA_signal_6523), .Z1_t (new_AGEMA_signal_6524), .Z1_f (new_AGEMA_signal_6525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T7), .A0_f (new_AGEMA_signal_6511), .A1_t (new_AGEMA_signal_6512), .A1_f (new_AGEMA_signal_6513), .B0_t (SubBytesIns_Inst_Sbox_5_T21), .B0_f (new_AGEMA_signal_6523), .B1_t (new_AGEMA_signal_6524), .B1_f (new_AGEMA_signal_6525), .Z0_t (SubBytesIns_Inst_Sbox_5_T22), .Z0_f (new_AGEMA_signal_7066), .Z1_t (new_AGEMA_signal_7067), .Z1_f (new_AGEMA_signal_7068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T2), .A0_f (new_AGEMA_signal_6499), .A1_t (new_AGEMA_signal_6500), .A1_f (new_AGEMA_signal_6501), .B0_t (SubBytesIns_Inst_Sbox_5_T22), .B0_f (new_AGEMA_signal_7066), .B1_t (new_AGEMA_signal_7067), .B1_f (new_AGEMA_signal_7068), .Z0_t (SubBytesIns_Inst_Sbox_5_T23), .Z0_f (new_AGEMA_signal_7682), .Z1_t (new_AGEMA_signal_7683), .Z1_f (new_AGEMA_signal_7684) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T2), .A0_f (new_AGEMA_signal_6499), .A1_t (new_AGEMA_signal_6500), .A1_f (new_AGEMA_signal_6501), .B0_t (SubBytesIns_Inst_Sbox_5_T10), .B0_f (new_AGEMA_signal_7670), .B1_t (new_AGEMA_signal_7671), .B1_f (new_AGEMA_signal_7672), .Z0_t (SubBytesIns_Inst_Sbox_5_T24), .Z0_f (new_AGEMA_signal_8339), .Z1_t (new_AGEMA_signal_8340), .Z1_f (new_AGEMA_signal_8341) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T20), .A0_f (new_AGEMA_signal_7679), .A1_t (new_AGEMA_signal_7680), .A1_f (new_AGEMA_signal_7681), .B0_t (SubBytesIns_Inst_Sbox_5_T17), .B0_f (new_AGEMA_signal_7676), .B1_t (new_AGEMA_signal_7677), .B1_f (new_AGEMA_signal_7678), .Z0_t (SubBytesIns_Inst_Sbox_5_T25), .Z0_f (new_AGEMA_signal_8342), .Z1_t (new_AGEMA_signal_8343), .Z1_f (new_AGEMA_signal_8344) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T3), .A0_f (new_AGEMA_signal_6502), .A1_t (new_AGEMA_signal_6503), .A1_f (new_AGEMA_signal_6504), .B0_t (SubBytesIns_Inst_Sbox_5_T16), .B0_f (new_AGEMA_signal_7060), .B1_t (new_AGEMA_signal_7061), .B1_f (new_AGEMA_signal_7062), .Z0_t (SubBytesIns_Inst_Sbox_5_T26), .Z0_f (new_AGEMA_signal_7685), .Z1_t (new_AGEMA_signal_7686), .Z1_f (new_AGEMA_signal_7687) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T1), .A0_f (new_AGEMA_signal_6496), .A1_t (new_AGEMA_signal_6497), .A1_f (new_AGEMA_signal_6498), .B0_t (SubBytesIns_Inst_Sbox_5_T12), .B0_f (new_AGEMA_signal_6517), .B1_t (new_AGEMA_signal_6518), .B1_f (new_AGEMA_signal_6519), .Z0_t (SubBytesIns_Inst_Sbox_5_T27), .Z0_f (new_AGEMA_signal_7069), .Z1_t (new_AGEMA_signal_7070), .Z1_f (new_AGEMA_signal_7071) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T13), .A0_f (new_AGEMA_signal_7054), .A1_t (new_AGEMA_signal_7055), .A1_f (new_AGEMA_signal_7056), .B0_t (SubBytesIns_Inst_Sbox_5_T6), .B0_f (new_AGEMA_signal_7048), .B1_t (new_AGEMA_signal_7049), .B1_f (new_AGEMA_signal_7050), .Z0_t (SubBytesIns_Inst_Sbox_5_M1), .Z0_f (new_AGEMA_signal_7688), .Z1_t (new_AGEMA_signal_7689), .Z1_f (new_AGEMA_signal_7690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T23), .A0_f (new_AGEMA_signal_7682), .A1_t (new_AGEMA_signal_7683), .A1_f (new_AGEMA_signal_7684), .B0_t (SubBytesIns_Inst_Sbox_5_T8), .B0_f (new_AGEMA_signal_7667), .B1_t (new_AGEMA_signal_7668), .B1_f (new_AGEMA_signal_7669), .Z0_t (SubBytesIns_Inst_Sbox_5_M2), .Z0_f (new_AGEMA_signal_8345), .Z1_t (new_AGEMA_signal_8346), .Z1_f (new_AGEMA_signal_8347) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T14), .A0_f (new_AGEMA_signal_7673), .A1_t (new_AGEMA_signal_7674), .A1_f (new_AGEMA_signal_7675), .B0_t (SubBytesIns_Inst_Sbox_5_M1), .B0_f (new_AGEMA_signal_7688), .B1_t (new_AGEMA_signal_7689), .B1_f (new_AGEMA_signal_7690), .Z0_t (SubBytesIns_Inst_Sbox_5_M3), .Z0_f (new_AGEMA_signal_8348), .Z1_t (new_AGEMA_signal_8349), .Z1_f (new_AGEMA_signal_8350) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T19), .A0_f (new_AGEMA_signal_7063), .A1_t (new_AGEMA_signal_7064), .A1_f (new_AGEMA_signal_7065), .B0_t (ciphertext_s0_t[40]), .B0_f (ciphertext_s0_f[40]), .B1_t (ciphertext_s1_t[40]), .B1_f (ciphertext_s1_f[40]), .Z0_t (SubBytesIns_Inst_Sbox_5_M4), .Z0_f (new_AGEMA_signal_7691), .Z1_t (new_AGEMA_signal_7692), .Z1_f (new_AGEMA_signal_7693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M4), .A0_f (new_AGEMA_signal_7691), .A1_t (new_AGEMA_signal_7692), .A1_f (new_AGEMA_signal_7693), .B0_t (SubBytesIns_Inst_Sbox_5_M1), .B0_f (new_AGEMA_signal_7688), .B1_t (new_AGEMA_signal_7689), .B1_f (new_AGEMA_signal_7690), .Z0_t (SubBytesIns_Inst_Sbox_5_M5), .Z0_f (new_AGEMA_signal_8351), .Z1_t (new_AGEMA_signal_8352), .Z1_f (new_AGEMA_signal_8353) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T3), .A0_f (new_AGEMA_signal_6502), .A1_t (new_AGEMA_signal_6503), .A1_f (new_AGEMA_signal_6504), .B0_t (SubBytesIns_Inst_Sbox_5_T16), .B0_f (new_AGEMA_signal_7060), .B1_t (new_AGEMA_signal_7061), .B1_f (new_AGEMA_signal_7062), .Z0_t (SubBytesIns_Inst_Sbox_5_M6), .Z0_f (new_AGEMA_signal_7694), .Z1_t (new_AGEMA_signal_7695), .Z1_f (new_AGEMA_signal_7696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T22), .A0_f (new_AGEMA_signal_7066), .A1_t (new_AGEMA_signal_7067), .A1_f (new_AGEMA_signal_7068), .B0_t (SubBytesIns_Inst_Sbox_5_T9), .B0_f (new_AGEMA_signal_7051), .B1_t (new_AGEMA_signal_7052), .B1_f (new_AGEMA_signal_7053), .Z0_t (SubBytesIns_Inst_Sbox_5_M7), .Z0_f (new_AGEMA_signal_7697), .Z1_t (new_AGEMA_signal_7698), .Z1_f (new_AGEMA_signal_7699) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T26), .A0_f (new_AGEMA_signal_7685), .A1_t (new_AGEMA_signal_7686), .A1_f (new_AGEMA_signal_7687), .B0_t (SubBytesIns_Inst_Sbox_5_M6), .B0_f (new_AGEMA_signal_7694), .B1_t (new_AGEMA_signal_7695), .B1_f (new_AGEMA_signal_7696), .Z0_t (SubBytesIns_Inst_Sbox_5_M8), .Z0_f (new_AGEMA_signal_8354), .Z1_t (new_AGEMA_signal_8355), .Z1_f (new_AGEMA_signal_8356) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T20), .A0_f (new_AGEMA_signal_7679), .A1_t (new_AGEMA_signal_7680), .A1_f (new_AGEMA_signal_7681), .B0_t (SubBytesIns_Inst_Sbox_5_T17), .B0_f (new_AGEMA_signal_7676), .B1_t (new_AGEMA_signal_7677), .B1_f (new_AGEMA_signal_7678), .Z0_t (SubBytesIns_Inst_Sbox_5_M9), .Z0_f (new_AGEMA_signal_8357), .Z1_t (new_AGEMA_signal_8358), .Z1_f (new_AGEMA_signal_8359) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M9), .A0_f (new_AGEMA_signal_8357), .A1_t (new_AGEMA_signal_8358), .A1_f (new_AGEMA_signal_8359), .B0_t (SubBytesIns_Inst_Sbox_5_M6), .B0_f (new_AGEMA_signal_7694), .B1_t (new_AGEMA_signal_7695), .B1_f (new_AGEMA_signal_7696), .Z0_t (SubBytesIns_Inst_Sbox_5_M10), .Z0_f (new_AGEMA_signal_8771), .Z1_t (new_AGEMA_signal_8772), .Z1_f (new_AGEMA_signal_8773) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T1), .A0_f (new_AGEMA_signal_6496), .A1_t (new_AGEMA_signal_6497), .A1_f (new_AGEMA_signal_6498), .B0_t (SubBytesIns_Inst_Sbox_5_T15), .B0_f (new_AGEMA_signal_7057), .B1_t (new_AGEMA_signal_7058), .B1_f (new_AGEMA_signal_7059), .Z0_t (SubBytesIns_Inst_Sbox_5_M11), .Z0_f (new_AGEMA_signal_7700), .Z1_t (new_AGEMA_signal_7701), .Z1_f (new_AGEMA_signal_7702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T4), .A0_f (new_AGEMA_signal_6505), .A1_t (new_AGEMA_signal_6506), .A1_f (new_AGEMA_signal_6507), .B0_t (SubBytesIns_Inst_Sbox_5_T27), .B0_f (new_AGEMA_signal_7069), .B1_t (new_AGEMA_signal_7070), .B1_f (new_AGEMA_signal_7071), .Z0_t (SubBytesIns_Inst_Sbox_5_M12), .Z0_f (new_AGEMA_signal_7703), .Z1_t (new_AGEMA_signal_7704), .Z1_f (new_AGEMA_signal_7705) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M12), .A0_f (new_AGEMA_signal_7703), .A1_t (new_AGEMA_signal_7704), .A1_f (new_AGEMA_signal_7705), .B0_t (SubBytesIns_Inst_Sbox_5_M11), .B0_f (new_AGEMA_signal_7700), .B1_t (new_AGEMA_signal_7701), .B1_f (new_AGEMA_signal_7702), .Z0_t (SubBytesIns_Inst_Sbox_5_M13), .Z0_f (new_AGEMA_signal_8360), .Z1_t (new_AGEMA_signal_8361), .Z1_f (new_AGEMA_signal_8362) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T2), .A0_f (new_AGEMA_signal_6499), .A1_t (new_AGEMA_signal_6500), .A1_f (new_AGEMA_signal_6501), .B0_t (SubBytesIns_Inst_Sbox_5_T10), .B0_f (new_AGEMA_signal_7670), .B1_t (new_AGEMA_signal_7671), .B1_f (new_AGEMA_signal_7672), .Z0_t (SubBytesIns_Inst_Sbox_5_M14), .Z0_f (new_AGEMA_signal_8363), .Z1_t (new_AGEMA_signal_8364), .Z1_f (new_AGEMA_signal_8365) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M14), .A0_f (new_AGEMA_signal_8363), .A1_t (new_AGEMA_signal_8364), .A1_f (new_AGEMA_signal_8365), .B0_t (SubBytesIns_Inst_Sbox_5_M11), .B0_f (new_AGEMA_signal_7700), .B1_t (new_AGEMA_signal_7701), .B1_f (new_AGEMA_signal_7702), .Z0_t (SubBytesIns_Inst_Sbox_5_M15), .Z0_f (new_AGEMA_signal_8774), .Z1_t (new_AGEMA_signal_8775), .Z1_f (new_AGEMA_signal_8776) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M3), .A0_f (new_AGEMA_signal_8348), .A1_t (new_AGEMA_signal_8349), .A1_f (new_AGEMA_signal_8350), .B0_t (SubBytesIns_Inst_Sbox_5_M2), .B0_f (new_AGEMA_signal_8345), .B1_t (new_AGEMA_signal_8346), .B1_f (new_AGEMA_signal_8347), .Z0_t (SubBytesIns_Inst_Sbox_5_M16), .Z0_f (new_AGEMA_signal_8777), .Z1_t (new_AGEMA_signal_8778), .Z1_f (new_AGEMA_signal_8779) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M5), .A0_f (new_AGEMA_signal_8351), .A1_t (new_AGEMA_signal_8352), .A1_f (new_AGEMA_signal_8353), .B0_t (SubBytesIns_Inst_Sbox_5_T24), .B0_f (new_AGEMA_signal_8339), .B1_t (new_AGEMA_signal_8340), .B1_f (new_AGEMA_signal_8341), .Z0_t (SubBytesIns_Inst_Sbox_5_M17), .Z0_f (new_AGEMA_signal_8780), .Z1_t (new_AGEMA_signal_8781), .Z1_f (new_AGEMA_signal_8782) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M8), .A0_f (new_AGEMA_signal_8354), .A1_t (new_AGEMA_signal_8355), .A1_f (new_AGEMA_signal_8356), .B0_t (SubBytesIns_Inst_Sbox_5_M7), .B0_f (new_AGEMA_signal_7697), .B1_t (new_AGEMA_signal_7698), .B1_f (new_AGEMA_signal_7699), .Z0_t (SubBytesIns_Inst_Sbox_5_M18), .Z0_f (new_AGEMA_signal_8783), .Z1_t (new_AGEMA_signal_8784), .Z1_f (new_AGEMA_signal_8785) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M10), .A0_f (new_AGEMA_signal_8771), .A1_t (new_AGEMA_signal_8772), .A1_f (new_AGEMA_signal_8773), .B0_t (SubBytesIns_Inst_Sbox_5_M15), .B0_f (new_AGEMA_signal_8774), .B1_t (new_AGEMA_signal_8775), .B1_f (new_AGEMA_signal_8776), .Z0_t (SubBytesIns_Inst_Sbox_5_M19), .Z0_f (new_AGEMA_signal_9044), .Z1_t (new_AGEMA_signal_9045), .Z1_f (new_AGEMA_signal_9046) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M16), .A0_f (new_AGEMA_signal_8777), .A1_t (new_AGEMA_signal_8778), .A1_f (new_AGEMA_signal_8779), .B0_t (SubBytesIns_Inst_Sbox_5_M13), .B0_f (new_AGEMA_signal_8360), .B1_t (new_AGEMA_signal_8361), .B1_f (new_AGEMA_signal_8362), .Z0_t (SubBytesIns_Inst_Sbox_5_M20), .Z0_f (new_AGEMA_signal_9047), .Z1_t (new_AGEMA_signal_9048), .Z1_f (new_AGEMA_signal_9049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M17), .A0_f (new_AGEMA_signal_8780), .A1_t (new_AGEMA_signal_8781), .A1_f (new_AGEMA_signal_8782), .B0_t (SubBytesIns_Inst_Sbox_5_M15), .B0_f (new_AGEMA_signal_8774), .B1_t (new_AGEMA_signal_8775), .B1_f (new_AGEMA_signal_8776), .Z0_t (SubBytesIns_Inst_Sbox_5_M21), .Z0_f (new_AGEMA_signal_9050), .Z1_t (new_AGEMA_signal_9051), .Z1_f (new_AGEMA_signal_9052) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M18), .A0_f (new_AGEMA_signal_8783), .A1_t (new_AGEMA_signal_8784), .A1_f (new_AGEMA_signal_8785), .B0_t (SubBytesIns_Inst_Sbox_5_M13), .B0_f (new_AGEMA_signal_8360), .B1_t (new_AGEMA_signal_8361), .B1_f (new_AGEMA_signal_8362), .Z0_t (SubBytesIns_Inst_Sbox_5_M22), .Z0_f (new_AGEMA_signal_9053), .Z1_t (new_AGEMA_signal_9054), .Z1_f (new_AGEMA_signal_9055) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M19), .A0_f (new_AGEMA_signal_9044), .A1_t (new_AGEMA_signal_9045), .A1_f (new_AGEMA_signal_9046), .B0_t (SubBytesIns_Inst_Sbox_5_T25), .B0_f (new_AGEMA_signal_8342), .B1_t (new_AGEMA_signal_8343), .B1_f (new_AGEMA_signal_8344), .Z0_t (SubBytesIns_Inst_Sbox_5_M23), .Z0_f (new_AGEMA_signal_9284), .Z1_t (new_AGEMA_signal_9285), .Z1_f (new_AGEMA_signal_9286) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M22), .A0_f (new_AGEMA_signal_9053), .A1_t (new_AGEMA_signal_9054), .A1_f (new_AGEMA_signal_9055), .B0_t (SubBytesIns_Inst_Sbox_5_M23), .B0_f (new_AGEMA_signal_9284), .B1_t (new_AGEMA_signal_9285), .B1_f (new_AGEMA_signal_9286), .Z0_t (SubBytesIns_Inst_Sbox_5_M24), .Z0_f (new_AGEMA_signal_9551), .Z1_t (new_AGEMA_signal_9552), .Z1_f (new_AGEMA_signal_9553) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M22), .A0_f (new_AGEMA_signal_9053), .A1_t (new_AGEMA_signal_9054), .A1_f (new_AGEMA_signal_9055), .B0_t (SubBytesIns_Inst_Sbox_5_M20), .B0_f (new_AGEMA_signal_9047), .B1_t (new_AGEMA_signal_9048), .B1_f (new_AGEMA_signal_9049), .Z0_t (SubBytesIns_Inst_Sbox_5_M25), .Z0_f (new_AGEMA_signal_9287), .Z1_t (new_AGEMA_signal_9288), .Z1_f (new_AGEMA_signal_9289) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M21), .A0_f (new_AGEMA_signal_9050), .A1_t (new_AGEMA_signal_9051), .A1_f (new_AGEMA_signal_9052), .B0_t (SubBytesIns_Inst_Sbox_5_M25), .B0_f (new_AGEMA_signal_9287), .B1_t (new_AGEMA_signal_9288), .B1_f (new_AGEMA_signal_9289), .Z0_t (SubBytesIns_Inst_Sbox_5_M26), .Z0_f (new_AGEMA_signal_9554), .Z1_t (new_AGEMA_signal_9555), .Z1_f (new_AGEMA_signal_9556) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M20), .A0_f (new_AGEMA_signal_9047), .A1_t (new_AGEMA_signal_9048), .A1_f (new_AGEMA_signal_9049), .B0_t (SubBytesIns_Inst_Sbox_5_M21), .B0_f (new_AGEMA_signal_9050), .B1_t (new_AGEMA_signal_9051), .B1_f (new_AGEMA_signal_9052), .Z0_t (SubBytesIns_Inst_Sbox_5_M27), .Z0_f (new_AGEMA_signal_9290), .Z1_t (new_AGEMA_signal_9291), .Z1_f (new_AGEMA_signal_9292) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M23), .A0_f (new_AGEMA_signal_9284), .A1_t (new_AGEMA_signal_9285), .A1_f (new_AGEMA_signal_9286), .B0_t (SubBytesIns_Inst_Sbox_5_M25), .B0_f (new_AGEMA_signal_9287), .B1_t (new_AGEMA_signal_9288), .B1_f (new_AGEMA_signal_9289), .Z0_t (SubBytesIns_Inst_Sbox_5_M28), .Z0_f (new_AGEMA_signal_9557), .Z1_t (new_AGEMA_signal_9558), .Z1_f (new_AGEMA_signal_9559) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M28), .A0_f (new_AGEMA_signal_9557), .A1_t (new_AGEMA_signal_9558), .A1_f (new_AGEMA_signal_9559), .B0_t (SubBytesIns_Inst_Sbox_5_M27), .B0_f (new_AGEMA_signal_9290), .B1_t (new_AGEMA_signal_9291), .B1_f (new_AGEMA_signal_9292), .Z0_t (SubBytesIns_Inst_Sbox_5_M29), .Z0_f (new_AGEMA_signal_9851), .Z1_t (new_AGEMA_signal_9852), .Z1_f (new_AGEMA_signal_9853) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M26), .A0_f (new_AGEMA_signal_9554), .A1_t (new_AGEMA_signal_9555), .A1_f (new_AGEMA_signal_9556), .B0_t (SubBytesIns_Inst_Sbox_5_M24), .B0_f (new_AGEMA_signal_9551), .B1_t (new_AGEMA_signal_9552), .B1_f (new_AGEMA_signal_9553), .Z0_t (SubBytesIns_Inst_Sbox_5_M30), .Z0_f (new_AGEMA_signal_9854), .Z1_t (new_AGEMA_signal_9855), .Z1_f (new_AGEMA_signal_9856) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M20), .A0_f (new_AGEMA_signal_9047), .A1_t (new_AGEMA_signal_9048), .A1_f (new_AGEMA_signal_9049), .B0_t (SubBytesIns_Inst_Sbox_5_M23), .B0_f (new_AGEMA_signal_9284), .B1_t (new_AGEMA_signal_9285), .B1_f (new_AGEMA_signal_9286), .Z0_t (SubBytesIns_Inst_Sbox_5_M31), .Z0_f (new_AGEMA_signal_9560), .Z1_t (new_AGEMA_signal_9561), .Z1_f (new_AGEMA_signal_9562) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M27), .A0_f (new_AGEMA_signal_9290), .A1_t (new_AGEMA_signal_9291), .A1_f (new_AGEMA_signal_9292), .B0_t (SubBytesIns_Inst_Sbox_5_M31), .B0_f (new_AGEMA_signal_9560), .B1_t (new_AGEMA_signal_9561), .B1_f (new_AGEMA_signal_9562), .Z0_t (SubBytesIns_Inst_Sbox_5_M32), .Z0_f (new_AGEMA_signal_9857), .Z1_t (new_AGEMA_signal_9858), .Z1_f (new_AGEMA_signal_9859) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M27), .A0_f (new_AGEMA_signal_9290), .A1_t (new_AGEMA_signal_9291), .A1_f (new_AGEMA_signal_9292), .B0_t (SubBytesIns_Inst_Sbox_5_M25), .B0_f (new_AGEMA_signal_9287), .B1_t (new_AGEMA_signal_9288), .B1_f (new_AGEMA_signal_9289), .Z0_t (SubBytesIns_Inst_Sbox_5_M33), .Z0_f (new_AGEMA_signal_9563), .Z1_t (new_AGEMA_signal_9564), .Z1_f (new_AGEMA_signal_9565) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M21), .A0_f (new_AGEMA_signal_9050), .A1_t (new_AGEMA_signal_9051), .A1_f (new_AGEMA_signal_9052), .B0_t (SubBytesIns_Inst_Sbox_5_M22), .B0_f (new_AGEMA_signal_9053), .B1_t (new_AGEMA_signal_9054), .B1_f (new_AGEMA_signal_9055), .Z0_t (SubBytesIns_Inst_Sbox_5_M34), .Z0_f (new_AGEMA_signal_9293), .Z1_t (new_AGEMA_signal_9294), .Z1_f (new_AGEMA_signal_9295) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M24), .A0_f (new_AGEMA_signal_9551), .A1_t (new_AGEMA_signal_9552), .A1_f (new_AGEMA_signal_9553), .B0_t (SubBytesIns_Inst_Sbox_5_M34), .B0_f (new_AGEMA_signal_9293), .B1_t (new_AGEMA_signal_9294), .B1_f (new_AGEMA_signal_9295), .Z0_t (SubBytesIns_Inst_Sbox_5_M35), .Z0_f (new_AGEMA_signal_9860), .Z1_t (new_AGEMA_signal_9861), .Z1_f (new_AGEMA_signal_9862) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M24), .A0_f (new_AGEMA_signal_9551), .A1_t (new_AGEMA_signal_9552), .A1_f (new_AGEMA_signal_9553), .B0_t (SubBytesIns_Inst_Sbox_5_M25), .B0_f (new_AGEMA_signal_9287), .B1_t (new_AGEMA_signal_9288), .B1_f (new_AGEMA_signal_9289), .Z0_t (SubBytesIns_Inst_Sbox_5_M36), .Z0_f (new_AGEMA_signal_9863), .Z1_t (new_AGEMA_signal_9864), .Z1_f (new_AGEMA_signal_9865) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M21), .A0_f (new_AGEMA_signal_9050), .A1_t (new_AGEMA_signal_9051), .A1_f (new_AGEMA_signal_9052), .B0_t (SubBytesIns_Inst_Sbox_5_M29), .B0_f (new_AGEMA_signal_9851), .B1_t (new_AGEMA_signal_9852), .B1_f (new_AGEMA_signal_9853), .Z0_t (SubBytesIns_Inst_Sbox_5_M37), .Z0_f (new_AGEMA_signal_10124), .Z1_t (new_AGEMA_signal_10125), .Z1_f (new_AGEMA_signal_10126) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M32), .A0_f (new_AGEMA_signal_9857), .A1_t (new_AGEMA_signal_9858), .A1_f (new_AGEMA_signal_9859), .B0_t (SubBytesIns_Inst_Sbox_5_M33), .B0_f (new_AGEMA_signal_9563), .B1_t (new_AGEMA_signal_9564), .B1_f (new_AGEMA_signal_9565), .Z0_t (SubBytesIns_Inst_Sbox_5_M38), .Z0_f (new_AGEMA_signal_10127), .Z1_t (new_AGEMA_signal_10128), .Z1_f (new_AGEMA_signal_10129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M23), .A0_f (new_AGEMA_signal_9284), .A1_t (new_AGEMA_signal_9285), .A1_f (new_AGEMA_signal_9286), .B0_t (SubBytesIns_Inst_Sbox_5_M30), .B0_f (new_AGEMA_signal_9854), .B1_t (new_AGEMA_signal_9855), .B1_f (new_AGEMA_signal_9856), .Z0_t (SubBytesIns_Inst_Sbox_5_M39), .Z0_f (new_AGEMA_signal_10130), .Z1_t (new_AGEMA_signal_10131), .Z1_f (new_AGEMA_signal_10132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M35), .A0_f (new_AGEMA_signal_9860), .A1_t (new_AGEMA_signal_9861), .A1_f (new_AGEMA_signal_9862), .B0_t (SubBytesIns_Inst_Sbox_5_M36), .B0_f (new_AGEMA_signal_9863), .B1_t (new_AGEMA_signal_9864), .B1_f (new_AGEMA_signal_9865), .Z0_t (SubBytesIns_Inst_Sbox_5_M40), .Z0_f (new_AGEMA_signal_10133), .Z1_t (new_AGEMA_signal_10134), .Z1_f (new_AGEMA_signal_10135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M38), .A0_f (new_AGEMA_signal_10127), .A1_t (new_AGEMA_signal_10128), .A1_f (new_AGEMA_signal_10129), .B0_t (SubBytesIns_Inst_Sbox_5_M40), .B0_f (new_AGEMA_signal_10133), .B1_t (new_AGEMA_signal_10134), .B1_f (new_AGEMA_signal_10135), .Z0_t (SubBytesIns_Inst_Sbox_5_M41), .Z0_f (new_AGEMA_signal_10580), .Z1_t (new_AGEMA_signal_10581), .Z1_f (new_AGEMA_signal_10582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M37), .A0_f (new_AGEMA_signal_10124), .A1_t (new_AGEMA_signal_10125), .A1_f (new_AGEMA_signal_10126), .B0_t (SubBytesIns_Inst_Sbox_5_M39), .B0_f (new_AGEMA_signal_10130), .B1_t (new_AGEMA_signal_10131), .B1_f (new_AGEMA_signal_10132), .Z0_t (SubBytesIns_Inst_Sbox_5_M42), .Z0_f (new_AGEMA_signal_10583), .Z1_t (new_AGEMA_signal_10584), .Z1_f (new_AGEMA_signal_10585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M37), .A0_f (new_AGEMA_signal_10124), .A1_t (new_AGEMA_signal_10125), .A1_f (new_AGEMA_signal_10126), .B0_t (SubBytesIns_Inst_Sbox_5_M38), .B0_f (new_AGEMA_signal_10127), .B1_t (new_AGEMA_signal_10128), .B1_f (new_AGEMA_signal_10129), .Z0_t (SubBytesIns_Inst_Sbox_5_M43), .Z0_f (new_AGEMA_signal_10586), .Z1_t (new_AGEMA_signal_10587), .Z1_f (new_AGEMA_signal_10588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M39), .A0_f (new_AGEMA_signal_10130), .A1_t (new_AGEMA_signal_10131), .A1_f (new_AGEMA_signal_10132), .B0_t (SubBytesIns_Inst_Sbox_5_M40), .B0_f (new_AGEMA_signal_10133), .B1_t (new_AGEMA_signal_10134), .B1_f (new_AGEMA_signal_10135), .Z0_t (SubBytesIns_Inst_Sbox_5_M44), .Z0_f (new_AGEMA_signal_10589), .Z1_t (new_AGEMA_signal_10590), .Z1_f (new_AGEMA_signal_10591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M42), .A0_f (new_AGEMA_signal_10583), .A1_t (new_AGEMA_signal_10584), .A1_f (new_AGEMA_signal_10585), .B0_t (SubBytesIns_Inst_Sbox_5_M41), .B0_f (new_AGEMA_signal_10580), .B1_t (new_AGEMA_signal_10581), .B1_f (new_AGEMA_signal_10582), .Z0_t (SubBytesIns_Inst_Sbox_5_M45), .Z0_f (new_AGEMA_signal_11300), .Z1_t (new_AGEMA_signal_11301), .Z1_f (new_AGEMA_signal_11302) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M44), .A0_f (new_AGEMA_signal_10589), .A1_t (new_AGEMA_signal_10590), .A1_f (new_AGEMA_signal_10591), .B0_t (SubBytesIns_Inst_Sbox_5_T6), .B0_f (new_AGEMA_signal_7048), .B1_t (new_AGEMA_signal_7049), .B1_f (new_AGEMA_signal_7050), .Z0_t (SubBytesIns_Inst_Sbox_5_M46), .Z0_f (new_AGEMA_signal_11303), .Z1_t (new_AGEMA_signal_11304), .Z1_f (new_AGEMA_signal_11305) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M40), .A0_f (new_AGEMA_signal_10133), .A1_t (new_AGEMA_signal_10134), .A1_f (new_AGEMA_signal_10135), .B0_t (SubBytesIns_Inst_Sbox_5_T8), .B0_f (new_AGEMA_signal_7667), .B1_t (new_AGEMA_signal_7668), .B1_f (new_AGEMA_signal_7669), .Z0_t (SubBytesIns_Inst_Sbox_5_M47), .Z0_f (new_AGEMA_signal_10592), .Z1_t (new_AGEMA_signal_10593), .Z1_f (new_AGEMA_signal_10594) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M39), .A0_f (new_AGEMA_signal_10130), .A1_t (new_AGEMA_signal_10131), .A1_f (new_AGEMA_signal_10132), .B0_t (ciphertext_s0_t[40]), .B0_f (ciphertext_s0_f[40]), .B1_t (ciphertext_s1_t[40]), .B1_f (ciphertext_s1_f[40]), .Z0_t (SubBytesIns_Inst_Sbox_5_M48), .Z0_f (new_AGEMA_signal_10595), .Z1_t (new_AGEMA_signal_10596), .Z1_f (new_AGEMA_signal_10597) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M43), .A0_f (new_AGEMA_signal_10586), .A1_t (new_AGEMA_signal_10587), .A1_f (new_AGEMA_signal_10588), .B0_t (SubBytesIns_Inst_Sbox_5_T16), .B0_f (new_AGEMA_signal_7060), .B1_t (new_AGEMA_signal_7061), .B1_f (new_AGEMA_signal_7062), .Z0_t (SubBytesIns_Inst_Sbox_5_M49), .Z0_f (new_AGEMA_signal_11306), .Z1_t (new_AGEMA_signal_11307), .Z1_f (new_AGEMA_signal_11308) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M38), .A0_f (new_AGEMA_signal_10127), .A1_t (new_AGEMA_signal_10128), .A1_f (new_AGEMA_signal_10129), .B0_t (SubBytesIns_Inst_Sbox_5_T9), .B0_f (new_AGEMA_signal_7051), .B1_t (new_AGEMA_signal_7052), .B1_f (new_AGEMA_signal_7053), .Z0_t (SubBytesIns_Inst_Sbox_5_M50), .Z0_f (new_AGEMA_signal_10598), .Z1_t (new_AGEMA_signal_10599), .Z1_f (new_AGEMA_signal_10600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M37), .A0_f (new_AGEMA_signal_10124), .A1_t (new_AGEMA_signal_10125), .A1_f (new_AGEMA_signal_10126), .B0_t (SubBytesIns_Inst_Sbox_5_T17), .B0_f (new_AGEMA_signal_7676), .B1_t (new_AGEMA_signal_7677), .B1_f (new_AGEMA_signal_7678), .Z0_t (SubBytesIns_Inst_Sbox_5_M51), .Z0_f (new_AGEMA_signal_10601), .Z1_t (new_AGEMA_signal_10602), .Z1_f (new_AGEMA_signal_10603) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M42), .A0_f (new_AGEMA_signal_10583), .A1_t (new_AGEMA_signal_10584), .A1_f (new_AGEMA_signal_10585), .B0_t (SubBytesIns_Inst_Sbox_5_T15), .B0_f (new_AGEMA_signal_7057), .B1_t (new_AGEMA_signal_7058), .B1_f (new_AGEMA_signal_7059), .Z0_t (SubBytesIns_Inst_Sbox_5_M52), .Z0_f (new_AGEMA_signal_11309), .Z1_t (new_AGEMA_signal_11310), .Z1_f (new_AGEMA_signal_11311) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M45), .A0_f (new_AGEMA_signal_11300), .A1_t (new_AGEMA_signal_11301), .A1_f (new_AGEMA_signal_11302), .B0_t (SubBytesIns_Inst_Sbox_5_T27), .B0_f (new_AGEMA_signal_7069), .B1_t (new_AGEMA_signal_7070), .B1_f (new_AGEMA_signal_7071), .Z0_t (SubBytesIns_Inst_Sbox_5_M53), .Z0_f (new_AGEMA_signal_11966), .Z1_t (new_AGEMA_signal_11967), .Z1_f (new_AGEMA_signal_11968) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M41), .A0_f (new_AGEMA_signal_10580), .A1_t (new_AGEMA_signal_10581), .A1_f (new_AGEMA_signal_10582), .B0_t (SubBytesIns_Inst_Sbox_5_T10), .B0_f (new_AGEMA_signal_7670), .B1_t (new_AGEMA_signal_7671), .B1_f (new_AGEMA_signal_7672), .Z0_t (SubBytesIns_Inst_Sbox_5_M54), .Z0_f (new_AGEMA_signal_11312), .Z1_t (new_AGEMA_signal_11313), .Z1_f (new_AGEMA_signal_11314) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M44), .A0_f (new_AGEMA_signal_10589), .A1_t (new_AGEMA_signal_10590), .A1_f (new_AGEMA_signal_10591), .B0_t (SubBytesIns_Inst_Sbox_5_T13), .B0_f (new_AGEMA_signal_7054), .B1_t (new_AGEMA_signal_7055), .B1_f (new_AGEMA_signal_7056), .Z0_t (SubBytesIns_Inst_Sbox_5_M55), .Z0_f (new_AGEMA_signal_11315), .Z1_t (new_AGEMA_signal_11316), .Z1_f (new_AGEMA_signal_11317) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M40), .A0_f (new_AGEMA_signal_10133), .A1_t (new_AGEMA_signal_10134), .A1_f (new_AGEMA_signal_10135), .B0_t (SubBytesIns_Inst_Sbox_5_T23), .B0_f (new_AGEMA_signal_7682), .B1_t (new_AGEMA_signal_7683), .B1_f (new_AGEMA_signal_7684), .Z0_t (SubBytesIns_Inst_Sbox_5_M56), .Z0_f (new_AGEMA_signal_10604), .Z1_t (new_AGEMA_signal_10605), .Z1_f (new_AGEMA_signal_10606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M39), .A0_f (new_AGEMA_signal_10130), .A1_t (new_AGEMA_signal_10131), .A1_f (new_AGEMA_signal_10132), .B0_t (SubBytesIns_Inst_Sbox_5_T19), .B0_f (new_AGEMA_signal_7063), .B1_t (new_AGEMA_signal_7064), .B1_f (new_AGEMA_signal_7065), .Z0_t (SubBytesIns_Inst_Sbox_5_M57), .Z0_f (new_AGEMA_signal_10607), .Z1_t (new_AGEMA_signal_10608), .Z1_f (new_AGEMA_signal_10609) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M43), .A0_f (new_AGEMA_signal_10586), .A1_t (new_AGEMA_signal_10587), .A1_f (new_AGEMA_signal_10588), .B0_t (SubBytesIns_Inst_Sbox_5_T3), .B0_f (new_AGEMA_signal_6502), .B1_t (new_AGEMA_signal_6503), .B1_f (new_AGEMA_signal_6504), .Z0_t (SubBytesIns_Inst_Sbox_5_M58), .Z0_f (new_AGEMA_signal_11318), .Z1_t (new_AGEMA_signal_11319), .Z1_f (new_AGEMA_signal_11320) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M38), .A0_f (new_AGEMA_signal_10127), .A1_t (new_AGEMA_signal_10128), .A1_f (new_AGEMA_signal_10129), .B0_t (SubBytesIns_Inst_Sbox_5_T22), .B0_f (new_AGEMA_signal_7066), .B1_t (new_AGEMA_signal_7067), .B1_f (new_AGEMA_signal_7068), .Z0_t (SubBytesIns_Inst_Sbox_5_M59), .Z0_f (new_AGEMA_signal_10610), .Z1_t (new_AGEMA_signal_10611), .Z1_f (new_AGEMA_signal_10612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M37), .A0_f (new_AGEMA_signal_10124), .A1_t (new_AGEMA_signal_10125), .A1_f (new_AGEMA_signal_10126), .B0_t (SubBytesIns_Inst_Sbox_5_T20), .B0_f (new_AGEMA_signal_7679), .B1_t (new_AGEMA_signal_7680), .B1_f (new_AGEMA_signal_7681), .Z0_t (SubBytesIns_Inst_Sbox_5_M60), .Z0_f (new_AGEMA_signal_10613), .Z1_t (new_AGEMA_signal_10614), .Z1_f (new_AGEMA_signal_10615) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M42), .A0_f (new_AGEMA_signal_10583), .A1_t (new_AGEMA_signal_10584), .A1_f (new_AGEMA_signal_10585), .B0_t (SubBytesIns_Inst_Sbox_5_T1), .B0_f (new_AGEMA_signal_6496), .B1_t (new_AGEMA_signal_6497), .B1_f (new_AGEMA_signal_6498), .Z0_t (SubBytesIns_Inst_Sbox_5_M61), .Z0_f (new_AGEMA_signal_11321), .Z1_t (new_AGEMA_signal_11322), .Z1_f (new_AGEMA_signal_11323) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M45), .A0_f (new_AGEMA_signal_11300), .A1_t (new_AGEMA_signal_11301), .A1_f (new_AGEMA_signal_11302), .B0_t (SubBytesIns_Inst_Sbox_5_T4), .B0_f (new_AGEMA_signal_6505), .B1_t (new_AGEMA_signal_6506), .B1_f (new_AGEMA_signal_6507), .Z0_t (SubBytesIns_Inst_Sbox_5_M62), .Z0_f (new_AGEMA_signal_11969), .Z1_t (new_AGEMA_signal_11970), .Z1_f (new_AGEMA_signal_11971) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M41), .A0_f (new_AGEMA_signal_10580), .A1_t (new_AGEMA_signal_10581), .A1_f (new_AGEMA_signal_10582), .B0_t (SubBytesIns_Inst_Sbox_5_T2), .B0_f (new_AGEMA_signal_6499), .B1_t (new_AGEMA_signal_6500), .B1_f (new_AGEMA_signal_6501), .Z0_t (SubBytesIns_Inst_Sbox_5_M63), .Z0_f (new_AGEMA_signal_11324), .Z1_t (new_AGEMA_signal_11325), .Z1_f (new_AGEMA_signal_11326) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M61), .A0_f (new_AGEMA_signal_11321), .A1_t (new_AGEMA_signal_11322), .A1_f (new_AGEMA_signal_11323), .B0_t (SubBytesIns_Inst_Sbox_5_M62), .B0_f (new_AGEMA_signal_11969), .B1_t (new_AGEMA_signal_11970), .B1_f (new_AGEMA_signal_11971), .Z0_t (SubBytesIns_Inst_Sbox_5_L0), .Z0_f (new_AGEMA_signal_12539), .Z1_t (new_AGEMA_signal_12540), .Z1_f (new_AGEMA_signal_12541) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M50), .A0_f (new_AGEMA_signal_10598), .A1_t (new_AGEMA_signal_10599), .A1_f (new_AGEMA_signal_10600), .B0_t (SubBytesIns_Inst_Sbox_5_M56), .B0_f (new_AGEMA_signal_10604), .B1_t (new_AGEMA_signal_10605), .B1_f (new_AGEMA_signal_10606), .Z0_t (SubBytesIns_Inst_Sbox_5_L1), .Z0_f (new_AGEMA_signal_11327), .Z1_t (new_AGEMA_signal_11328), .Z1_f (new_AGEMA_signal_11329) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M46), .A0_f (new_AGEMA_signal_11303), .A1_t (new_AGEMA_signal_11304), .A1_f (new_AGEMA_signal_11305), .B0_t (SubBytesIns_Inst_Sbox_5_M48), .B0_f (new_AGEMA_signal_10595), .B1_t (new_AGEMA_signal_10596), .B1_f (new_AGEMA_signal_10597), .Z0_t (SubBytesIns_Inst_Sbox_5_L2), .Z0_f (new_AGEMA_signal_11972), .Z1_t (new_AGEMA_signal_11973), .Z1_f (new_AGEMA_signal_11974) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M47), .A0_f (new_AGEMA_signal_10592), .A1_t (new_AGEMA_signal_10593), .A1_f (new_AGEMA_signal_10594), .B0_t (SubBytesIns_Inst_Sbox_5_M55), .B0_f (new_AGEMA_signal_11315), .B1_t (new_AGEMA_signal_11316), .B1_f (new_AGEMA_signal_11317), .Z0_t (SubBytesIns_Inst_Sbox_5_L3), .Z0_f (new_AGEMA_signal_11975), .Z1_t (new_AGEMA_signal_11976), .Z1_f (new_AGEMA_signal_11977) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M54), .A0_f (new_AGEMA_signal_11312), .A1_t (new_AGEMA_signal_11313), .A1_f (new_AGEMA_signal_11314), .B0_t (SubBytesIns_Inst_Sbox_5_M58), .B0_f (new_AGEMA_signal_11318), .B1_t (new_AGEMA_signal_11319), .B1_f (new_AGEMA_signal_11320), .Z0_t (SubBytesIns_Inst_Sbox_5_L4), .Z0_f (new_AGEMA_signal_11978), .Z1_t (new_AGEMA_signal_11979), .Z1_f (new_AGEMA_signal_11980) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M49), .A0_f (new_AGEMA_signal_11306), .A1_t (new_AGEMA_signal_11307), .A1_f (new_AGEMA_signal_11308), .B0_t (SubBytesIns_Inst_Sbox_5_M61), .B0_f (new_AGEMA_signal_11321), .B1_t (new_AGEMA_signal_11322), .B1_f (new_AGEMA_signal_11323), .Z0_t (SubBytesIns_Inst_Sbox_5_L5), .Z0_f (new_AGEMA_signal_11981), .Z1_t (new_AGEMA_signal_11982), .Z1_f (new_AGEMA_signal_11983) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M62), .A0_f (new_AGEMA_signal_11969), .A1_t (new_AGEMA_signal_11970), .A1_f (new_AGEMA_signal_11971), .B0_t (SubBytesIns_Inst_Sbox_5_L5), .B0_f (new_AGEMA_signal_11981), .B1_t (new_AGEMA_signal_11982), .B1_f (new_AGEMA_signal_11983), .Z0_t (SubBytesIns_Inst_Sbox_5_L6), .Z0_f (new_AGEMA_signal_12542), .Z1_t (new_AGEMA_signal_12543), .Z1_f (new_AGEMA_signal_12544) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M46), .A0_f (new_AGEMA_signal_11303), .A1_t (new_AGEMA_signal_11304), .A1_f (new_AGEMA_signal_11305), .B0_t (SubBytesIns_Inst_Sbox_5_L3), .B0_f (new_AGEMA_signal_11975), .B1_t (new_AGEMA_signal_11976), .B1_f (new_AGEMA_signal_11977), .Z0_t (SubBytesIns_Inst_Sbox_5_L7), .Z0_f (new_AGEMA_signal_12545), .Z1_t (new_AGEMA_signal_12546), .Z1_f (new_AGEMA_signal_12547) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M51), .A0_f (new_AGEMA_signal_10601), .A1_t (new_AGEMA_signal_10602), .A1_f (new_AGEMA_signal_10603), .B0_t (SubBytesIns_Inst_Sbox_5_M59), .B0_f (new_AGEMA_signal_10610), .B1_t (new_AGEMA_signal_10611), .B1_f (new_AGEMA_signal_10612), .Z0_t (SubBytesIns_Inst_Sbox_5_L8), .Z0_f (new_AGEMA_signal_11330), .Z1_t (new_AGEMA_signal_11331), .Z1_f (new_AGEMA_signal_11332) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M52), .A0_f (new_AGEMA_signal_11309), .A1_t (new_AGEMA_signal_11310), .A1_f (new_AGEMA_signal_11311), .B0_t (SubBytesIns_Inst_Sbox_5_M53), .B0_f (new_AGEMA_signal_11966), .B1_t (new_AGEMA_signal_11967), .B1_f (new_AGEMA_signal_11968), .Z0_t (SubBytesIns_Inst_Sbox_5_L9), .Z0_f (new_AGEMA_signal_12548), .Z1_t (new_AGEMA_signal_12549), .Z1_f (new_AGEMA_signal_12550) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M53), .A0_f (new_AGEMA_signal_11966), .A1_t (new_AGEMA_signal_11967), .A1_f (new_AGEMA_signal_11968), .B0_t (SubBytesIns_Inst_Sbox_5_L4), .B0_f (new_AGEMA_signal_11978), .B1_t (new_AGEMA_signal_11979), .B1_f (new_AGEMA_signal_11980), .Z0_t (SubBytesIns_Inst_Sbox_5_L10), .Z0_f (new_AGEMA_signal_12551), .Z1_t (new_AGEMA_signal_12552), .Z1_f (new_AGEMA_signal_12553) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M60), .A0_f (new_AGEMA_signal_10613), .A1_t (new_AGEMA_signal_10614), .A1_f (new_AGEMA_signal_10615), .B0_t (SubBytesIns_Inst_Sbox_5_L2), .B0_f (new_AGEMA_signal_11972), .B1_t (new_AGEMA_signal_11973), .B1_f (new_AGEMA_signal_11974), .Z0_t (SubBytesIns_Inst_Sbox_5_L11), .Z0_f (new_AGEMA_signal_12554), .Z1_t (new_AGEMA_signal_12555), .Z1_f (new_AGEMA_signal_12556) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M48), .A0_f (new_AGEMA_signal_10595), .A1_t (new_AGEMA_signal_10596), .A1_f (new_AGEMA_signal_10597), .B0_t (SubBytesIns_Inst_Sbox_5_M51), .B0_f (new_AGEMA_signal_10601), .B1_t (new_AGEMA_signal_10602), .B1_f (new_AGEMA_signal_10603), .Z0_t (SubBytesIns_Inst_Sbox_5_L12), .Z0_f (new_AGEMA_signal_11333), .Z1_t (new_AGEMA_signal_11334), .Z1_f (new_AGEMA_signal_11335) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M50), .A0_f (new_AGEMA_signal_10598), .A1_t (new_AGEMA_signal_10599), .A1_f (new_AGEMA_signal_10600), .B0_t (SubBytesIns_Inst_Sbox_5_L0), .B0_f (new_AGEMA_signal_12539), .B1_t (new_AGEMA_signal_12540), .B1_f (new_AGEMA_signal_12541), .Z0_t (SubBytesIns_Inst_Sbox_5_L13), .Z0_f (new_AGEMA_signal_13133), .Z1_t (new_AGEMA_signal_13134), .Z1_f (new_AGEMA_signal_13135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M52), .A0_f (new_AGEMA_signal_11309), .A1_t (new_AGEMA_signal_11310), .A1_f (new_AGEMA_signal_11311), .B0_t (SubBytesIns_Inst_Sbox_5_M61), .B0_f (new_AGEMA_signal_11321), .B1_t (new_AGEMA_signal_11322), .B1_f (new_AGEMA_signal_11323), .Z0_t (SubBytesIns_Inst_Sbox_5_L14), .Z0_f (new_AGEMA_signal_11984), .Z1_t (new_AGEMA_signal_11985), .Z1_f (new_AGEMA_signal_11986) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M55), .A0_f (new_AGEMA_signal_11315), .A1_t (new_AGEMA_signal_11316), .A1_f (new_AGEMA_signal_11317), .B0_t (SubBytesIns_Inst_Sbox_5_L1), .B0_f (new_AGEMA_signal_11327), .B1_t (new_AGEMA_signal_11328), .B1_f (new_AGEMA_signal_11329), .Z0_t (SubBytesIns_Inst_Sbox_5_L15), .Z0_f (new_AGEMA_signal_11987), .Z1_t (new_AGEMA_signal_11988), .Z1_f (new_AGEMA_signal_11989) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M56), .A0_f (new_AGEMA_signal_10604), .A1_t (new_AGEMA_signal_10605), .A1_f (new_AGEMA_signal_10606), .B0_t (SubBytesIns_Inst_Sbox_5_L0), .B0_f (new_AGEMA_signal_12539), .B1_t (new_AGEMA_signal_12540), .B1_f (new_AGEMA_signal_12541), .Z0_t (SubBytesIns_Inst_Sbox_5_L16), .Z0_f (new_AGEMA_signal_13136), .Z1_t (new_AGEMA_signal_13137), .Z1_f (new_AGEMA_signal_13138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M57), .A0_f (new_AGEMA_signal_10607), .A1_t (new_AGEMA_signal_10608), .A1_f (new_AGEMA_signal_10609), .B0_t (SubBytesIns_Inst_Sbox_5_L1), .B0_f (new_AGEMA_signal_11327), .B1_t (new_AGEMA_signal_11328), .B1_f (new_AGEMA_signal_11329), .Z0_t (SubBytesIns_Inst_Sbox_5_L17), .Z0_f (new_AGEMA_signal_11990), .Z1_t (new_AGEMA_signal_11991), .Z1_f (new_AGEMA_signal_11992) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M58), .A0_f (new_AGEMA_signal_11318), .A1_t (new_AGEMA_signal_11319), .A1_f (new_AGEMA_signal_11320), .B0_t (SubBytesIns_Inst_Sbox_5_L8), .B0_f (new_AGEMA_signal_11330), .B1_t (new_AGEMA_signal_11331), .B1_f (new_AGEMA_signal_11332), .Z0_t (SubBytesIns_Inst_Sbox_5_L18), .Z0_f (new_AGEMA_signal_11993), .Z1_t (new_AGEMA_signal_11994), .Z1_f (new_AGEMA_signal_11995) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M63), .A0_f (new_AGEMA_signal_11324), .A1_t (new_AGEMA_signal_11325), .A1_f (new_AGEMA_signal_11326), .B0_t (SubBytesIns_Inst_Sbox_5_L4), .B0_f (new_AGEMA_signal_11978), .B1_t (new_AGEMA_signal_11979), .B1_f (new_AGEMA_signal_11980), .Z0_t (SubBytesIns_Inst_Sbox_5_L19), .Z0_f (new_AGEMA_signal_12557), .Z1_t (new_AGEMA_signal_12558), .Z1_f (new_AGEMA_signal_12559) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L0), .A0_f (new_AGEMA_signal_12539), .A1_t (new_AGEMA_signal_12540), .A1_f (new_AGEMA_signal_12541), .B0_t (SubBytesIns_Inst_Sbox_5_L1), .B0_f (new_AGEMA_signal_11327), .B1_t (new_AGEMA_signal_11328), .B1_f (new_AGEMA_signal_11329), .Z0_t (SubBytesIns_Inst_Sbox_5_L20), .Z0_f (new_AGEMA_signal_13139), .Z1_t (new_AGEMA_signal_13140), .Z1_f (new_AGEMA_signal_13141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L1), .A0_f (new_AGEMA_signal_11327), .A1_t (new_AGEMA_signal_11328), .A1_f (new_AGEMA_signal_11329), .B0_t (SubBytesIns_Inst_Sbox_5_L7), .B0_f (new_AGEMA_signal_12545), .B1_t (new_AGEMA_signal_12546), .B1_f (new_AGEMA_signal_12547), .Z0_t (SubBytesIns_Inst_Sbox_5_L21), .Z0_f (new_AGEMA_signal_13142), .Z1_t (new_AGEMA_signal_13143), .Z1_f (new_AGEMA_signal_13144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L3), .A0_f (new_AGEMA_signal_11975), .A1_t (new_AGEMA_signal_11976), .A1_f (new_AGEMA_signal_11977), .B0_t (SubBytesIns_Inst_Sbox_5_L12), .B0_f (new_AGEMA_signal_11333), .B1_t (new_AGEMA_signal_11334), .B1_f (new_AGEMA_signal_11335), .Z0_t (SubBytesIns_Inst_Sbox_5_L22), .Z0_f (new_AGEMA_signal_12560), .Z1_t (new_AGEMA_signal_12561), .Z1_f (new_AGEMA_signal_12562) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L18), .A0_f (new_AGEMA_signal_11993), .A1_t (new_AGEMA_signal_11994), .A1_f (new_AGEMA_signal_11995), .B0_t (SubBytesIns_Inst_Sbox_5_L2), .B0_f (new_AGEMA_signal_11972), .B1_t (new_AGEMA_signal_11973), .B1_f (new_AGEMA_signal_11974), .Z0_t (SubBytesIns_Inst_Sbox_5_L23), .Z0_f (new_AGEMA_signal_12563), .Z1_t (new_AGEMA_signal_12564), .Z1_f (new_AGEMA_signal_12565) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L15), .A0_f (new_AGEMA_signal_11987), .A1_t (new_AGEMA_signal_11988), .A1_f (new_AGEMA_signal_11989), .B0_t (SubBytesIns_Inst_Sbox_5_L9), .B0_f (new_AGEMA_signal_12548), .B1_t (new_AGEMA_signal_12549), .B1_f (new_AGEMA_signal_12550), .Z0_t (SubBytesIns_Inst_Sbox_5_L24), .Z0_f (new_AGEMA_signal_13145), .Z1_t (new_AGEMA_signal_13146), .Z1_f (new_AGEMA_signal_13147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L6), .A0_f (new_AGEMA_signal_12542), .A1_t (new_AGEMA_signal_12543), .A1_f (new_AGEMA_signal_12544), .B0_t (SubBytesIns_Inst_Sbox_5_L10), .B0_f (new_AGEMA_signal_12551), .B1_t (new_AGEMA_signal_12552), .B1_f (new_AGEMA_signal_12553), .Z0_t (SubBytesIns_Inst_Sbox_5_L25), .Z0_f (new_AGEMA_signal_13148), .Z1_t (new_AGEMA_signal_13149), .Z1_f (new_AGEMA_signal_13150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L7), .A0_f (new_AGEMA_signal_12545), .A1_t (new_AGEMA_signal_12546), .A1_f (new_AGEMA_signal_12547), .B0_t (SubBytesIns_Inst_Sbox_5_L9), .B0_f (new_AGEMA_signal_12548), .B1_t (new_AGEMA_signal_12549), .B1_f (new_AGEMA_signal_12550), .Z0_t (SubBytesIns_Inst_Sbox_5_L26), .Z0_f (new_AGEMA_signal_13151), .Z1_t (new_AGEMA_signal_13152), .Z1_f (new_AGEMA_signal_13153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L8), .A0_f (new_AGEMA_signal_11330), .A1_t (new_AGEMA_signal_11331), .A1_f (new_AGEMA_signal_11332), .B0_t (SubBytesIns_Inst_Sbox_5_L10), .B0_f (new_AGEMA_signal_12551), .B1_t (new_AGEMA_signal_12552), .B1_f (new_AGEMA_signal_12553), .Z0_t (SubBytesIns_Inst_Sbox_5_L27), .Z0_f (new_AGEMA_signal_13154), .Z1_t (new_AGEMA_signal_13155), .Z1_f (new_AGEMA_signal_13156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L11), .A0_f (new_AGEMA_signal_12554), .A1_t (new_AGEMA_signal_12555), .A1_f (new_AGEMA_signal_12556), .B0_t (SubBytesIns_Inst_Sbox_5_L14), .B0_f (new_AGEMA_signal_11984), .B1_t (new_AGEMA_signal_11985), .B1_f (new_AGEMA_signal_11986), .Z0_t (SubBytesIns_Inst_Sbox_5_L28), .Z0_f (new_AGEMA_signal_13157), .Z1_t (new_AGEMA_signal_13158), .Z1_f (new_AGEMA_signal_13159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L11), .A0_f (new_AGEMA_signal_12554), .A1_t (new_AGEMA_signal_12555), .A1_f (new_AGEMA_signal_12556), .B0_t (SubBytesIns_Inst_Sbox_5_L17), .B0_f (new_AGEMA_signal_11990), .B1_t (new_AGEMA_signal_11991), .B1_f (new_AGEMA_signal_11992), .Z0_t (SubBytesIns_Inst_Sbox_5_L29), .Z0_f (new_AGEMA_signal_13160), .Z1_t (new_AGEMA_signal_13161), .Z1_f (new_AGEMA_signal_13162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L6), .A0_f (new_AGEMA_signal_12542), .A1_t (new_AGEMA_signal_12543), .A1_f (new_AGEMA_signal_12544), .B0_t (SubBytesIns_Inst_Sbox_5_L24), .B0_f (new_AGEMA_signal_13145), .B1_t (new_AGEMA_signal_13146), .B1_f (new_AGEMA_signal_13147), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .Z0_f (new_AGEMA_signal_13745), .Z1_t (new_AGEMA_signal_13746), .Z1_f (new_AGEMA_signal_13747) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L16), .A0_f (new_AGEMA_signal_13136), .A1_t (new_AGEMA_signal_13137), .A1_f (new_AGEMA_signal_13138), .B0_t (SubBytesIns_Inst_Sbox_5_L26), .B0_f (new_AGEMA_signal_13151), .B1_t (new_AGEMA_signal_13152), .B1_f (new_AGEMA_signal_13153), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .Z0_f (new_AGEMA_signal_13748), .Z1_t (new_AGEMA_signal_13749), .Z1_f (new_AGEMA_signal_13750) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L19), .A0_f (new_AGEMA_signal_12557), .A1_t (new_AGEMA_signal_12558), .A1_f (new_AGEMA_signal_12559), .B0_t (SubBytesIns_Inst_Sbox_5_L28), .B0_f (new_AGEMA_signal_13157), .B1_t (new_AGEMA_signal_13158), .B1_f (new_AGEMA_signal_13159), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .Z0_f (new_AGEMA_signal_13751), .Z1_t (new_AGEMA_signal_13752), .Z1_f (new_AGEMA_signal_13753) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L6), .A0_f (new_AGEMA_signal_12542), .A1_t (new_AGEMA_signal_12543), .A1_f (new_AGEMA_signal_12544), .B0_t (SubBytesIns_Inst_Sbox_5_L21), .B0_f (new_AGEMA_signal_13142), .B1_t (new_AGEMA_signal_13143), .B1_f (new_AGEMA_signal_13144), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .Z0_f (new_AGEMA_signal_13754), .Z1_t (new_AGEMA_signal_13755), .Z1_f (new_AGEMA_signal_13756) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L20), .A0_f (new_AGEMA_signal_13139), .A1_t (new_AGEMA_signal_13140), .A1_f (new_AGEMA_signal_13141), .B0_t (SubBytesIns_Inst_Sbox_5_L22), .B0_f (new_AGEMA_signal_12560), .B1_t (new_AGEMA_signal_12561), .B1_f (new_AGEMA_signal_12562), .Z0_t (MixColumnsInput[107]), .Z0_f (new_AGEMA_signal_13757), .Z1_t (new_AGEMA_signal_13758), .Z1_f (new_AGEMA_signal_13759) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L25), .A0_f (new_AGEMA_signal_13148), .A1_t (new_AGEMA_signal_13149), .A1_f (new_AGEMA_signal_13150), .B0_t (SubBytesIns_Inst_Sbox_5_L29), .B0_f (new_AGEMA_signal_13160), .B1_t (new_AGEMA_signal_13161), .B1_f (new_AGEMA_signal_13162), .Z0_t (MixColumnsInput[106]), .Z0_f (new_AGEMA_signal_13760), .Z1_t (new_AGEMA_signal_13761), .Z1_f (new_AGEMA_signal_13762) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L13), .A0_f (new_AGEMA_signal_13133), .A1_t (new_AGEMA_signal_13134), .A1_f (new_AGEMA_signal_13135), .B0_t (SubBytesIns_Inst_Sbox_5_L27), .B0_f (new_AGEMA_signal_13154), .B1_t (new_AGEMA_signal_13155), .B1_f (new_AGEMA_signal_13156), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .Z0_f (new_AGEMA_signal_13763), .Z1_t (new_AGEMA_signal_13764), .Z1_f (new_AGEMA_signal_13765) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L6), .A0_f (new_AGEMA_signal_12542), .A1_t (new_AGEMA_signal_12543), .A1_f (new_AGEMA_signal_12544), .B0_t (SubBytesIns_Inst_Sbox_5_L23), .B0_f (new_AGEMA_signal_12563), .B1_t (new_AGEMA_signal_12564), .B1_f (new_AGEMA_signal_12565), .Z0_t (MixColumnsInput[104]), .Z0_f (new_AGEMA_signal_13163), .Z1_t (new_AGEMA_signal_13164), .Z1_f (new_AGEMA_signal_13165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[55]), .A0_f (ciphertext_s0_f[55]), .A1_t (ciphertext_s1_t[55]), .A1_f (ciphertext_s1_f[55]), .B0_t (ciphertext_s0_t[52]), .B0_f (ciphertext_s0_f[52]), .B1_t (ciphertext_s1_t[52]), .B1_f (ciphertext_s1_f[52]), .Z0_t (SubBytesIns_Inst_Sbox_6_T1), .Z0_f (new_AGEMA_signal_6526), .Z1_t (new_AGEMA_signal_6527), .Z1_f (new_AGEMA_signal_6528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[55]), .A0_f (ciphertext_s0_f[55]), .A1_t (ciphertext_s1_t[55]), .A1_f (ciphertext_s1_f[55]), .B0_t (ciphertext_s0_t[50]), .B0_f (ciphertext_s0_f[50]), .B1_t (ciphertext_s1_t[50]), .B1_f (ciphertext_s1_f[50]), .Z0_t (SubBytesIns_Inst_Sbox_6_T2), .Z0_f (new_AGEMA_signal_6529), .Z1_t (new_AGEMA_signal_6530), .Z1_f (new_AGEMA_signal_6531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[55]), .A0_f (ciphertext_s0_f[55]), .A1_t (ciphertext_s1_t[55]), .A1_f (ciphertext_s1_f[55]), .B0_t (ciphertext_s0_t[49]), .B0_f (ciphertext_s0_f[49]), .B1_t (ciphertext_s1_t[49]), .B1_f (ciphertext_s1_f[49]), .Z0_t (SubBytesIns_Inst_Sbox_6_T3), .Z0_f (new_AGEMA_signal_6532), .Z1_t (new_AGEMA_signal_6533), .Z1_f (new_AGEMA_signal_6534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[52]), .A0_f (ciphertext_s0_f[52]), .A1_t (ciphertext_s1_t[52]), .A1_f (ciphertext_s1_f[52]), .B0_t (ciphertext_s0_t[50]), .B0_f (ciphertext_s0_f[50]), .B1_t (ciphertext_s1_t[50]), .B1_f (ciphertext_s1_f[50]), .Z0_t (SubBytesIns_Inst_Sbox_6_T4), .Z0_f (new_AGEMA_signal_6535), .Z1_t (new_AGEMA_signal_6536), .Z1_f (new_AGEMA_signal_6537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[51]), .A0_f (ciphertext_s0_f[51]), .A1_t (ciphertext_s1_t[51]), .A1_f (ciphertext_s1_f[51]), .B0_t (ciphertext_s0_t[49]), .B0_f (ciphertext_s0_f[49]), .B1_t (ciphertext_s1_t[49]), .B1_f (ciphertext_s1_f[49]), .Z0_t (SubBytesIns_Inst_Sbox_6_T5), .Z0_f (new_AGEMA_signal_6538), .Z1_t (new_AGEMA_signal_6539), .Z1_f (new_AGEMA_signal_6540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T1), .A0_f (new_AGEMA_signal_6526), .A1_t (new_AGEMA_signal_6527), .A1_f (new_AGEMA_signal_6528), .B0_t (SubBytesIns_Inst_Sbox_6_T5), .B0_f (new_AGEMA_signal_6538), .B1_t (new_AGEMA_signal_6539), .B1_f (new_AGEMA_signal_6540), .Z0_t (SubBytesIns_Inst_Sbox_6_T6), .Z0_f (new_AGEMA_signal_7072), .Z1_t (new_AGEMA_signal_7073), .Z1_f (new_AGEMA_signal_7074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[54]), .A0_f (ciphertext_s0_f[54]), .A1_t (ciphertext_s1_t[54]), .A1_f (ciphertext_s1_f[54]), .B0_t (ciphertext_s0_t[53]), .B0_f (ciphertext_s0_f[53]), .B1_t (ciphertext_s1_t[53]), .B1_f (ciphertext_s1_f[53]), .Z0_t (SubBytesIns_Inst_Sbox_6_T7), .Z0_f (new_AGEMA_signal_6541), .Z1_t (new_AGEMA_signal_6542), .Z1_f (new_AGEMA_signal_6543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[48]), .A0_f (ciphertext_s0_f[48]), .A1_t (ciphertext_s1_t[48]), .A1_f (ciphertext_s1_f[48]), .B0_t (SubBytesIns_Inst_Sbox_6_T6), .B0_f (new_AGEMA_signal_7072), .B1_t (new_AGEMA_signal_7073), .B1_f (new_AGEMA_signal_7074), .Z0_t (SubBytesIns_Inst_Sbox_6_T8), .Z0_f (new_AGEMA_signal_7706), .Z1_t (new_AGEMA_signal_7707), .Z1_f (new_AGEMA_signal_7708) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[48]), .A0_f (ciphertext_s0_f[48]), .A1_t (ciphertext_s1_t[48]), .A1_f (ciphertext_s1_f[48]), .B0_t (SubBytesIns_Inst_Sbox_6_T7), .B0_f (new_AGEMA_signal_6541), .B1_t (new_AGEMA_signal_6542), .B1_f (new_AGEMA_signal_6543), .Z0_t (SubBytesIns_Inst_Sbox_6_T9), .Z0_f (new_AGEMA_signal_7075), .Z1_t (new_AGEMA_signal_7076), .Z1_f (new_AGEMA_signal_7077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T6), .A0_f (new_AGEMA_signal_7072), .A1_t (new_AGEMA_signal_7073), .A1_f (new_AGEMA_signal_7074), .B0_t (SubBytesIns_Inst_Sbox_6_T7), .B0_f (new_AGEMA_signal_6541), .B1_t (new_AGEMA_signal_6542), .B1_f (new_AGEMA_signal_6543), .Z0_t (SubBytesIns_Inst_Sbox_6_T10), .Z0_f (new_AGEMA_signal_7709), .Z1_t (new_AGEMA_signal_7710), .Z1_f (new_AGEMA_signal_7711) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[54]), .A0_f (ciphertext_s0_f[54]), .A1_t (ciphertext_s1_t[54]), .A1_f (ciphertext_s1_f[54]), .B0_t (ciphertext_s0_t[50]), .B0_f (ciphertext_s0_f[50]), .B1_t (ciphertext_s1_t[50]), .B1_f (ciphertext_s1_f[50]), .Z0_t (SubBytesIns_Inst_Sbox_6_T11), .Z0_f (new_AGEMA_signal_6544), .Z1_t (new_AGEMA_signal_6545), .Z1_f (new_AGEMA_signal_6546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[53]), .A0_f (ciphertext_s0_f[53]), .A1_t (ciphertext_s1_t[53]), .A1_f (ciphertext_s1_f[53]), .B0_t (ciphertext_s0_t[50]), .B0_f (ciphertext_s0_f[50]), .B1_t (ciphertext_s1_t[50]), .B1_f (ciphertext_s1_f[50]), .Z0_t (SubBytesIns_Inst_Sbox_6_T12), .Z0_f (new_AGEMA_signal_6547), .Z1_t (new_AGEMA_signal_6548), .Z1_f (new_AGEMA_signal_6549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T3), .A0_f (new_AGEMA_signal_6532), .A1_t (new_AGEMA_signal_6533), .A1_f (new_AGEMA_signal_6534), .B0_t (SubBytesIns_Inst_Sbox_6_T4), .B0_f (new_AGEMA_signal_6535), .B1_t (new_AGEMA_signal_6536), .B1_f (new_AGEMA_signal_6537), .Z0_t (SubBytesIns_Inst_Sbox_6_T13), .Z0_f (new_AGEMA_signal_7078), .Z1_t (new_AGEMA_signal_7079), .Z1_f (new_AGEMA_signal_7080) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T6), .A0_f (new_AGEMA_signal_7072), .A1_t (new_AGEMA_signal_7073), .A1_f (new_AGEMA_signal_7074), .B0_t (SubBytesIns_Inst_Sbox_6_T11), .B0_f (new_AGEMA_signal_6544), .B1_t (new_AGEMA_signal_6545), .B1_f (new_AGEMA_signal_6546), .Z0_t (SubBytesIns_Inst_Sbox_6_T14), .Z0_f (new_AGEMA_signal_7712), .Z1_t (new_AGEMA_signal_7713), .Z1_f (new_AGEMA_signal_7714) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T5), .A0_f (new_AGEMA_signal_6538), .A1_t (new_AGEMA_signal_6539), .A1_f (new_AGEMA_signal_6540), .B0_t (SubBytesIns_Inst_Sbox_6_T11), .B0_f (new_AGEMA_signal_6544), .B1_t (new_AGEMA_signal_6545), .B1_f (new_AGEMA_signal_6546), .Z0_t (SubBytesIns_Inst_Sbox_6_T15), .Z0_f (new_AGEMA_signal_7081), .Z1_t (new_AGEMA_signal_7082), .Z1_f (new_AGEMA_signal_7083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T5), .A0_f (new_AGEMA_signal_6538), .A1_t (new_AGEMA_signal_6539), .A1_f (new_AGEMA_signal_6540), .B0_t (SubBytesIns_Inst_Sbox_6_T12), .B0_f (new_AGEMA_signal_6547), .B1_t (new_AGEMA_signal_6548), .B1_f (new_AGEMA_signal_6549), .Z0_t (SubBytesIns_Inst_Sbox_6_T16), .Z0_f (new_AGEMA_signal_7084), .Z1_t (new_AGEMA_signal_7085), .Z1_f (new_AGEMA_signal_7086) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T9), .A0_f (new_AGEMA_signal_7075), .A1_t (new_AGEMA_signal_7076), .A1_f (new_AGEMA_signal_7077), .B0_t (SubBytesIns_Inst_Sbox_6_T16), .B0_f (new_AGEMA_signal_7084), .B1_t (new_AGEMA_signal_7085), .B1_f (new_AGEMA_signal_7086), .Z0_t (SubBytesIns_Inst_Sbox_6_T17), .Z0_f (new_AGEMA_signal_7715), .Z1_t (new_AGEMA_signal_7716), .Z1_f (new_AGEMA_signal_7717) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[52]), .A0_f (ciphertext_s0_f[52]), .A1_t (ciphertext_s1_t[52]), .A1_f (ciphertext_s1_f[52]), .B0_t (ciphertext_s0_t[48]), .B0_f (ciphertext_s0_f[48]), .B1_t (ciphertext_s1_t[48]), .B1_f (ciphertext_s1_f[48]), .Z0_t (SubBytesIns_Inst_Sbox_6_T18), .Z0_f (new_AGEMA_signal_6550), .Z1_t (new_AGEMA_signal_6551), .Z1_f (new_AGEMA_signal_6552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T7), .A0_f (new_AGEMA_signal_6541), .A1_t (new_AGEMA_signal_6542), .A1_f (new_AGEMA_signal_6543), .B0_t (SubBytesIns_Inst_Sbox_6_T18), .B0_f (new_AGEMA_signal_6550), .B1_t (new_AGEMA_signal_6551), .B1_f (new_AGEMA_signal_6552), .Z0_t (SubBytesIns_Inst_Sbox_6_T19), .Z0_f (new_AGEMA_signal_7087), .Z1_t (new_AGEMA_signal_7088), .Z1_f (new_AGEMA_signal_7089) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T1), .A0_f (new_AGEMA_signal_6526), .A1_t (new_AGEMA_signal_6527), .A1_f (new_AGEMA_signal_6528), .B0_t (SubBytesIns_Inst_Sbox_6_T19), .B0_f (new_AGEMA_signal_7087), .B1_t (new_AGEMA_signal_7088), .B1_f (new_AGEMA_signal_7089), .Z0_t (SubBytesIns_Inst_Sbox_6_T20), .Z0_f (new_AGEMA_signal_7718), .Z1_t (new_AGEMA_signal_7719), .Z1_f (new_AGEMA_signal_7720) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[49]), .A0_f (ciphertext_s0_f[49]), .A1_t (ciphertext_s1_t[49]), .A1_f (ciphertext_s1_f[49]), .B0_t (ciphertext_s0_t[48]), .B0_f (ciphertext_s0_f[48]), .B1_t (ciphertext_s1_t[48]), .B1_f (ciphertext_s1_f[48]), .Z0_t (SubBytesIns_Inst_Sbox_6_T21), .Z0_f (new_AGEMA_signal_6553), .Z1_t (new_AGEMA_signal_6554), .Z1_f (new_AGEMA_signal_6555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T7), .A0_f (new_AGEMA_signal_6541), .A1_t (new_AGEMA_signal_6542), .A1_f (new_AGEMA_signal_6543), .B0_t (SubBytesIns_Inst_Sbox_6_T21), .B0_f (new_AGEMA_signal_6553), .B1_t (new_AGEMA_signal_6554), .B1_f (new_AGEMA_signal_6555), .Z0_t (SubBytesIns_Inst_Sbox_6_T22), .Z0_f (new_AGEMA_signal_7090), .Z1_t (new_AGEMA_signal_7091), .Z1_f (new_AGEMA_signal_7092) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T2), .A0_f (new_AGEMA_signal_6529), .A1_t (new_AGEMA_signal_6530), .A1_f (new_AGEMA_signal_6531), .B0_t (SubBytesIns_Inst_Sbox_6_T22), .B0_f (new_AGEMA_signal_7090), .B1_t (new_AGEMA_signal_7091), .B1_f (new_AGEMA_signal_7092), .Z0_t (SubBytesIns_Inst_Sbox_6_T23), .Z0_f (new_AGEMA_signal_7721), .Z1_t (new_AGEMA_signal_7722), .Z1_f (new_AGEMA_signal_7723) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T2), .A0_f (new_AGEMA_signal_6529), .A1_t (new_AGEMA_signal_6530), .A1_f (new_AGEMA_signal_6531), .B0_t (SubBytesIns_Inst_Sbox_6_T10), .B0_f (new_AGEMA_signal_7709), .B1_t (new_AGEMA_signal_7710), .B1_f (new_AGEMA_signal_7711), .Z0_t (SubBytesIns_Inst_Sbox_6_T24), .Z0_f (new_AGEMA_signal_8366), .Z1_t (new_AGEMA_signal_8367), .Z1_f (new_AGEMA_signal_8368) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T20), .A0_f (new_AGEMA_signal_7718), .A1_t (new_AGEMA_signal_7719), .A1_f (new_AGEMA_signal_7720), .B0_t (SubBytesIns_Inst_Sbox_6_T17), .B0_f (new_AGEMA_signal_7715), .B1_t (new_AGEMA_signal_7716), .B1_f (new_AGEMA_signal_7717), .Z0_t (SubBytesIns_Inst_Sbox_6_T25), .Z0_f (new_AGEMA_signal_8369), .Z1_t (new_AGEMA_signal_8370), .Z1_f (new_AGEMA_signal_8371) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T3), .A0_f (new_AGEMA_signal_6532), .A1_t (new_AGEMA_signal_6533), .A1_f (new_AGEMA_signal_6534), .B0_t (SubBytesIns_Inst_Sbox_6_T16), .B0_f (new_AGEMA_signal_7084), .B1_t (new_AGEMA_signal_7085), .B1_f (new_AGEMA_signal_7086), .Z0_t (SubBytesIns_Inst_Sbox_6_T26), .Z0_f (new_AGEMA_signal_7724), .Z1_t (new_AGEMA_signal_7725), .Z1_f (new_AGEMA_signal_7726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T1), .A0_f (new_AGEMA_signal_6526), .A1_t (new_AGEMA_signal_6527), .A1_f (new_AGEMA_signal_6528), .B0_t (SubBytesIns_Inst_Sbox_6_T12), .B0_f (new_AGEMA_signal_6547), .B1_t (new_AGEMA_signal_6548), .B1_f (new_AGEMA_signal_6549), .Z0_t (SubBytesIns_Inst_Sbox_6_T27), .Z0_f (new_AGEMA_signal_7093), .Z1_t (new_AGEMA_signal_7094), .Z1_f (new_AGEMA_signal_7095) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T13), .A0_f (new_AGEMA_signal_7078), .A1_t (new_AGEMA_signal_7079), .A1_f (new_AGEMA_signal_7080), .B0_t (SubBytesIns_Inst_Sbox_6_T6), .B0_f (new_AGEMA_signal_7072), .B1_t (new_AGEMA_signal_7073), .B1_f (new_AGEMA_signal_7074), .Z0_t (SubBytesIns_Inst_Sbox_6_M1), .Z0_f (new_AGEMA_signal_7727), .Z1_t (new_AGEMA_signal_7728), .Z1_f (new_AGEMA_signal_7729) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T23), .A0_f (new_AGEMA_signal_7721), .A1_t (new_AGEMA_signal_7722), .A1_f (new_AGEMA_signal_7723), .B0_t (SubBytesIns_Inst_Sbox_6_T8), .B0_f (new_AGEMA_signal_7706), .B1_t (new_AGEMA_signal_7707), .B1_f (new_AGEMA_signal_7708), .Z0_t (SubBytesIns_Inst_Sbox_6_M2), .Z0_f (new_AGEMA_signal_8372), .Z1_t (new_AGEMA_signal_8373), .Z1_f (new_AGEMA_signal_8374) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T14), .A0_f (new_AGEMA_signal_7712), .A1_t (new_AGEMA_signal_7713), .A1_f (new_AGEMA_signal_7714), .B0_t (SubBytesIns_Inst_Sbox_6_M1), .B0_f (new_AGEMA_signal_7727), .B1_t (new_AGEMA_signal_7728), .B1_f (new_AGEMA_signal_7729), .Z0_t (SubBytesIns_Inst_Sbox_6_M3), .Z0_f (new_AGEMA_signal_8375), .Z1_t (new_AGEMA_signal_8376), .Z1_f (new_AGEMA_signal_8377) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T19), .A0_f (new_AGEMA_signal_7087), .A1_t (new_AGEMA_signal_7088), .A1_f (new_AGEMA_signal_7089), .B0_t (ciphertext_s0_t[48]), .B0_f (ciphertext_s0_f[48]), .B1_t (ciphertext_s1_t[48]), .B1_f (ciphertext_s1_f[48]), .Z0_t (SubBytesIns_Inst_Sbox_6_M4), .Z0_f (new_AGEMA_signal_7730), .Z1_t (new_AGEMA_signal_7731), .Z1_f (new_AGEMA_signal_7732) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M4), .A0_f (new_AGEMA_signal_7730), .A1_t (new_AGEMA_signal_7731), .A1_f (new_AGEMA_signal_7732), .B0_t (SubBytesIns_Inst_Sbox_6_M1), .B0_f (new_AGEMA_signal_7727), .B1_t (new_AGEMA_signal_7728), .B1_f (new_AGEMA_signal_7729), .Z0_t (SubBytesIns_Inst_Sbox_6_M5), .Z0_f (new_AGEMA_signal_8378), .Z1_t (new_AGEMA_signal_8379), .Z1_f (new_AGEMA_signal_8380) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T3), .A0_f (new_AGEMA_signal_6532), .A1_t (new_AGEMA_signal_6533), .A1_f (new_AGEMA_signal_6534), .B0_t (SubBytesIns_Inst_Sbox_6_T16), .B0_f (new_AGEMA_signal_7084), .B1_t (new_AGEMA_signal_7085), .B1_f (new_AGEMA_signal_7086), .Z0_t (SubBytesIns_Inst_Sbox_6_M6), .Z0_f (new_AGEMA_signal_7733), .Z1_t (new_AGEMA_signal_7734), .Z1_f (new_AGEMA_signal_7735) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T22), .A0_f (new_AGEMA_signal_7090), .A1_t (new_AGEMA_signal_7091), .A1_f (new_AGEMA_signal_7092), .B0_t (SubBytesIns_Inst_Sbox_6_T9), .B0_f (new_AGEMA_signal_7075), .B1_t (new_AGEMA_signal_7076), .B1_f (new_AGEMA_signal_7077), .Z0_t (SubBytesIns_Inst_Sbox_6_M7), .Z0_f (new_AGEMA_signal_7736), .Z1_t (new_AGEMA_signal_7737), .Z1_f (new_AGEMA_signal_7738) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T26), .A0_f (new_AGEMA_signal_7724), .A1_t (new_AGEMA_signal_7725), .A1_f (new_AGEMA_signal_7726), .B0_t (SubBytesIns_Inst_Sbox_6_M6), .B0_f (new_AGEMA_signal_7733), .B1_t (new_AGEMA_signal_7734), .B1_f (new_AGEMA_signal_7735), .Z0_t (SubBytesIns_Inst_Sbox_6_M8), .Z0_f (new_AGEMA_signal_8381), .Z1_t (new_AGEMA_signal_8382), .Z1_f (new_AGEMA_signal_8383) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T20), .A0_f (new_AGEMA_signal_7718), .A1_t (new_AGEMA_signal_7719), .A1_f (new_AGEMA_signal_7720), .B0_t (SubBytesIns_Inst_Sbox_6_T17), .B0_f (new_AGEMA_signal_7715), .B1_t (new_AGEMA_signal_7716), .B1_f (new_AGEMA_signal_7717), .Z0_t (SubBytesIns_Inst_Sbox_6_M9), .Z0_f (new_AGEMA_signal_8384), .Z1_t (new_AGEMA_signal_8385), .Z1_f (new_AGEMA_signal_8386) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M9), .A0_f (new_AGEMA_signal_8384), .A1_t (new_AGEMA_signal_8385), .A1_f (new_AGEMA_signal_8386), .B0_t (SubBytesIns_Inst_Sbox_6_M6), .B0_f (new_AGEMA_signal_7733), .B1_t (new_AGEMA_signal_7734), .B1_f (new_AGEMA_signal_7735), .Z0_t (SubBytesIns_Inst_Sbox_6_M10), .Z0_f (new_AGEMA_signal_8786), .Z1_t (new_AGEMA_signal_8787), .Z1_f (new_AGEMA_signal_8788) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T1), .A0_f (new_AGEMA_signal_6526), .A1_t (new_AGEMA_signal_6527), .A1_f (new_AGEMA_signal_6528), .B0_t (SubBytesIns_Inst_Sbox_6_T15), .B0_f (new_AGEMA_signal_7081), .B1_t (new_AGEMA_signal_7082), .B1_f (new_AGEMA_signal_7083), .Z0_t (SubBytesIns_Inst_Sbox_6_M11), .Z0_f (new_AGEMA_signal_7739), .Z1_t (new_AGEMA_signal_7740), .Z1_f (new_AGEMA_signal_7741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T4), .A0_f (new_AGEMA_signal_6535), .A1_t (new_AGEMA_signal_6536), .A1_f (new_AGEMA_signal_6537), .B0_t (SubBytesIns_Inst_Sbox_6_T27), .B0_f (new_AGEMA_signal_7093), .B1_t (new_AGEMA_signal_7094), .B1_f (new_AGEMA_signal_7095), .Z0_t (SubBytesIns_Inst_Sbox_6_M12), .Z0_f (new_AGEMA_signal_7742), .Z1_t (new_AGEMA_signal_7743), .Z1_f (new_AGEMA_signal_7744) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M12), .A0_f (new_AGEMA_signal_7742), .A1_t (new_AGEMA_signal_7743), .A1_f (new_AGEMA_signal_7744), .B0_t (SubBytesIns_Inst_Sbox_6_M11), .B0_f (new_AGEMA_signal_7739), .B1_t (new_AGEMA_signal_7740), .B1_f (new_AGEMA_signal_7741), .Z0_t (SubBytesIns_Inst_Sbox_6_M13), .Z0_f (new_AGEMA_signal_8387), .Z1_t (new_AGEMA_signal_8388), .Z1_f (new_AGEMA_signal_8389) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T2), .A0_f (new_AGEMA_signal_6529), .A1_t (new_AGEMA_signal_6530), .A1_f (new_AGEMA_signal_6531), .B0_t (SubBytesIns_Inst_Sbox_6_T10), .B0_f (new_AGEMA_signal_7709), .B1_t (new_AGEMA_signal_7710), .B1_f (new_AGEMA_signal_7711), .Z0_t (SubBytesIns_Inst_Sbox_6_M14), .Z0_f (new_AGEMA_signal_8390), .Z1_t (new_AGEMA_signal_8391), .Z1_f (new_AGEMA_signal_8392) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M14), .A0_f (new_AGEMA_signal_8390), .A1_t (new_AGEMA_signal_8391), .A1_f (new_AGEMA_signal_8392), .B0_t (SubBytesIns_Inst_Sbox_6_M11), .B0_f (new_AGEMA_signal_7739), .B1_t (new_AGEMA_signal_7740), .B1_f (new_AGEMA_signal_7741), .Z0_t (SubBytesIns_Inst_Sbox_6_M15), .Z0_f (new_AGEMA_signal_8789), .Z1_t (new_AGEMA_signal_8790), .Z1_f (new_AGEMA_signal_8791) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M3), .A0_f (new_AGEMA_signal_8375), .A1_t (new_AGEMA_signal_8376), .A1_f (new_AGEMA_signal_8377), .B0_t (SubBytesIns_Inst_Sbox_6_M2), .B0_f (new_AGEMA_signal_8372), .B1_t (new_AGEMA_signal_8373), .B1_f (new_AGEMA_signal_8374), .Z0_t (SubBytesIns_Inst_Sbox_6_M16), .Z0_f (new_AGEMA_signal_8792), .Z1_t (new_AGEMA_signal_8793), .Z1_f (new_AGEMA_signal_8794) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M5), .A0_f (new_AGEMA_signal_8378), .A1_t (new_AGEMA_signal_8379), .A1_f (new_AGEMA_signal_8380), .B0_t (SubBytesIns_Inst_Sbox_6_T24), .B0_f (new_AGEMA_signal_8366), .B1_t (new_AGEMA_signal_8367), .B1_f (new_AGEMA_signal_8368), .Z0_t (SubBytesIns_Inst_Sbox_6_M17), .Z0_f (new_AGEMA_signal_8795), .Z1_t (new_AGEMA_signal_8796), .Z1_f (new_AGEMA_signal_8797) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M8), .A0_f (new_AGEMA_signal_8381), .A1_t (new_AGEMA_signal_8382), .A1_f (new_AGEMA_signal_8383), .B0_t (SubBytesIns_Inst_Sbox_6_M7), .B0_f (new_AGEMA_signal_7736), .B1_t (new_AGEMA_signal_7737), .B1_f (new_AGEMA_signal_7738), .Z0_t (SubBytesIns_Inst_Sbox_6_M18), .Z0_f (new_AGEMA_signal_8798), .Z1_t (new_AGEMA_signal_8799), .Z1_f (new_AGEMA_signal_8800) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M10), .A0_f (new_AGEMA_signal_8786), .A1_t (new_AGEMA_signal_8787), .A1_f (new_AGEMA_signal_8788), .B0_t (SubBytesIns_Inst_Sbox_6_M15), .B0_f (new_AGEMA_signal_8789), .B1_t (new_AGEMA_signal_8790), .B1_f (new_AGEMA_signal_8791), .Z0_t (SubBytesIns_Inst_Sbox_6_M19), .Z0_f (new_AGEMA_signal_9056), .Z1_t (new_AGEMA_signal_9057), .Z1_f (new_AGEMA_signal_9058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M16), .A0_f (new_AGEMA_signal_8792), .A1_t (new_AGEMA_signal_8793), .A1_f (new_AGEMA_signal_8794), .B0_t (SubBytesIns_Inst_Sbox_6_M13), .B0_f (new_AGEMA_signal_8387), .B1_t (new_AGEMA_signal_8388), .B1_f (new_AGEMA_signal_8389), .Z0_t (SubBytesIns_Inst_Sbox_6_M20), .Z0_f (new_AGEMA_signal_9059), .Z1_t (new_AGEMA_signal_9060), .Z1_f (new_AGEMA_signal_9061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M17), .A0_f (new_AGEMA_signal_8795), .A1_t (new_AGEMA_signal_8796), .A1_f (new_AGEMA_signal_8797), .B0_t (SubBytesIns_Inst_Sbox_6_M15), .B0_f (new_AGEMA_signal_8789), .B1_t (new_AGEMA_signal_8790), .B1_f (new_AGEMA_signal_8791), .Z0_t (SubBytesIns_Inst_Sbox_6_M21), .Z0_f (new_AGEMA_signal_9062), .Z1_t (new_AGEMA_signal_9063), .Z1_f (new_AGEMA_signal_9064) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M18), .A0_f (new_AGEMA_signal_8798), .A1_t (new_AGEMA_signal_8799), .A1_f (new_AGEMA_signal_8800), .B0_t (SubBytesIns_Inst_Sbox_6_M13), .B0_f (new_AGEMA_signal_8387), .B1_t (new_AGEMA_signal_8388), .B1_f (new_AGEMA_signal_8389), .Z0_t (SubBytesIns_Inst_Sbox_6_M22), .Z0_f (new_AGEMA_signal_9065), .Z1_t (new_AGEMA_signal_9066), .Z1_f (new_AGEMA_signal_9067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M19), .A0_f (new_AGEMA_signal_9056), .A1_t (new_AGEMA_signal_9057), .A1_f (new_AGEMA_signal_9058), .B0_t (SubBytesIns_Inst_Sbox_6_T25), .B0_f (new_AGEMA_signal_8369), .B1_t (new_AGEMA_signal_8370), .B1_f (new_AGEMA_signal_8371), .Z0_t (SubBytesIns_Inst_Sbox_6_M23), .Z0_f (new_AGEMA_signal_9296), .Z1_t (new_AGEMA_signal_9297), .Z1_f (new_AGEMA_signal_9298) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M22), .A0_f (new_AGEMA_signal_9065), .A1_t (new_AGEMA_signal_9066), .A1_f (new_AGEMA_signal_9067), .B0_t (SubBytesIns_Inst_Sbox_6_M23), .B0_f (new_AGEMA_signal_9296), .B1_t (new_AGEMA_signal_9297), .B1_f (new_AGEMA_signal_9298), .Z0_t (SubBytesIns_Inst_Sbox_6_M24), .Z0_f (new_AGEMA_signal_9566), .Z1_t (new_AGEMA_signal_9567), .Z1_f (new_AGEMA_signal_9568) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M22), .A0_f (new_AGEMA_signal_9065), .A1_t (new_AGEMA_signal_9066), .A1_f (new_AGEMA_signal_9067), .B0_t (SubBytesIns_Inst_Sbox_6_M20), .B0_f (new_AGEMA_signal_9059), .B1_t (new_AGEMA_signal_9060), .B1_f (new_AGEMA_signal_9061), .Z0_t (SubBytesIns_Inst_Sbox_6_M25), .Z0_f (new_AGEMA_signal_9299), .Z1_t (new_AGEMA_signal_9300), .Z1_f (new_AGEMA_signal_9301) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M21), .A0_f (new_AGEMA_signal_9062), .A1_t (new_AGEMA_signal_9063), .A1_f (new_AGEMA_signal_9064), .B0_t (SubBytesIns_Inst_Sbox_6_M25), .B0_f (new_AGEMA_signal_9299), .B1_t (new_AGEMA_signal_9300), .B1_f (new_AGEMA_signal_9301), .Z0_t (SubBytesIns_Inst_Sbox_6_M26), .Z0_f (new_AGEMA_signal_9569), .Z1_t (new_AGEMA_signal_9570), .Z1_f (new_AGEMA_signal_9571) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M20), .A0_f (new_AGEMA_signal_9059), .A1_t (new_AGEMA_signal_9060), .A1_f (new_AGEMA_signal_9061), .B0_t (SubBytesIns_Inst_Sbox_6_M21), .B0_f (new_AGEMA_signal_9062), .B1_t (new_AGEMA_signal_9063), .B1_f (new_AGEMA_signal_9064), .Z0_t (SubBytesIns_Inst_Sbox_6_M27), .Z0_f (new_AGEMA_signal_9302), .Z1_t (new_AGEMA_signal_9303), .Z1_f (new_AGEMA_signal_9304) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M23), .A0_f (new_AGEMA_signal_9296), .A1_t (new_AGEMA_signal_9297), .A1_f (new_AGEMA_signal_9298), .B0_t (SubBytesIns_Inst_Sbox_6_M25), .B0_f (new_AGEMA_signal_9299), .B1_t (new_AGEMA_signal_9300), .B1_f (new_AGEMA_signal_9301), .Z0_t (SubBytesIns_Inst_Sbox_6_M28), .Z0_f (new_AGEMA_signal_9572), .Z1_t (new_AGEMA_signal_9573), .Z1_f (new_AGEMA_signal_9574) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M28), .A0_f (new_AGEMA_signal_9572), .A1_t (new_AGEMA_signal_9573), .A1_f (new_AGEMA_signal_9574), .B0_t (SubBytesIns_Inst_Sbox_6_M27), .B0_f (new_AGEMA_signal_9302), .B1_t (new_AGEMA_signal_9303), .B1_f (new_AGEMA_signal_9304), .Z0_t (SubBytesIns_Inst_Sbox_6_M29), .Z0_f (new_AGEMA_signal_9866), .Z1_t (new_AGEMA_signal_9867), .Z1_f (new_AGEMA_signal_9868) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M26), .A0_f (new_AGEMA_signal_9569), .A1_t (new_AGEMA_signal_9570), .A1_f (new_AGEMA_signal_9571), .B0_t (SubBytesIns_Inst_Sbox_6_M24), .B0_f (new_AGEMA_signal_9566), .B1_t (new_AGEMA_signal_9567), .B1_f (new_AGEMA_signal_9568), .Z0_t (SubBytesIns_Inst_Sbox_6_M30), .Z0_f (new_AGEMA_signal_9869), .Z1_t (new_AGEMA_signal_9870), .Z1_f (new_AGEMA_signal_9871) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M20), .A0_f (new_AGEMA_signal_9059), .A1_t (new_AGEMA_signal_9060), .A1_f (new_AGEMA_signal_9061), .B0_t (SubBytesIns_Inst_Sbox_6_M23), .B0_f (new_AGEMA_signal_9296), .B1_t (new_AGEMA_signal_9297), .B1_f (new_AGEMA_signal_9298), .Z0_t (SubBytesIns_Inst_Sbox_6_M31), .Z0_f (new_AGEMA_signal_9575), .Z1_t (new_AGEMA_signal_9576), .Z1_f (new_AGEMA_signal_9577) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M27), .A0_f (new_AGEMA_signal_9302), .A1_t (new_AGEMA_signal_9303), .A1_f (new_AGEMA_signal_9304), .B0_t (SubBytesIns_Inst_Sbox_6_M31), .B0_f (new_AGEMA_signal_9575), .B1_t (new_AGEMA_signal_9576), .B1_f (new_AGEMA_signal_9577), .Z0_t (SubBytesIns_Inst_Sbox_6_M32), .Z0_f (new_AGEMA_signal_9872), .Z1_t (new_AGEMA_signal_9873), .Z1_f (new_AGEMA_signal_9874) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M27), .A0_f (new_AGEMA_signal_9302), .A1_t (new_AGEMA_signal_9303), .A1_f (new_AGEMA_signal_9304), .B0_t (SubBytesIns_Inst_Sbox_6_M25), .B0_f (new_AGEMA_signal_9299), .B1_t (new_AGEMA_signal_9300), .B1_f (new_AGEMA_signal_9301), .Z0_t (SubBytesIns_Inst_Sbox_6_M33), .Z0_f (new_AGEMA_signal_9578), .Z1_t (new_AGEMA_signal_9579), .Z1_f (new_AGEMA_signal_9580) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M21), .A0_f (new_AGEMA_signal_9062), .A1_t (new_AGEMA_signal_9063), .A1_f (new_AGEMA_signal_9064), .B0_t (SubBytesIns_Inst_Sbox_6_M22), .B0_f (new_AGEMA_signal_9065), .B1_t (new_AGEMA_signal_9066), .B1_f (new_AGEMA_signal_9067), .Z0_t (SubBytesIns_Inst_Sbox_6_M34), .Z0_f (new_AGEMA_signal_9305), .Z1_t (new_AGEMA_signal_9306), .Z1_f (new_AGEMA_signal_9307) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M24), .A0_f (new_AGEMA_signal_9566), .A1_t (new_AGEMA_signal_9567), .A1_f (new_AGEMA_signal_9568), .B0_t (SubBytesIns_Inst_Sbox_6_M34), .B0_f (new_AGEMA_signal_9305), .B1_t (new_AGEMA_signal_9306), .B1_f (new_AGEMA_signal_9307), .Z0_t (SubBytesIns_Inst_Sbox_6_M35), .Z0_f (new_AGEMA_signal_9875), .Z1_t (new_AGEMA_signal_9876), .Z1_f (new_AGEMA_signal_9877) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M24), .A0_f (new_AGEMA_signal_9566), .A1_t (new_AGEMA_signal_9567), .A1_f (new_AGEMA_signal_9568), .B0_t (SubBytesIns_Inst_Sbox_6_M25), .B0_f (new_AGEMA_signal_9299), .B1_t (new_AGEMA_signal_9300), .B1_f (new_AGEMA_signal_9301), .Z0_t (SubBytesIns_Inst_Sbox_6_M36), .Z0_f (new_AGEMA_signal_9878), .Z1_t (new_AGEMA_signal_9879), .Z1_f (new_AGEMA_signal_9880) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M21), .A0_f (new_AGEMA_signal_9062), .A1_t (new_AGEMA_signal_9063), .A1_f (new_AGEMA_signal_9064), .B0_t (SubBytesIns_Inst_Sbox_6_M29), .B0_f (new_AGEMA_signal_9866), .B1_t (new_AGEMA_signal_9867), .B1_f (new_AGEMA_signal_9868), .Z0_t (SubBytesIns_Inst_Sbox_6_M37), .Z0_f (new_AGEMA_signal_10136), .Z1_t (new_AGEMA_signal_10137), .Z1_f (new_AGEMA_signal_10138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M32), .A0_f (new_AGEMA_signal_9872), .A1_t (new_AGEMA_signal_9873), .A1_f (new_AGEMA_signal_9874), .B0_t (SubBytesIns_Inst_Sbox_6_M33), .B0_f (new_AGEMA_signal_9578), .B1_t (new_AGEMA_signal_9579), .B1_f (new_AGEMA_signal_9580), .Z0_t (SubBytesIns_Inst_Sbox_6_M38), .Z0_f (new_AGEMA_signal_10139), .Z1_t (new_AGEMA_signal_10140), .Z1_f (new_AGEMA_signal_10141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M23), .A0_f (new_AGEMA_signal_9296), .A1_t (new_AGEMA_signal_9297), .A1_f (new_AGEMA_signal_9298), .B0_t (SubBytesIns_Inst_Sbox_6_M30), .B0_f (new_AGEMA_signal_9869), .B1_t (new_AGEMA_signal_9870), .B1_f (new_AGEMA_signal_9871), .Z0_t (SubBytesIns_Inst_Sbox_6_M39), .Z0_f (new_AGEMA_signal_10142), .Z1_t (new_AGEMA_signal_10143), .Z1_f (new_AGEMA_signal_10144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M35), .A0_f (new_AGEMA_signal_9875), .A1_t (new_AGEMA_signal_9876), .A1_f (new_AGEMA_signal_9877), .B0_t (SubBytesIns_Inst_Sbox_6_M36), .B0_f (new_AGEMA_signal_9878), .B1_t (new_AGEMA_signal_9879), .B1_f (new_AGEMA_signal_9880), .Z0_t (SubBytesIns_Inst_Sbox_6_M40), .Z0_f (new_AGEMA_signal_10145), .Z1_t (new_AGEMA_signal_10146), .Z1_f (new_AGEMA_signal_10147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M38), .A0_f (new_AGEMA_signal_10139), .A1_t (new_AGEMA_signal_10140), .A1_f (new_AGEMA_signal_10141), .B0_t (SubBytesIns_Inst_Sbox_6_M40), .B0_f (new_AGEMA_signal_10145), .B1_t (new_AGEMA_signal_10146), .B1_f (new_AGEMA_signal_10147), .Z0_t (SubBytesIns_Inst_Sbox_6_M41), .Z0_f (new_AGEMA_signal_10616), .Z1_t (new_AGEMA_signal_10617), .Z1_f (new_AGEMA_signal_10618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M37), .A0_f (new_AGEMA_signal_10136), .A1_t (new_AGEMA_signal_10137), .A1_f (new_AGEMA_signal_10138), .B0_t (SubBytesIns_Inst_Sbox_6_M39), .B0_f (new_AGEMA_signal_10142), .B1_t (new_AGEMA_signal_10143), .B1_f (new_AGEMA_signal_10144), .Z0_t (SubBytesIns_Inst_Sbox_6_M42), .Z0_f (new_AGEMA_signal_10619), .Z1_t (new_AGEMA_signal_10620), .Z1_f (new_AGEMA_signal_10621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M37), .A0_f (new_AGEMA_signal_10136), .A1_t (new_AGEMA_signal_10137), .A1_f (new_AGEMA_signal_10138), .B0_t (SubBytesIns_Inst_Sbox_6_M38), .B0_f (new_AGEMA_signal_10139), .B1_t (new_AGEMA_signal_10140), .B1_f (new_AGEMA_signal_10141), .Z0_t (SubBytesIns_Inst_Sbox_6_M43), .Z0_f (new_AGEMA_signal_10622), .Z1_t (new_AGEMA_signal_10623), .Z1_f (new_AGEMA_signal_10624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M39), .A0_f (new_AGEMA_signal_10142), .A1_t (new_AGEMA_signal_10143), .A1_f (new_AGEMA_signal_10144), .B0_t (SubBytesIns_Inst_Sbox_6_M40), .B0_f (new_AGEMA_signal_10145), .B1_t (new_AGEMA_signal_10146), .B1_f (new_AGEMA_signal_10147), .Z0_t (SubBytesIns_Inst_Sbox_6_M44), .Z0_f (new_AGEMA_signal_10625), .Z1_t (new_AGEMA_signal_10626), .Z1_f (new_AGEMA_signal_10627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M42), .A0_f (new_AGEMA_signal_10619), .A1_t (new_AGEMA_signal_10620), .A1_f (new_AGEMA_signal_10621), .B0_t (SubBytesIns_Inst_Sbox_6_M41), .B0_f (new_AGEMA_signal_10616), .B1_t (new_AGEMA_signal_10617), .B1_f (new_AGEMA_signal_10618), .Z0_t (SubBytesIns_Inst_Sbox_6_M45), .Z0_f (new_AGEMA_signal_11336), .Z1_t (new_AGEMA_signal_11337), .Z1_f (new_AGEMA_signal_11338) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M44), .A0_f (new_AGEMA_signal_10625), .A1_t (new_AGEMA_signal_10626), .A1_f (new_AGEMA_signal_10627), .B0_t (SubBytesIns_Inst_Sbox_6_T6), .B0_f (new_AGEMA_signal_7072), .B1_t (new_AGEMA_signal_7073), .B1_f (new_AGEMA_signal_7074), .Z0_t (SubBytesIns_Inst_Sbox_6_M46), .Z0_f (new_AGEMA_signal_11339), .Z1_t (new_AGEMA_signal_11340), .Z1_f (new_AGEMA_signal_11341) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M40), .A0_f (new_AGEMA_signal_10145), .A1_t (new_AGEMA_signal_10146), .A1_f (new_AGEMA_signal_10147), .B0_t (SubBytesIns_Inst_Sbox_6_T8), .B0_f (new_AGEMA_signal_7706), .B1_t (new_AGEMA_signal_7707), .B1_f (new_AGEMA_signal_7708), .Z0_t (SubBytesIns_Inst_Sbox_6_M47), .Z0_f (new_AGEMA_signal_10628), .Z1_t (new_AGEMA_signal_10629), .Z1_f (new_AGEMA_signal_10630) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M39), .A0_f (new_AGEMA_signal_10142), .A1_t (new_AGEMA_signal_10143), .A1_f (new_AGEMA_signal_10144), .B0_t (ciphertext_s0_t[48]), .B0_f (ciphertext_s0_f[48]), .B1_t (ciphertext_s1_t[48]), .B1_f (ciphertext_s1_f[48]), .Z0_t (SubBytesIns_Inst_Sbox_6_M48), .Z0_f (new_AGEMA_signal_10631), .Z1_t (new_AGEMA_signal_10632), .Z1_f (new_AGEMA_signal_10633) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M43), .A0_f (new_AGEMA_signal_10622), .A1_t (new_AGEMA_signal_10623), .A1_f (new_AGEMA_signal_10624), .B0_t (SubBytesIns_Inst_Sbox_6_T16), .B0_f (new_AGEMA_signal_7084), .B1_t (new_AGEMA_signal_7085), .B1_f (new_AGEMA_signal_7086), .Z0_t (SubBytesIns_Inst_Sbox_6_M49), .Z0_f (new_AGEMA_signal_11342), .Z1_t (new_AGEMA_signal_11343), .Z1_f (new_AGEMA_signal_11344) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M38), .A0_f (new_AGEMA_signal_10139), .A1_t (new_AGEMA_signal_10140), .A1_f (new_AGEMA_signal_10141), .B0_t (SubBytesIns_Inst_Sbox_6_T9), .B0_f (new_AGEMA_signal_7075), .B1_t (new_AGEMA_signal_7076), .B1_f (new_AGEMA_signal_7077), .Z0_t (SubBytesIns_Inst_Sbox_6_M50), .Z0_f (new_AGEMA_signal_10634), .Z1_t (new_AGEMA_signal_10635), .Z1_f (new_AGEMA_signal_10636) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M37), .A0_f (new_AGEMA_signal_10136), .A1_t (new_AGEMA_signal_10137), .A1_f (new_AGEMA_signal_10138), .B0_t (SubBytesIns_Inst_Sbox_6_T17), .B0_f (new_AGEMA_signal_7715), .B1_t (new_AGEMA_signal_7716), .B1_f (new_AGEMA_signal_7717), .Z0_t (SubBytesIns_Inst_Sbox_6_M51), .Z0_f (new_AGEMA_signal_10637), .Z1_t (new_AGEMA_signal_10638), .Z1_f (new_AGEMA_signal_10639) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M42), .A0_f (new_AGEMA_signal_10619), .A1_t (new_AGEMA_signal_10620), .A1_f (new_AGEMA_signal_10621), .B0_t (SubBytesIns_Inst_Sbox_6_T15), .B0_f (new_AGEMA_signal_7081), .B1_t (new_AGEMA_signal_7082), .B1_f (new_AGEMA_signal_7083), .Z0_t (SubBytesIns_Inst_Sbox_6_M52), .Z0_f (new_AGEMA_signal_11345), .Z1_t (new_AGEMA_signal_11346), .Z1_f (new_AGEMA_signal_11347) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M45), .A0_f (new_AGEMA_signal_11336), .A1_t (new_AGEMA_signal_11337), .A1_f (new_AGEMA_signal_11338), .B0_t (SubBytesIns_Inst_Sbox_6_T27), .B0_f (new_AGEMA_signal_7093), .B1_t (new_AGEMA_signal_7094), .B1_f (new_AGEMA_signal_7095), .Z0_t (SubBytesIns_Inst_Sbox_6_M53), .Z0_f (new_AGEMA_signal_11996), .Z1_t (new_AGEMA_signal_11997), .Z1_f (new_AGEMA_signal_11998) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M41), .A0_f (new_AGEMA_signal_10616), .A1_t (new_AGEMA_signal_10617), .A1_f (new_AGEMA_signal_10618), .B0_t (SubBytesIns_Inst_Sbox_6_T10), .B0_f (new_AGEMA_signal_7709), .B1_t (new_AGEMA_signal_7710), .B1_f (new_AGEMA_signal_7711), .Z0_t (SubBytesIns_Inst_Sbox_6_M54), .Z0_f (new_AGEMA_signal_11348), .Z1_t (new_AGEMA_signal_11349), .Z1_f (new_AGEMA_signal_11350) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M44), .A0_f (new_AGEMA_signal_10625), .A1_t (new_AGEMA_signal_10626), .A1_f (new_AGEMA_signal_10627), .B0_t (SubBytesIns_Inst_Sbox_6_T13), .B0_f (new_AGEMA_signal_7078), .B1_t (new_AGEMA_signal_7079), .B1_f (new_AGEMA_signal_7080), .Z0_t (SubBytesIns_Inst_Sbox_6_M55), .Z0_f (new_AGEMA_signal_11351), .Z1_t (new_AGEMA_signal_11352), .Z1_f (new_AGEMA_signal_11353) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M40), .A0_f (new_AGEMA_signal_10145), .A1_t (new_AGEMA_signal_10146), .A1_f (new_AGEMA_signal_10147), .B0_t (SubBytesIns_Inst_Sbox_6_T23), .B0_f (new_AGEMA_signal_7721), .B1_t (new_AGEMA_signal_7722), .B1_f (new_AGEMA_signal_7723), .Z0_t (SubBytesIns_Inst_Sbox_6_M56), .Z0_f (new_AGEMA_signal_10640), .Z1_t (new_AGEMA_signal_10641), .Z1_f (new_AGEMA_signal_10642) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M39), .A0_f (new_AGEMA_signal_10142), .A1_t (new_AGEMA_signal_10143), .A1_f (new_AGEMA_signal_10144), .B0_t (SubBytesIns_Inst_Sbox_6_T19), .B0_f (new_AGEMA_signal_7087), .B1_t (new_AGEMA_signal_7088), .B1_f (new_AGEMA_signal_7089), .Z0_t (SubBytesIns_Inst_Sbox_6_M57), .Z0_f (new_AGEMA_signal_10643), .Z1_t (new_AGEMA_signal_10644), .Z1_f (new_AGEMA_signal_10645) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M43), .A0_f (new_AGEMA_signal_10622), .A1_t (new_AGEMA_signal_10623), .A1_f (new_AGEMA_signal_10624), .B0_t (SubBytesIns_Inst_Sbox_6_T3), .B0_f (new_AGEMA_signal_6532), .B1_t (new_AGEMA_signal_6533), .B1_f (new_AGEMA_signal_6534), .Z0_t (SubBytesIns_Inst_Sbox_6_M58), .Z0_f (new_AGEMA_signal_11354), .Z1_t (new_AGEMA_signal_11355), .Z1_f (new_AGEMA_signal_11356) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M38), .A0_f (new_AGEMA_signal_10139), .A1_t (new_AGEMA_signal_10140), .A1_f (new_AGEMA_signal_10141), .B0_t (SubBytesIns_Inst_Sbox_6_T22), .B0_f (new_AGEMA_signal_7090), .B1_t (new_AGEMA_signal_7091), .B1_f (new_AGEMA_signal_7092), .Z0_t (SubBytesIns_Inst_Sbox_6_M59), .Z0_f (new_AGEMA_signal_10646), .Z1_t (new_AGEMA_signal_10647), .Z1_f (new_AGEMA_signal_10648) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M37), .A0_f (new_AGEMA_signal_10136), .A1_t (new_AGEMA_signal_10137), .A1_f (new_AGEMA_signal_10138), .B0_t (SubBytesIns_Inst_Sbox_6_T20), .B0_f (new_AGEMA_signal_7718), .B1_t (new_AGEMA_signal_7719), .B1_f (new_AGEMA_signal_7720), .Z0_t (SubBytesIns_Inst_Sbox_6_M60), .Z0_f (new_AGEMA_signal_10649), .Z1_t (new_AGEMA_signal_10650), .Z1_f (new_AGEMA_signal_10651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M42), .A0_f (new_AGEMA_signal_10619), .A1_t (new_AGEMA_signal_10620), .A1_f (new_AGEMA_signal_10621), .B0_t (SubBytesIns_Inst_Sbox_6_T1), .B0_f (new_AGEMA_signal_6526), .B1_t (new_AGEMA_signal_6527), .B1_f (new_AGEMA_signal_6528), .Z0_t (SubBytesIns_Inst_Sbox_6_M61), .Z0_f (new_AGEMA_signal_11357), .Z1_t (new_AGEMA_signal_11358), .Z1_f (new_AGEMA_signal_11359) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M45), .A0_f (new_AGEMA_signal_11336), .A1_t (new_AGEMA_signal_11337), .A1_f (new_AGEMA_signal_11338), .B0_t (SubBytesIns_Inst_Sbox_6_T4), .B0_f (new_AGEMA_signal_6535), .B1_t (new_AGEMA_signal_6536), .B1_f (new_AGEMA_signal_6537), .Z0_t (SubBytesIns_Inst_Sbox_6_M62), .Z0_f (new_AGEMA_signal_11999), .Z1_t (new_AGEMA_signal_12000), .Z1_f (new_AGEMA_signal_12001) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M41), .A0_f (new_AGEMA_signal_10616), .A1_t (new_AGEMA_signal_10617), .A1_f (new_AGEMA_signal_10618), .B0_t (SubBytesIns_Inst_Sbox_6_T2), .B0_f (new_AGEMA_signal_6529), .B1_t (new_AGEMA_signal_6530), .B1_f (new_AGEMA_signal_6531), .Z0_t (SubBytesIns_Inst_Sbox_6_M63), .Z0_f (new_AGEMA_signal_11360), .Z1_t (new_AGEMA_signal_11361), .Z1_f (new_AGEMA_signal_11362) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M61), .A0_f (new_AGEMA_signal_11357), .A1_t (new_AGEMA_signal_11358), .A1_f (new_AGEMA_signal_11359), .B0_t (SubBytesIns_Inst_Sbox_6_M62), .B0_f (new_AGEMA_signal_11999), .B1_t (new_AGEMA_signal_12000), .B1_f (new_AGEMA_signal_12001), .Z0_t (SubBytesIns_Inst_Sbox_6_L0), .Z0_f (new_AGEMA_signal_12566), .Z1_t (new_AGEMA_signal_12567), .Z1_f (new_AGEMA_signal_12568) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M50), .A0_f (new_AGEMA_signal_10634), .A1_t (new_AGEMA_signal_10635), .A1_f (new_AGEMA_signal_10636), .B0_t (SubBytesIns_Inst_Sbox_6_M56), .B0_f (new_AGEMA_signal_10640), .B1_t (new_AGEMA_signal_10641), .B1_f (new_AGEMA_signal_10642), .Z0_t (SubBytesIns_Inst_Sbox_6_L1), .Z0_f (new_AGEMA_signal_11363), .Z1_t (new_AGEMA_signal_11364), .Z1_f (new_AGEMA_signal_11365) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M46), .A0_f (new_AGEMA_signal_11339), .A1_t (new_AGEMA_signal_11340), .A1_f (new_AGEMA_signal_11341), .B0_t (SubBytesIns_Inst_Sbox_6_M48), .B0_f (new_AGEMA_signal_10631), .B1_t (new_AGEMA_signal_10632), .B1_f (new_AGEMA_signal_10633), .Z0_t (SubBytesIns_Inst_Sbox_6_L2), .Z0_f (new_AGEMA_signal_12002), .Z1_t (new_AGEMA_signal_12003), .Z1_f (new_AGEMA_signal_12004) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M47), .A0_f (new_AGEMA_signal_10628), .A1_t (new_AGEMA_signal_10629), .A1_f (new_AGEMA_signal_10630), .B0_t (SubBytesIns_Inst_Sbox_6_M55), .B0_f (new_AGEMA_signal_11351), .B1_t (new_AGEMA_signal_11352), .B1_f (new_AGEMA_signal_11353), .Z0_t (SubBytesIns_Inst_Sbox_6_L3), .Z0_f (new_AGEMA_signal_12005), .Z1_t (new_AGEMA_signal_12006), .Z1_f (new_AGEMA_signal_12007) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M54), .A0_f (new_AGEMA_signal_11348), .A1_t (new_AGEMA_signal_11349), .A1_f (new_AGEMA_signal_11350), .B0_t (SubBytesIns_Inst_Sbox_6_M58), .B0_f (new_AGEMA_signal_11354), .B1_t (new_AGEMA_signal_11355), .B1_f (new_AGEMA_signal_11356), .Z0_t (SubBytesIns_Inst_Sbox_6_L4), .Z0_f (new_AGEMA_signal_12008), .Z1_t (new_AGEMA_signal_12009), .Z1_f (new_AGEMA_signal_12010) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M49), .A0_f (new_AGEMA_signal_11342), .A1_t (new_AGEMA_signal_11343), .A1_f (new_AGEMA_signal_11344), .B0_t (SubBytesIns_Inst_Sbox_6_M61), .B0_f (new_AGEMA_signal_11357), .B1_t (new_AGEMA_signal_11358), .B1_f (new_AGEMA_signal_11359), .Z0_t (SubBytesIns_Inst_Sbox_6_L5), .Z0_f (new_AGEMA_signal_12011), .Z1_t (new_AGEMA_signal_12012), .Z1_f (new_AGEMA_signal_12013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M62), .A0_f (new_AGEMA_signal_11999), .A1_t (new_AGEMA_signal_12000), .A1_f (new_AGEMA_signal_12001), .B0_t (SubBytesIns_Inst_Sbox_6_L5), .B0_f (new_AGEMA_signal_12011), .B1_t (new_AGEMA_signal_12012), .B1_f (new_AGEMA_signal_12013), .Z0_t (SubBytesIns_Inst_Sbox_6_L6), .Z0_f (new_AGEMA_signal_12569), .Z1_t (new_AGEMA_signal_12570), .Z1_f (new_AGEMA_signal_12571) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M46), .A0_f (new_AGEMA_signal_11339), .A1_t (new_AGEMA_signal_11340), .A1_f (new_AGEMA_signal_11341), .B0_t (SubBytesIns_Inst_Sbox_6_L3), .B0_f (new_AGEMA_signal_12005), .B1_t (new_AGEMA_signal_12006), .B1_f (new_AGEMA_signal_12007), .Z0_t (SubBytesIns_Inst_Sbox_6_L7), .Z0_f (new_AGEMA_signal_12572), .Z1_t (new_AGEMA_signal_12573), .Z1_f (new_AGEMA_signal_12574) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M51), .A0_f (new_AGEMA_signal_10637), .A1_t (new_AGEMA_signal_10638), .A1_f (new_AGEMA_signal_10639), .B0_t (SubBytesIns_Inst_Sbox_6_M59), .B0_f (new_AGEMA_signal_10646), .B1_t (new_AGEMA_signal_10647), .B1_f (new_AGEMA_signal_10648), .Z0_t (SubBytesIns_Inst_Sbox_6_L8), .Z0_f (new_AGEMA_signal_11366), .Z1_t (new_AGEMA_signal_11367), .Z1_f (new_AGEMA_signal_11368) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M52), .A0_f (new_AGEMA_signal_11345), .A1_t (new_AGEMA_signal_11346), .A1_f (new_AGEMA_signal_11347), .B0_t (SubBytesIns_Inst_Sbox_6_M53), .B0_f (new_AGEMA_signal_11996), .B1_t (new_AGEMA_signal_11997), .B1_f (new_AGEMA_signal_11998), .Z0_t (SubBytesIns_Inst_Sbox_6_L9), .Z0_f (new_AGEMA_signal_12575), .Z1_t (new_AGEMA_signal_12576), .Z1_f (new_AGEMA_signal_12577) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M53), .A0_f (new_AGEMA_signal_11996), .A1_t (new_AGEMA_signal_11997), .A1_f (new_AGEMA_signal_11998), .B0_t (SubBytesIns_Inst_Sbox_6_L4), .B0_f (new_AGEMA_signal_12008), .B1_t (new_AGEMA_signal_12009), .B1_f (new_AGEMA_signal_12010), .Z0_t (SubBytesIns_Inst_Sbox_6_L10), .Z0_f (new_AGEMA_signal_12578), .Z1_t (new_AGEMA_signal_12579), .Z1_f (new_AGEMA_signal_12580) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M60), .A0_f (new_AGEMA_signal_10649), .A1_t (new_AGEMA_signal_10650), .A1_f (new_AGEMA_signal_10651), .B0_t (SubBytesIns_Inst_Sbox_6_L2), .B0_f (new_AGEMA_signal_12002), .B1_t (new_AGEMA_signal_12003), .B1_f (new_AGEMA_signal_12004), .Z0_t (SubBytesIns_Inst_Sbox_6_L11), .Z0_f (new_AGEMA_signal_12581), .Z1_t (new_AGEMA_signal_12582), .Z1_f (new_AGEMA_signal_12583) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M48), .A0_f (new_AGEMA_signal_10631), .A1_t (new_AGEMA_signal_10632), .A1_f (new_AGEMA_signal_10633), .B0_t (SubBytesIns_Inst_Sbox_6_M51), .B0_f (new_AGEMA_signal_10637), .B1_t (new_AGEMA_signal_10638), .B1_f (new_AGEMA_signal_10639), .Z0_t (SubBytesIns_Inst_Sbox_6_L12), .Z0_f (new_AGEMA_signal_11369), .Z1_t (new_AGEMA_signal_11370), .Z1_f (new_AGEMA_signal_11371) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M50), .A0_f (new_AGEMA_signal_10634), .A1_t (new_AGEMA_signal_10635), .A1_f (new_AGEMA_signal_10636), .B0_t (SubBytesIns_Inst_Sbox_6_L0), .B0_f (new_AGEMA_signal_12566), .B1_t (new_AGEMA_signal_12567), .B1_f (new_AGEMA_signal_12568), .Z0_t (SubBytesIns_Inst_Sbox_6_L13), .Z0_f (new_AGEMA_signal_13166), .Z1_t (new_AGEMA_signal_13167), .Z1_f (new_AGEMA_signal_13168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M52), .A0_f (new_AGEMA_signal_11345), .A1_t (new_AGEMA_signal_11346), .A1_f (new_AGEMA_signal_11347), .B0_t (SubBytesIns_Inst_Sbox_6_M61), .B0_f (new_AGEMA_signal_11357), .B1_t (new_AGEMA_signal_11358), .B1_f (new_AGEMA_signal_11359), .Z0_t (SubBytesIns_Inst_Sbox_6_L14), .Z0_f (new_AGEMA_signal_12014), .Z1_t (new_AGEMA_signal_12015), .Z1_f (new_AGEMA_signal_12016) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M55), .A0_f (new_AGEMA_signal_11351), .A1_t (new_AGEMA_signal_11352), .A1_f (new_AGEMA_signal_11353), .B0_t (SubBytesIns_Inst_Sbox_6_L1), .B0_f (new_AGEMA_signal_11363), .B1_t (new_AGEMA_signal_11364), .B1_f (new_AGEMA_signal_11365), .Z0_t (SubBytesIns_Inst_Sbox_6_L15), .Z0_f (new_AGEMA_signal_12017), .Z1_t (new_AGEMA_signal_12018), .Z1_f (new_AGEMA_signal_12019) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M56), .A0_f (new_AGEMA_signal_10640), .A1_t (new_AGEMA_signal_10641), .A1_f (new_AGEMA_signal_10642), .B0_t (SubBytesIns_Inst_Sbox_6_L0), .B0_f (new_AGEMA_signal_12566), .B1_t (new_AGEMA_signal_12567), .B1_f (new_AGEMA_signal_12568), .Z0_t (SubBytesIns_Inst_Sbox_6_L16), .Z0_f (new_AGEMA_signal_13169), .Z1_t (new_AGEMA_signal_13170), .Z1_f (new_AGEMA_signal_13171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M57), .A0_f (new_AGEMA_signal_10643), .A1_t (new_AGEMA_signal_10644), .A1_f (new_AGEMA_signal_10645), .B0_t (SubBytesIns_Inst_Sbox_6_L1), .B0_f (new_AGEMA_signal_11363), .B1_t (new_AGEMA_signal_11364), .B1_f (new_AGEMA_signal_11365), .Z0_t (SubBytesIns_Inst_Sbox_6_L17), .Z0_f (new_AGEMA_signal_12020), .Z1_t (new_AGEMA_signal_12021), .Z1_f (new_AGEMA_signal_12022) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M58), .A0_f (new_AGEMA_signal_11354), .A1_t (new_AGEMA_signal_11355), .A1_f (new_AGEMA_signal_11356), .B0_t (SubBytesIns_Inst_Sbox_6_L8), .B0_f (new_AGEMA_signal_11366), .B1_t (new_AGEMA_signal_11367), .B1_f (new_AGEMA_signal_11368), .Z0_t (SubBytesIns_Inst_Sbox_6_L18), .Z0_f (new_AGEMA_signal_12023), .Z1_t (new_AGEMA_signal_12024), .Z1_f (new_AGEMA_signal_12025) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M63), .A0_f (new_AGEMA_signal_11360), .A1_t (new_AGEMA_signal_11361), .A1_f (new_AGEMA_signal_11362), .B0_t (SubBytesIns_Inst_Sbox_6_L4), .B0_f (new_AGEMA_signal_12008), .B1_t (new_AGEMA_signal_12009), .B1_f (new_AGEMA_signal_12010), .Z0_t (SubBytesIns_Inst_Sbox_6_L19), .Z0_f (new_AGEMA_signal_12584), .Z1_t (new_AGEMA_signal_12585), .Z1_f (new_AGEMA_signal_12586) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L0), .A0_f (new_AGEMA_signal_12566), .A1_t (new_AGEMA_signal_12567), .A1_f (new_AGEMA_signal_12568), .B0_t (SubBytesIns_Inst_Sbox_6_L1), .B0_f (new_AGEMA_signal_11363), .B1_t (new_AGEMA_signal_11364), .B1_f (new_AGEMA_signal_11365), .Z0_t (SubBytesIns_Inst_Sbox_6_L20), .Z0_f (new_AGEMA_signal_13172), .Z1_t (new_AGEMA_signal_13173), .Z1_f (new_AGEMA_signal_13174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L1), .A0_f (new_AGEMA_signal_11363), .A1_t (new_AGEMA_signal_11364), .A1_f (new_AGEMA_signal_11365), .B0_t (SubBytesIns_Inst_Sbox_6_L7), .B0_f (new_AGEMA_signal_12572), .B1_t (new_AGEMA_signal_12573), .B1_f (new_AGEMA_signal_12574), .Z0_t (SubBytesIns_Inst_Sbox_6_L21), .Z0_f (new_AGEMA_signal_13175), .Z1_t (new_AGEMA_signal_13176), .Z1_f (new_AGEMA_signal_13177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L3), .A0_f (new_AGEMA_signal_12005), .A1_t (new_AGEMA_signal_12006), .A1_f (new_AGEMA_signal_12007), .B0_t (SubBytesIns_Inst_Sbox_6_L12), .B0_f (new_AGEMA_signal_11369), .B1_t (new_AGEMA_signal_11370), .B1_f (new_AGEMA_signal_11371), .Z0_t (SubBytesIns_Inst_Sbox_6_L22), .Z0_f (new_AGEMA_signal_12587), .Z1_t (new_AGEMA_signal_12588), .Z1_f (new_AGEMA_signal_12589) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L18), .A0_f (new_AGEMA_signal_12023), .A1_t (new_AGEMA_signal_12024), .A1_f (new_AGEMA_signal_12025), .B0_t (SubBytesIns_Inst_Sbox_6_L2), .B0_f (new_AGEMA_signal_12002), .B1_t (new_AGEMA_signal_12003), .B1_f (new_AGEMA_signal_12004), .Z0_t (SubBytesIns_Inst_Sbox_6_L23), .Z0_f (new_AGEMA_signal_12590), .Z1_t (new_AGEMA_signal_12591), .Z1_f (new_AGEMA_signal_12592) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L15), .A0_f (new_AGEMA_signal_12017), .A1_t (new_AGEMA_signal_12018), .A1_f (new_AGEMA_signal_12019), .B0_t (SubBytesIns_Inst_Sbox_6_L9), .B0_f (new_AGEMA_signal_12575), .B1_t (new_AGEMA_signal_12576), .B1_f (new_AGEMA_signal_12577), .Z0_t (SubBytesIns_Inst_Sbox_6_L24), .Z0_f (new_AGEMA_signal_13178), .Z1_t (new_AGEMA_signal_13179), .Z1_f (new_AGEMA_signal_13180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L6), .A0_f (new_AGEMA_signal_12569), .A1_t (new_AGEMA_signal_12570), .A1_f (new_AGEMA_signal_12571), .B0_t (SubBytesIns_Inst_Sbox_6_L10), .B0_f (new_AGEMA_signal_12578), .B1_t (new_AGEMA_signal_12579), .B1_f (new_AGEMA_signal_12580), .Z0_t (SubBytesIns_Inst_Sbox_6_L25), .Z0_f (new_AGEMA_signal_13181), .Z1_t (new_AGEMA_signal_13182), .Z1_f (new_AGEMA_signal_13183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L7), .A0_f (new_AGEMA_signal_12572), .A1_t (new_AGEMA_signal_12573), .A1_f (new_AGEMA_signal_12574), .B0_t (SubBytesIns_Inst_Sbox_6_L9), .B0_f (new_AGEMA_signal_12575), .B1_t (new_AGEMA_signal_12576), .B1_f (new_AGEMA_signal_12577), .Z0_t (SubBytesIns_Inst_Sbox_6_L26), .Z0_f (new_AGEMA_signal_13184), .Z1_t (new_AGEMA_signal_13185), .Z1_f (new_AGEMA_signal_13186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L8), .A0_f (new_AGEMA_signal_11366), .A1_t (new_AGEMA_signal_11367), .A1_f (new_AGEMA_signal_11368), .B0_t (SubBytesIns_Inst_Sbox_6_L10), .B0_f (new_AGEMA_signal_12578), .B1_t (new_AGEMA_signal_12579), .B1_f (new_AGEMA_signal_12580), .Z0_t (SubBytesIns_Inst_Sbox_6_L27), .Z0_f (new_AGEMA_signal_13187), .Z1_t (new_AGEMA_signal_13188), .Z1_f (new_AGEMA_signal_13189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L11), .A0_f (new_AGEMA_signal_12581), .A1_t (new_AGEMA_signal_12582), .A1_f (new_AGEMA_signal_12583), .B0_t (SubBytesIns_Inst_Sbox_6_L14), .B0_f (new_AGEMA_signal_12014), .B1_t (new_AGEMA_signal_12015), .B1_f (new_AGEMA_signal_12016), .Z0_t (SubBytesIns_Inst_Sbox_6_L28), .Z0_f (new_AGEMA_signal_13190), .Z1_t (new_AGEMA_signal_13191), .Z1_f (new_AGEMA_signal_13192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L11), .A0_f (new_AGEMA_signal_12581), .A1_t (new_AGEMA_signal_12582), .A1_f (new_AGEMA_signal_12583), .B0_t (SubBytesIns_Inst_Sbox_6_L17), .B0_f (new_AGEMA_signal_12020), .B1_t (new_AGEMA_signal_12021), .B1_f (new_AGEMA_signal_12022), .Z0_t (SubBytesIns_Inst_Sbox_6_L29), .Z0_f (new_AGEMA_signal_13193), .Z1_t (new_AGEMA_signal_13194), .Z1_f (new_AGEMA_signal_13195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L6), .A0_f (new_AGEMA_signal_12569), .A1_t (new_AGEMA_signal_12570), .A1_f (new_AGEMA_signal_12571), .B0_t (SubBytesIns_Inst_Sbox_6_L24), .B0_f (new_AGEMA_signal_13178), .B1_t (new_AGEMA_signal_13179), .B1_f (new_AGEMA_signal_13180), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .Z0_f (new_AGEMA_signal_13766), .Z1_t (new_AGEMA_signal_13767), .Z1_f (new_AGEMA_signal_13768) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L16), .A0_f (new_AGEMA_signal_13169), .A1_t (new_AGEMA_signal_13170), .A1_f (new_AGEMA_signal_13171), .B0_t (SubBytesIns_Inst_Sbox_6_L26), .B0_f (new_AGEMA_signal_13184), .B1_t (new_AGEMA_signal_13185), .B1_f (new_AGEMA_signal_13186), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .Z0_f (new_AGEMA_signal_13769), .Z1_t (new_AGEMA_signal_13770), .Z1_f (new_AGEMA_signal_13771) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L19), .A0_f (new_AGEMA_signal_12584), .A1_t (new_AGEMA_signal_12585), .A1_f (new_AGEMA_signal_12586), .B0_t (SubBytesIns_Inst_Sbox_6_L28), .B0_f (new_AGEMA_signal_13190), .B1_t (new_AGEMA_signal_13191), .B1_f (new_AGEMA_signal_13192), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .Z0_f (new_AGEMA_signal_13772), .Z1_t (new_AGEMA_signal_13773), .Z1_f (new_AGEMA_signal_13774) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L6), .A0_f (new_AGEMA_signal_12569), .A1_t (new_AGEMA_signal_12570), .A1_f (new_AGEMA_signal_12571), .B0_t (SubBytesIns_Inst_Sbox_6_L21), .B0_f (new_AGEMA_signal_13175), .B1_t (new_AGEMA_signal_13176), .B1_f (new_AGEMA_signal_13177), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .Z0_f (new_AGEMA_signal_13775), .Z1_t (new_AGEMA_signal_13776), .Z1_f (new_AGEMA_signal_13777) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L20), .A0_f (new_AGEMA_signal_13172), .A1_t (new_AGEMA_signal_13173), .A1_f (new_AGEMA_signal_13174), .B0_t (SubBytesIns_Inst_Sbox_6_L22), .B0_f (new_AGEMA_signal_12587), .B1_t (new_AGEMA_signal_12588), .B1_f (new_AGEMA_signal_12589), .Z0_t (MixColumnsInput[83]), .Z0_f (new_AGEMA_signal_13778), .Z1_t (new_AGEMA_signal_13779), .Z1_f (new_AGEMA_signal_13780) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L25), .A0_f (new_AGEMA_signal_13181), .A1_t (new_AGEMA_signal_13182), .A1_f (new_AGEMA_signal_13183), .B0_t (SubBytesIns_Inst_Sbox_6_L29), .B0_f (new_AGEMA_signal_13193), .B1_t (new_AGEMA_signal_13194), .B1_f (new_AGEMA_signal_13195), .Z0_t (MixColumnsInput[82]), .Z0_f (new_AGEMA_signal_13781), .Z1_t (new_AGEMA_signal_13782), .Z1_f (new_AGEMA_signal_13783) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L13), .A0_f (new_AGEMA_signal_13166), .A1_t (new_AGEMA_signal_13167), .A1_f (new_AGEMA_signal_13168), .B0_t (SubBytesIns_Inst_Sbox_6_L27), .B0_f (new_AGEMA_signal_13187), .B1_t (new_AGEMA_signal_13188), .B1_f (new_AGEMA_signal_13189), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .Z0_f (new_AGEMA_signal_13784), .Z1_t (new_AGEMA_signal_13785), .Z1_f (new_AGEMA_signal_13786) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L6), .A0_f (new_AGEMA_signal_12569), .A1_t (new_AGEMA_signal_12570), .A1_f (new_AGEMA_signal_12571), .B0_t (SubBytesIns_Inst_Sbox_6_L23), .B0_f (new_AGEMA_signal_12590), .B1_t (new_AGEMA_signal_12591), .B1_f (new_AGEMA_signal_12592), .Z0_t (MixColumnsInput[80]), .Z0_f (new_AGEMA_signal_13196), .Z1_t (new_AGEMA_signal_13197), .Z1_f (new_AGEMA_signal_13198) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[63]), .A0_f (ciphertext_s0_f[63]), .A1_t (ciphertext_s1_t[63]), .A1_f (ciphertext_s1_f[63]), .B0_t (ciphertext_s0_t[60]), .B0_f (ciphertext_s0_f[60]), .B1_t (ciphertext_s1_t[60]), .B1_f (ciphertext_s1_f[60]), .Z0_t (SubBytesIns_Inst_Sbox_7_T1), .Z0_f (new_AGEMA_signal_6556), .Z1_t (new_AGEMA_signal_6557), .Z1_f (new_AGEMA_signal_6558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[63]), .A0_f (ciphertext_s0_f[63]), .A1_t (ciphertext_s1_t[63]), .A1_f (ciphertext_s1_f[63]), .B0_t (ciphertext_s0_t[58]), .B0_f (ciphertext_s0_f[58]), .B1_t (ciphertext_s1_t[58]), .B1_f (ciphertext_s1_f[58]), .Z0_t (SubBytesIns_Inst_Sbox_7_T2), .Z0_f (new_AGEMA_signal_6559), .Z1_t (new_AGEMA_signal_6560), .Z1_f (new_AGEMA_signal_6561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[63]), .A0_f (ciphertext_s0_f[63]), .A1_t (ciphertext_s1_t[63]), .A1_f (ciphertext_s1_f[63]), .B0_t (ciphertext_s0_t[57]), .B0_f (ciphertext_s0_f[57]), .B1_t (ciphertext_s1_t[57]), .B1_f (ciphertext_s1_f[57]), .Z0_t (SubBytesIns_Inst_Sbox_7_T3), .Z0_f (new_AGEMA_signal_6562), .Z1_t (new_AGEMA_signal_6563), .Z1_f (new_AGEMA_signal_6564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[60]), .A0_f (ciphertext_s0_f[60]), .A1_t (ciphertext_s1_t[60]), .A1_f (ciphertext_s1_f[60]), .B0_t (ciphertext_s0_t[58]), .B0_f (ciphertext_s0_f[58]), .B1_t (ciphertext_s1_t[58]), .B1_f (ciphertext_s1_f[58]), .Z0_t (SubBytesIns_Inst_Sbox_7_T4), .Z0_f (new_AGEMA_signal_6565), .Z1_t (new_AGEMA_signal_6566), .Z1_f (new_AGEMA_signal_6567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[59]), .A0_f (ciphertext_s0_f[59]), .A1_t (ciphertext_s1_t[59]), .A1_f (ciphertext_s1_f[59]), .B0_t (ciphertext_s0_t[57]), .B0_f (ciphertext_s0_f[57]), .B1_t (ciphertext_s1_t[57]), .B1_f (ciphertext_s1_f[57]), .Z0_t (SubBytesIns_Inst_Sbox_7_T5), .Z0_f (new_AGEMA_signal_6568), .Z1_t (new_AGEMA_signal_6569), .Z1_f (new_AGEMA_signal_6570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T1), .A0_f (new_AGEMA_signal_6556), .A1_t (new_AGEMA_signal_6557), .A1_f (new_AGEMA_signal_6558), .B0_t (SubBytesIns_Inst_Sbox_7_T5), .B0_f (new_AGEMA_signal_6568), .B1_t (new_AGEMA_signal_6569), .B1_f (new_AGEMA_signal_6570), .Z0_t (SubBytesIns_Inst_Sbox_7_T6), .Z0_f (new_AGEMA_signal_7096), .Z1_t (new_AGEMA_signal_7097), .Z1_f (new_AGEMA_signal_7098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[62]), .A0_f (ciphertext_s0_f[62]), .A1_t (ciphertext_s1_t[62]), .A1_f (ciphertext_s1_f[62]), .B0_t (ciphertext_s0_t[61]), .B0_f (ciphertext_s0_f[61]), .B1_t (ciphertext_s1_t[61]), .B1_f (ciphertext_s1_f[61]), .Z0_t (SubBytesIns_Inst_Sbox_7_T7), .Z0_f (new_AGEMA_signal_6571), .Z1_t (new_AGEMA_signal_6572), .Z1_f (new_AGEMA_signal_6573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[56]), .A0_f (ciphertext_s0_f[56]), .A1_t (ciphertext_s1_t[56]), .A1_f (ciphertext_s1_f[56]), .B0_t (SubBytesIns_Inst_Sbox_7_T6), .B0_f (new_AGEMA_signal_7096), .B1_t (new_AGEMA_signal_7097), .B1_f (new_AGEMA_signal_7098), .Z0_t (SubBytesIns_Inst_Sbox_7_T8), .Z0_f (new_AGEMA_signal_7745), .Z1_t (new_AGEMA_signal_7746), .Z1_f (new_AGEMA_signal_7747) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[56]), .A0_f (ciphertext_s0_f[56]), .A1_t (ciphertext_s1_t[56]), .A1_f (ciphertext_s1_f[56]), .B0_t (SubBytesIns_Inst_Sbox_7_T7), .B0_f (new_AGEMA_signal_6571), .B1_t (new_AGEMA_signal_6572), .B1_f (new_AGEMA_signal_6573), .Z0_t (SubBytesIns_Inst_Sbox_7_T9), .Z0_f (new_AGEMA_signal_7099), .Z1_t (new_AGEMA_signal_7100), .Z1_f (new_AGEMA_signal_7101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T6), .A0_f (new_AGEMA_signal_7096), .A1_t (new_AGEMA_signal_7097), .A1_f (new_AGEMA_signal_7098), .B0_t (SubBytesIns_Inst_Sbox_7_T7), .B0_f (new_AGEMA_signal_6571), .B1_t (new_AGEMA_signal_6572), .B1_f (new_AGEMA_signal_6573), .Z0_t (SubBytesIns_Inst_Sbox_7_T10), .Z0_f (new_AGEMA_signal_7748), .Z1_t (new_AGEMA_signal_7749), .Z1_f (new_AGEMA_signal_7750) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[62]), .A0_f (ciphertext_s0_f[62]), .A1_t (ciphertext_s1_t[62]), .A1_f (ciphertext_s1_f[62]), .B0_t (ciphertext_s0_t[58]), .B0_f (ciphertext_s0_f[58]), .B1_t (ciphertext_s1_t[58]), .B1_f (ciphertext_s1_f[58]), .Z0_t (SubBytesIns_Inst_Sbox_7_T11), .Z0_f (new_AGEMA_signal_6574), .Z1_t (new_AGEMA_signal_6575), .Z1_f (new_AGEMA_signal_6576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[61]), .A0_f (ciphertext_s0_f[61]), .A1_t (ciphertext_s1_t[61]), .A1_f (ciphertext_s1_f[61]), .B0_t (ciphertext_s0_t[58]), .B0_f (ciphertext_s0_f[58]), .B1_t (ciphertext_s1_t[58]), .B1_f (ciphertext_s1_f[58]), .Z0_t (SubBytesIns_Inst_Sbox_7_T12), .Z0_f (new_AGEMA_signal_6577), .Z1_t (new_AGEMA_signal_6578), .Z1_f (new_AGEMA_signal_6579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T3), .A0_f (new_AGEMA_signal_6562), .A1_t (new_AGEMA_signal_6563), .A1_f (new_AGEMA_signal_6564), .B0_t (SubBytesIns_Inst_Sbox_7_T4), .B0_f (new_AGEMA_signal_6565), .B1_t (new_AGEMA_signal_6566), .B1_f (new_AGEMA_signal_6567), .Z0_t (SubBytesIns_Inst_Sbox_7_T13), .Z0_f (new_AGEMA_signal_7102), .Z1_t (new_AGEMA_signal_7103), .Z1_f (new_AGEMA_signal_7104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T6), .A0_f (new_AGEMA_signal_7096), .A1_t (new_AGEMA_signal_7097), .A1_f (new_AGEMA_signal_7098), .B0_t (SubBytesIns_Inst_Sbox_7_T11), .B0_f (new_AGEMA_signal_6574), .B1_t (new_AGEMA_signal_6575), .B1_f (new_AGEMA_signal_6576), .Z0_t (SubBytesIns_Inst_Sbox_7_T14), .Z0_f (new_AGEMA_signal_7751), .Z1_t (new_AGEMA_signal_7752), .Z1_f (new_AGEMA_signal_7753) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T5), .A0_f (new_AGEMA_signal_6568), .A1_t (new_AGEMA_signal_6569), .A1_f (new_AGEMA_signal_6570), .B0_t (SubBytesIns_Inst_Sbox_7_T11), .B0_f (new_AGEMA_signal_6574), .B1_t (new_AGEMA_signal_6575), .B1_f (new_AGEMA_signal_6576), .Z0_t (SubBytesIns_Inst_Sbox_7_T15), .Z0_f (new_AGEMA_signal_7105), .Z1_t (new_AGEMA_signal_7106), .Z1_f (new_AGEMA_signal_7107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T5), .A0_f (new_AGEMA_signal_6568), .A1_t (new_AGEMA_signal_6569), .A1_f (new_AGEMA_signal_6570), .B0_t (SubBytesIns_Inst_Sbox_7_T12), .B0_f (new_AGEMA_signal_6577), .B1_t (new_AGEMA_signal_6578), .B1_f (new_AGEMA_signal_6579), .Z0_t (SubBytesIns_Inst_Sbox_7_T16), .Z0_f (new_AGEMA_signal_7108), .Z1_t (new_AGEMA_signal_7109), .Z1_f (new_AGEMA_signal_7110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T9), .A0_f (new_AGEMA_signal_7099), .A1_t (new_AGEMA_signal_7100), .A1_f (new_AGEMA_signal_7101), .B0_t (SubBytesIns_Inst_Sbox_7_T16), .B0_f (new_AGEMA_signal_7108), .B1_t (new_AGEMA_signal_7109), .B1_f (new_AGEMA_signal_7110), .Z0_t (SubBytesIns_Inst_Sbox_7_T17), .Z0_f (new_AGEMA_signal_7754), .Z1_t (new_AGEMA_signal_7755), .Z1_f (new_AGEMA_signal_7756) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[60]), .A0_f (ciphertext_s0_f[60]), .A1_t (ciphertext_s1_t[60]), .A1_f (ciphertext_s1_f[60]), .B0_t (ciphertext_s0_t[56]), .B0_f (ciphertext_s0_f[56]), .B1_t (ciphertext_s1_t[56]), .B1_f (ciphertext_s1_f[56]), .Z0_t (SubBytesIns_Inst_Sbox_7_T18), .Z0_f (new_AGEMA_signal_6580), .Z1_t (new_AGEMA_signal_6581), .Z1_f (new_AGEMA_signal_6582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T7), .A0_f (new_AGEMA_signal_6571), .A1_t (new_AGEMA_signal_6572), .A1_f (new_AGEMA_signal_6573), .B0_t (SubBytesIns_Inst_Sbox_7_T18), .B0_f (new_AGEMA_signal_6580), .B1_t (new_AGEMA_signal_6581), .B1_f (new_AGEMA_signal_6582), .Z0_t (SubBytesIns_Inst_Sbox_7_T19), .Z0_f (new_AGEMA_signal_7111), .Z1_t (new_AGEMA_signal_7112), .Z1_f (new_AGEMA_signal_7113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T1), .A0_f (new_AGEMA_signal_6556), .A1_t (new_AGEMA_signal_6557), .A1_f (new_AGEMA_signal_6558), .B0_t (SubBytesIns_Inst_Sbox_7_T19), .B0_f (new_AGEMA_signal_7111), .B1_t (new_AGEMA_signal_7112), .B1_f (new_AGEMA_signal_7113), .Z0_t (SubBytesIns_Inst_Sbox_7_T20), .Z0_f (new_AGEMA_signal_7757), .Z1_t (new_AGEMA_signal_7758), .Z1_f (new_AGEMA_signal_7759) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[57]), .A0_f (ciphertext_s0_f[57]), .A1_t (ciphertext_s1_t[57]), .A1_f (ciphertext_s1_f[57]), .B0_t (ciphertext_s0_t[56]), .B0_f (ciphertext_s0_f[56]), .B1_t (ciphertext_s1_t[56]), .B1_f (ciphertext_s1_f[56]), .Z0_t (SubBytesIns_Inst_Sbox_7_T21), .Z0_f (new_AGEMA_signal_6583), .Z1_t (new_AGEMA_signal_6584), .Z1_f (new_AGEMA_signal_6585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T7), .A0_f (new_AGEMA_signal_6571), .A1_t (new_AGEMA_signal_6572), .A1_f (new_AGEMA_signal_6573), .B0_t (SubBytesIns_Inst_Sbox_7_T21), .B0_f (new_AGEMA_signal_6583), .B1_t (new_AGEMA_signal_6584), .B1_f (new_AGEMA_signal_6585), .Z0_t (SubBytesIns_Inst_Sbox_7_T22), .Z0_f (new_AGEMA_signal_7114), .Z1_t (new_AGEMA_signal_7115), .Z1_f (new_AGEMA_signal_7116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T2), .A0_f (new_AGEMA_signal_6559), .A1_t (new_AGEMA_signal_6560), .A1_f (new_AGEMA_signal_6561), .B0_t (SubBytesIns_Inst_Sbox_7_T22), .B0_f (new_AGEMA_signal_7114), .B1_t (new_AGEMA_signal_7115), .B1_f (new_AGEMA_signal_7116), .Z0_t (SubBytesIns_Inst_Sbox_7_T23), .Z0_f (new_AGEMA_signal_7760), .Z1_t (new_AGEMA_signal_7761), .Z1_f (new_AGEMA_signal_7762) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T2), .A0_f (new_AGEMA_signal_6559), .A1_t (new_AGEMA_signal_6560), .A1_f (new_AGEMA_signal_6561), .B0_t (SubBytesIns_Inst_Sbox_7_T10), .B0_f (new_AGEMA_signal_7748), .B1_t (new_AGEMA_signal_7749), .B1_f (new_AGEMA_signal_7750), .Z0_t (SubBytesIns_Inst_Sbox_7_T24), .Z0_f (new_AGEMA_signal_8393), .Z1_t (new_AGEMA_signal_8394), .Z1_f (new_AGEMA_signal_8395) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T20), .A0_f (new_AGEMA_signal_7757), .A1_t (new_AGEMA_signal_7758), .A1_f (new_AGEMA_signal_7759), .B0_t (SubBytesIns_Inst_Sbox_7_T17), .B0_f (new_AGEMA_signal_7754), .B1_t (new_AGEMA_signal_7755), .B1_f (new_AGEMA_signal_7756), .Z0_t (SubBytesIns_Inst_Sbox_7_T25), .Z0_f (new_AGEMA_signal_8396), .Z1_t (new_AGEMA_signal_8397), .Z1_f (new_AGEMA_signal_8398) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T3), .A0_f (new_AGEMA_signal_6562), .A1_t (new_AGEMA_signal_6563), .A1_f (new_AGEMA_signal_6564), .B0_t (SubBytesIns_Inst_Sbox_7_T16), .B0_f (new_AGEMA_signal_7108), .B1_t (new_AGEMA_signal_7109), .B1_f (new_AGEMA_signal_7110), .Z0_t (SubBytesIns_Inst_Sbox_7_T26), .Z0_f (new_AGEMA_signal_7763), .Z1_t (new_AGEMA_signal_7764), .Z1_f (new_AGEMA_signal_7765) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T1), .A0_f (new_AGEMA_signal_6556), .A1_t (new_AGEMA_signal_6557), .A1_f (new_AGEMA_signal_6558), .B0_t (SubBytesIns_Inst_Sbox_7_T12), .B0_f (new_AGEMA_signal_6577), .B1_t (new_AGEMA_signal_6578), .B1_f (new_AGEMA_signal_6579), .Z0_t (SubBytesIns_Inst_Sbox_7_T27), .Z0_f (new_AGEMA_signal_7117), .Z1_t (new_AGEMA_signal_7118), .Z1_f (new_AGEMA_signal_7119) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T13), .A0_f (new_AGEMA_signal_7102), .A1_t (new_AGEMA_signal_7103), .A1_f (new_AGEMA_signal_7104), .B0_t (SubBytesIns_Inst_Sbox_7_T6), .B0_f (new_AGEMA_signal_7096), .B1_t (new_AGEMA_signal_7097), .B1_f (new_AGEMA_signal_7098), .Z0_t (SubBytesIns_Inst_Sbox_7_M1), .Z0_f (new_AGEMA_signal_7766), .Z1_t (new_AGEMA_signal_7767), .Z1_f (new_AGEMA_signal_7768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T23), .A0_f (new_AGEMA_signal_7760), .A1_t (new_AGEMA_signal_7761), .A1_f (new_AGEMA_signal_7762), .B0_t (SubBytesIns_Inst_Sbox_7_T8), .B0_f (new_AGEMA_signal_7745), .B1_t (new_AGEMA_signal_7746), .B1_f (new_AGEMA_signal_7747), .Z0_t (SubBytesIns_Inst_Sbox_7_M2), .Z0_f (new_AGEMA_signal_8399), .Z1_t (new_AGEMA_signal_8400), .Z1_f (new_AGEMA_signal_8401) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T14), .A0_f (new_AGEMA_signal_7751), .A1_t (new_AGEMA_signal_7752), .A1_f (new_AGEMA_signal_7753), .B0_t (SubBytesIns_Inst_Sbox_7_M1), .B0_f (new_AGEMA_signal_7766), .B1_t (new_AGEMA_signal_7767), .B1_f (new_AGEMA_signal_7768), .Z0_t (SubBytesIns_Inst_Sbox_7_M3), .Z0_f (new_AGEMA_signal_8402), .Z1_t (new_AGEMA_signal_8403), .Z1_f (new_AGEMA_signal_8404) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T19), .A0_f (new_AGEMA_signal_7111), .A1_t (new_AGEMA_signal_7112), .A1_f (new_AGEMA_signal_7113), .B0_t (ciphertext_s0_t[56]), .B0_f (ciphertext_s0_f[56]), .B1_t (ciphertext_s1_t[56]), .B1_f (ciphertext_s1_f[56]), .Z0_t (SubBytesIns_Inst_Sbox_7_M4), .Z0_f (new_AGEMA_signal_7769), .Z1_t (new_AGEMA_signal_7770), .Z1_f (new_AGEMA_signal_7771) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M4), .A0_f (new_AGEMA_signal_7769), .A1_t (new_AGEMA_signal_7770), .A1_f (new_AGEMA_signal_7771), .B0_t (SubBytesIns_Inst_Sbox_7_M1), .B0_f (new_AGEMA_signal_7766), .B1_t (new_AGEMA_signal_7767), .B1_f (new_AGEMA_signal_7768), .Z0_t (SubBytesIns_Inst_Sbox_7_M5), .Z0_f (new_AGEMA_signal_8405), .Z1_t (new_AGEMA_signal_8406), .Z1_f (new_AGEMA_signal_8407) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T3), .A0_f (new_AGEMA_signal_6562), .A1_t (new_AGEMA_signal_6563), .A1_f (new_AGEMA_signal_6564), .B0_t (SubBytesIns_Inst_Sbox_7_T16), .B0_f (new_AGEMA_signal_7108), .B1_t (new_AGEMA_signal_7109), .B1_f (new_AGEMA_signal_7110), .Z0_t (SubBytesIns_Inst_Sbox_7_M6), .Z0_f (new_AGEMA_signal_7772), .Z1_t (new_AGEMA_signal_7773), .Z1_f (new_AGEMA_signal_7774) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T22), .A0_f (new_AGEMA_signal_7114), .A1_t (new_AGEMA_signal_7115), .A1_f (new_AGEMA_signal_7116), .B0_t (SubBytesIns_Inst_Sbox_7_T9), .B0_f (new_AGEMA_signal_7099), .B1_t (new_AGEMA_signal_7100), .B1_f (new_AGEMA_signal_7101), .Z0_t (SubBytesIns_Inst_Sbox_7_M7), .Z0_f (new_AGEMA_signal_7775), .Z1_t (new_AGEMA_signal_7776), .Z1_f (new_AGEMA_signal_7777) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T26), .A0_f (new_AGEMA_signal_7763), .A1_t (new_AGEMA_signal_7764), .A1_f (new_AGEMA_signal_7765), .B0_t (SubBytesIns_Inst_Sbox_7_M6), .B0_f (new_AGEMA_signal_7772), .B1_t (new_AGEMA_signal_7773), .B1_f (new_AGEMA_signal_7774), .Z0_t (SubBytesIns_Inst_Sbox_7_M8), .Z0_f (new_AGEMA_signal_8408), .Z1_t (new_AGEMA_signal_8409), .Z1_f (new_AGEMA_signal_8410) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T20), .A0_f (new_AGEMA_signal_7757), .A1_t (new_AGEMA_signal_7758), .A1_f (new_AGEMA_signal_7759), .B0_t (SubBytesIns_Inst_Sbox_7_T17), .B0_f (new_AGEMA_signal_7754), .B1_t (new_AGEMA_signal_7755), .B1_f (new_AGEMA_signal_7756), .Z0_t (SubBytesIns_Inst_Sbox_7_M9), .Z0_f (new_AGEMA_signal_8411), .Z1_t (new_AGEMA_signal_8412), .Z1_f (new_AGEMA_signal_8413) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M9), .A0_f (new_AGEMA_signal_8411), .A1_t (new_AGEMA_signal_8412), .A1_f (new_AGEMA_signal_8413), .B0_t (SubBytesIns_Inst_Sbox_7_M6), .B0_f (new_AGEMA_signal_7772), .B1_t (new_AGEMA_signal_7773), .B1_f (new_AGEMA_signal_7774), .Z0_t (SubBytesIns_Inst_Sbox_7_M10), .Z0_f (new_AGEMA_signal_8801), .Z1_t (new_AGEMA_signal_8802), .Z1_f (new_AGEMA_signal_8803) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T1), .A0_f (new_AGEMA_signal_6556), .A1_t (new_AGEMA_signal_6557), .A1_f (new_AGEMA_signal_6558), .B0_t (SubBytesIns_Inst_Sbox_7_T15), .B0_f (new_AGEMA_signal_7105), .B1_t (new_AGEMA_signal_7106), .B1_f (new_AGEMA_signal_7107), .Z0_t (SubBytesIns_Inst_Sbox_7_M11), .Z0_f (new_AGEMA_signal_7778), .Z1_t (new_AGEMA_signal_7779), .Z1_f (new_AGEMA_signal_7780) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T4), .A0_f (new_AGEMA_signal_6565), .A1_t (new_AGEMA_signal_6566), .A1_f (new_AGEMA_signal_6567), .B0_t (SubBytesIns_Inst_Sbox_7_T27), .B0_f (new_AGEMA_signal_7117), .B1_t (new_AGEMA_signal_7118), .B1_f (new_AGEMA_signal_7119), .Z0_t (SubBytesIns_Inst_Sbox_7_M12), .Z0_f (new_AGEMA_signal_7781), .Z1_t (new_AGEMA_signal_7782), .Z1_f (new_AGEMA_signal_7783) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M12), .A0_f (new_AGEMA_signal_7781), .A1_t (new_AGEMA_signal_7782), .A1_f (new_AGEMA_signal_7783), .B0_t (SubBytesIns_Inst_Sbox_7_M11), .B0_f (new_AGEMA_signal_7778), .B1_t (new_AGEMA_signal_7779), .B1_f (new_AGEMA_signal_7780), .Z0_t (SubBytesIns_Inst_Sbox_7_M13), .Z0_f (new_AGEMA_signal_8414), .Z1_t (new_AGEMA_signal_8415), .Z1_f (new_AGEMA_signal_8416) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T2), .A0_f (new_AGEMA_signal_6559), .A1_t (new_AGEMA_signal_6560), .A1_f (new_AGEMA_signal_6561), .B0_t (SubBytesIns_Inst_Sbox_7_T10), .B0_f (new_AGEMA_signal_7748), .B1_t (new_AGEMA_signal_7749), .B1_f (new_AGEMA_signal_7750), .Z0_t (SubBytesIns_Inst_Sbox_7_M14), .Z0_f (new_AGEMA_signal_8417), .Z1_t (new_AGEMA_signal_8418), .Z1_f (new_AGEMA_signal_8419) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M14), .A0_f (new_AGEMA_signal_8417), .A1_t (new_AGEMA_signal_8418), .A1_f (new_AGEMA_signal_8419), .B0_t (SubBytesIns_Inst_Sbox_7_M11), .B0_f (new_AGEMA_signal_7778), .B1_t (new_AGEMA_signal_7779), .B1_f (new_AGEMA_signal_7780), .Z0_t (SubBytesIns_Inst_Sbox_7_M15), .Z0_f (new_AGEMA_signal_8804), .Z1_t (new_AGEMA_signal_8805), .Z1_f (new_AGEMA_signal_8806) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M3), .A0_f (new_AGEMA_signal_8402), .A1_t (new_AGEMA_signal_8403), .A1_f (new_AGEMA_signal_8404), .B0_t (SubBytesIns_Inst_Sbox_7_M2), .B0_f (new_AGEMA_signal_8399), .B1_t (new_AGEMA_signal_8400), .B1_f (new_AGEMA_signal_8401), .Z0_t (SubBytesIns_Inst_Sbox_7_M16), .Z0_f (new_AGEMA_signal_8807), .Z1_t (new_AGEMA_signal_8808), .Z1_f (new_AGEMA_signal_8809) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M5), .A0_f (new_AGEMA_signal_8405), .A1_t (new_AGEMA_signal_8406), .A1_f (new_AGEMA_signal_8407), .B0_t (SubBytesIns_Inst_Sbox_7_T24), .B0_f (new_AGEMA_signal_8393), .B1_t (new_AGEMA_signal_8394), .B1_f (new_AGEMA_signal_8395), .Z0_t (SubBytesIns_Inst_Sbox_7_M17), .Z0_f (new_AGEMA_signal_8810), .Z1_t (new_AGEMA_signal_8811), .Z1_f (new_AGEMA_signal_8812) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M8), .A0_f (new_AGEMA_signal_8408), .A1_t (new_AGEMA_signal_8409), .A1_f (new_AGEMA_signal_8410), .B0_t (SubBytesIns_Inst_Sbox_7_M7), .B0_f (new_AGEMA_signal_7775), .B1_t (new_AGEMA_signal_7776), .B1_f (new_AGEMA_signal_7777), .Z0_t (SubBytesIns_Inst_Sbox_7_M18), .Z0_f (new_AGEMA_signal_8813), .Z1_t (new_AGEMA_signal_8814), .Z1_f (new_AGEMA_signal_8815) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M10), .A0_f (new_AGEMA_signal_8801), .A1_t (new_AGEMA_signal_8802), .A1_f (new_AGEMA_signal_8803), .B0_t (SubBytesIns_Inst_Sbox_7_M15), .B0_f (new_AGEMA_signal_8804), .B1_t (new_AGEMA_signal_8805), .B1_f (new_AGEMA_signal_8806), .Z0_t (SubBytesIns_Inst_Sbox_7_M19), .Z0_f (new_AGEMA_signal_9068), .Z1_t (new_AGEMA_signal_9069), .Z1_f (new_AGEMA_signal_9070) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M16), .A0_f (new_AGEMA_signal_8807), .A1_t (new_AGEMA_signal_8808), .A1_f (new_AGEMA_signal_8809), .B0_t (SubBytesIns_Inst_Sbox_7_M13), .B0_f (new_AGEMA_signal_8414), .B1_t (new_AGEMA_signal_8415), .B1_f (new_AGEMA_signal_8416), .Z0_t (SubBytesIns_Inst_Sbox_7_M20), .Z0_f (new_AGEMA_signal_9071), .Z1_t (new_AGEMA_signal_9072), .Z1_f (new_AGEMA_signal_9073) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M17), .A0_f (new_AGEMA_signal_8810), .A1_t (new_AGEMA_signal_8811), .A1_f (new_AGEMA_signal_8812), .B0_t (SubBytesIns_Inst_Sbox_7_M15), .B0_f (new_AGEMA_signal_8804), .B1_t (new_AGEMA_signal_8805), .B1_f (new_AGEMA_signal_8806), .Z0_t (SubBytesIns_Inst_Sbox_7_M21), .Z0_f (new_AGEMA_signal_9074), .Z1_t (new_AGEMA_signal_9075), .Z1_f (new_AGEMA_signal_9076) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M18), .A0_f (new_AGEMA_signal_8813), .A1_t (new_AGEMA_signal_8814), .A1_f (new_AGEMA_signal_8815), .B0_t (SubBytesIns_Inst_Sbox_7_M13), .B0_f (new_AGEMA_signal_8414), .B1_t (new_AGEMA_signal_8415), .B1_f (new_AGEMA_signal_8416), .Z0_t (SubBytesIns_Inst_Sbox_7_M22), .Z0_f (new_AGEMA_signal_9077), .Z1_t (new_AGEMA_signal_9078), .Z1_f (new_AGEMA_signal_9079) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M19), .A0_f (new_AGEMA_signal_9068), .A1_t (new_AGEMA_signal_9069), .A1_f (new_AGEMA_signal_9070), .B0_t (SubBytesIns_Inst_Sbox_7_T25), .B0_f (new_AGEMA_signal_8396), .B1_t (new_AGEMA_signal_8397), .B1_f (new_AGEMA_signal_8398), .Z0_t (SubBytesIns_Inst_Sbox_7_M23), .Z0_f (new_AGEMA_signal_9308), .Z1_t (new_AGEMA_signal_9309), .Z1_f (new_AGEMA_signal_9310) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M22), .A0_f (new_AGEMA_signal_9077), .A1_t (new_AGEMA_signal_9078), .A1_f (new_AGEMA_signal_9079), .B0_t (SubBytesIns_Inst_Sbox_7_M23), .B0_f (new_AGEMA_signal_9308), .B1_t (new_AGEMA_signal_9309), .B1_f (new_AGEMA_signal_9310), .Z0_t (SubBytesIns_Inst_Sbox_7_M24), .Z0_f (new_AGEMA_signal_9581), .Z1_t (new_AGEMA_signal_9582), .Z1_f (new_AGEMA_signal_9583) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M22), .A0_f (new_AGEMA_signal_9077), .A1_t (new_AGEMA_signal_9078), .A1_f (new_AGEMA_signal_9079), .B0_t (SubBytesIns_Inst_Sbox_7_M20), .B0_f (new_AGEMA_signal_9071), .B1_t (new_AGEMA_signal_9072), .B1_f (new_AGEMA_signal_9073), .Z0_t (SubBytesIns_Inst_Sbox_7_M25), .Z0_f (new_AGEMA_signal_9311), .Z1_t (new_AGEMA_signal_9312), .Z1_f (new_AGEMA_signal_9313) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M21), .A0_f (new_AGEMA_signal_9074), .A1_t (new_AGEMA_signal_9075), .A1_f (new_AGEMA_signal_9076), .B0_t (SubBytesIns_Inst_Sbox_7_M25), .B0_f (new_AGEMA_signal_9311), .B1_t (new_AGEMA_signal_9312), .B1_f (new_AGEMA_signal_9313), .Z0_t (SubBytesIns_Inst_Sbox_7_M26), .Z0_f (new_AGEMA_signal_9584), .Z1_t (new_AGEMA_signal_9585), .Z1_f (new_AGEMA_signal_9586) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M20), .A0_f (new_AGEMA_signal_9071), .A1_t (new_AGEMA_signal_9072), .A1_f (new_AGEMA_signal_9073), .B0_t (SubBytesIns_Inst_Sbox_7_M21), .B0_f (new_AGEMA_signal_9074), .B1_t (new_AGEMA_signal_9075), .B1_f (new_AGEMA_signal_9076), .Z0_t (SubBytesIns_Inst_Sbox_7_M27), .Z0_f (new_AGEMA_signal_9314), .Z1_t (new_AGEMA_signal_9315), .Z1_f (new_AGEMA_signal_9316) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M23), .A0_f (new_AGEMA_signal_9308), .A1_t (new_AGEMA_signal_9309), .A1_f (new_AGEMA_signal_9310), .B0_t (SubBytesIns_Inst_Sbox_7_M25), .B0_f (new_AGEMA_signal_9311), .B1_t (new_AGEMA_signal_9312), .B1_f (new_AGEMA_signal_9313), .Z0_t (SubBytesIns_Inst_Sbox_7_M28), .Z0_f (new_AGEMA_signal_9587), .Z1_t (new_AGEMA_signal_9588), .Z1_f (new_AGEMA_signal_9589) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M28), .A0_f (new_AGEMA_signal_9587), .A1_t (new_AGEMA_signal_9588), .A1_f (new_AGEMA_signal_9589), .B0_t (SubBytesIns_Inst_Sbox_7_M27), .B0_f (new_AGEMA_signal_9314), .B1_t (new_AGEMA_signal_9315), .B1_f (new_AGEMA_signal_9316), .Z0_t (SubBytesIns_Inst_Sbox_7_M29), .Z0_f (new_AGEMA_signal_9881), .Z1_t (new_AGEMA_signal_9882), .Z1_f (new_AGEMA_signal_9883) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M26), .A0_f (new_AGEMA_signal_9584), .A1_t (new_AGEMA_signal_9585), .A1_f (new_AGEMA_signal_9586), .B0_t (SubBytesIns_Inst_Sbox_7_M24), .B0_f (new_AGEMA_signal_9581), .B1_t (new_AGEMA_signal_9582), .B1_f (new_AGEMA_signal_9583), .Z0_t (SubBytesIns_Inst_Sbox_7_M30), .Z0_f (new_AGEMA_signal_9884), .Z1_t (new_AGEMA_signal_9885), .Z1_f (new_AGEMA_signal_9886) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M20), .A0_f (new_AGEMA_signal_9071), .A1_t (new_AGEMA_signal_9072), .A1_f (new_AGEMA_signal_9073), .B0_t (SubBytesIns_Inst_Sbox_7_M23), .B0_f (new_AGEMA_signal_9308), .B1_t (new_AGEMA_signal_9309), .B1_f (new_AGEMA_signal_9310), .Z0_t (SubBytesIns_Inst_Sbox_7_M31), .Z0_f (new_AGEMA_signal_9590), .Z1_t (new_AGEMA_signal_9591), .Z1_f (new_AGEMA_signal_9592) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M27), .A0_f (new_AGEMA_signal_9314), .A1_t (new_AGEMA_signal_9315), .A1_f (new_AGEMA_signal_9316), .B0_t (SubBytesIns_Inst_Sbox_7_M31), .B0_f (new_AGEMA_signal_9590), .B1_t (new_AGEMA_signal_9591), .B1_f (new_AGEMA_signal_9592), .Z0_t (SubBytesIns_Inst_Sbox_7_M32), .Z0_f (new_AGEMA_signal_9887), .Z1_t (new_AGEMA_signal_9888), .Z1_f (new_AGEMA_signal_9889) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M27), .A0_f (new_AGEMA_signal_9314), .A1_t (new_AGEMA_signal_9315), .A1_f (new_AGEMA_signal_9316), .B0_t (SubBytesIns_Inst_Sbox_7_M25), .B0_f (new_AGEMA_signal_9311), .B1_t (new_AGEMA_signal_9312), .B1_f (new_AGEMA_signal_9313), .Z0_t (SubBytesIns_Inst_Sbox_7_M33), .Z0_f (new_AGEMA_signal_9593), .Z1_t (new_AGEMA_signal_9594), .Z1_f (new_AGEMA_signal_9595) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M21), .A0_f (new_AGEMA_signal_9074), .A1_t (new_AGEMA_signal_9075), .A1_f (new_AGEMA_signal_9076), .B0_t (SubBytesIns_Inst_Sbox_7_M22), .B0_f (new_AGEMA_signal_9077), .B1_t (new_AGEMA_signal_9078), .B1_f (new_AGEMA_signal_9079), .Z0_t (SubBytesIns_Inst_Sbox_7_M34), .Z0_f (new_AGEMA_signal_9317), .Z1_t (new_AGEMA_signal_9318), .Z1_f (new_AGEMA_signal_9319) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M24), .A0_f (new_AGEMA_signal_9581), .A1_t (new_AGEMA_signal_9582), .A1_f (new_AGEMA_signal_9583), .B0_t (SubBytesIns_Inst_Sbox_7_M34), .B0_f (new_AGEMA_signal_9317), .B1_t (new_AGEMA_signal_9318), .B1_f (new_AGEMA_signal_9319), .Z0_t (SubBytesIns_Inst_Sbox_7_M35), .Z0_f (new_AGEMA_signal_9890), .Z1_t (new_AGEMA_signal_9891), .Z1_f (new_AGEMA_signal_9892) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M24), .A0_f (new_AGEMA_signal_9581), .A1_t (new_AGEMA_signal_9582), .A1_f (new_AGEMA_signal_9583), .B0_t (SubBytesIns_Inst_Sbox_7_M25), .B0_f (new_AGEMA_signal_9311), .B1_t (new_AGEMA_signal_9312), .B1_f (new_AGEMA_signal_9313), .Z0_t (SubBytesIns_Inst_Sbox_7_M36), .Z0_f (new_AGEMA_signal_9893), .Z1_t (new_AGEMA_signal_9894), .Z1_f (new_AGEMA_signal_9895) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M21), .A0_f (new_AGEMA_signal_9074), .A1_t (new_AGEMA_signal_9075), .A1_f (new_AGEMA_signal_9076), .B0_t (SubBytesIns_Inst_Sbox_7_M29), .B0_f (new_AGEMA_signal_9881), .B1_t (new_AGEMA_signal_9882), .B1_f (new_AGEMA_signal_9883), .Z0_t (SubBytesIns_Inst_Sbox_7_M37), .Z0_f (new_AGEMA_signal_10148), .Z1_t (new_AGEMA_signal_10149), .Z1_f (new_AGEMA_signal_10150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M32), .A0_f (new_AGEMA_signal_9887), .A1_t (new_AGEMA_signal_9888), .A1_f (new_AGEMA_signal_9889), .B0_t (SubBytesIns_Inst_Sbox_7_M33), .B0_f (new_AGEMA_signal_9593), .B1_t (new_AGEMA_signal_9594), .B1_f (new_AGEMA_signal_9595), .Z0_t (SubBytesIns_Inst_Sbox_7_M38), .Z0_f (new_AGEMA_signal_10151), .Z1_t (new_AGEMA_signal_10152), .Z1_f (new_AGEMA_signal_10153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M23), .A0_f (new_AGEMA_signal_9308), .A1_t (new_AGEMA_signal_9309), .A1_f (new_AGEMA_signal_9310), .B0_t (SubBytesIns_Inst_Sbox_7_M30), .B0_f (new_AGEMA_signal_9884), .B1_t (new_AGEMA_signal_9885), .B1_f (new_AGEMA_signal_9886), .Z0_t (SubBytesIns_Inst_Sbox_7_M39), .Z0_f (new_AGEMA_signal_10154), .Z1_t (new_AGEMA_signal_10155), .Z1_f (new_AGEMA_signal_10156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M35), .A0_f (new_AGEMA_signal_9890), .A1_t (new_AGEMA_signal_9891), .A1_f (new_AGEMA_signal_9892), .B0_t (SubBytesIns_Inst_Sbox_7_M36), .B0_f (new_AGEMA_signal_9893), .B1_t (new_AGEMA_signal_9894), .B1_f (new_AGEMA_signal_9895), .Z0_t (SubBytesIns_Inst_Sbox_7_M40), .Z0_f (new_AGEMA_signal_10157), .Z1_t (new_AGEMA_signal_10158), .Z1_f (new_AGEMA_signal_10159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M38), .A0_f (new_AGEMA_signal_10151), .A1_t (new_AGEMA_signal_10152), .A1_f (new_AGEMA_signal_10153), .B0_t (SubBytesIns_Inst_Sbox_7_M40), .B0_f (new_AGEMA_signal_10157), .B1_t (new_AGEMA_signal_10158), .B1_f (new_AGEMA_signal_10159), .Z0_t (SubBytesIns_Inst_Sbox_7_M41), .Z0_f (new_AGEMA_signal_10652), .Z1_t (new_AGEMA_signal_10653), .Z1_f (new_AGEMA_signal_10654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M37), .A0_f (new_AGEMA_signal_10148), .A1_t (new_AGEMA_signal_10149), .A1_f (new_AGEMA_signal_10150), .B0_t (SubBytesIns_Inst_Sbox_7_M39), .B0_f (new_AGEMA_signal_10154), .B1_t (new_AGEMA_signal_10155), .B1_f (new_AGEMA_signal_10156), .Z0_t (SubBytesIns_Inst_Sbox_7_M42), .Z0_f (new_AGEMA_signal_10655), .Z1_t (new_AGEMA_signal_10656), .Z1_f (new_AGEMA_signal_10657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M37), .A0_f (new_AGEMA_signal_10148), .A1_t (new_AGEMA_signal_10149), .A1_f (new_AGEMA_signal_10150), .B0_t (SubBytesIns_Inst_Sbox_7_M38), .B0_f (new_AGEMA_signal_10151), .B1_t (new_AGEMA_signal_10152), .B1_f (new_AGEMA_signal_10153), .Z0_t (SubBytesIns_Inst_Sbox_7_M43), .Z0_f (new_AGEMA_signal_10658), .Z1_t (new_AGEMA_signal_10659), .Z1_f (new_AGEMA_signal_10660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M39), .A0_f (new_AGEMA_signal_10154), .A1_t (new_AGEMA_signal_10155), .A1_f (new_AGEMA_signal_10156), .B0_t (SubBytesIns_Inst_Sbox_7_M40), .B0_f (new_AGEMA_signal_10157), .B1_t (new_AGEMA_signal_10158), .B1_f (new_AGEMA_signal_10159), .Z0_t (SubBytesIns_Inst_Sbox_7_M44), .Z0_f (new_AGEMA_signal_10661), .Z1_t (new_AGEMA_signal_10662), .Z1_f (new_AGEMA_signal_10663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M42), .A0_f (new_AGEMA_signal_10655), .A1_t (new_AGEMA_signal_10656), .A1_f (new_AGEMA_signal_10657), .B0_t (SubBytesIns_Inst_Sbox_7_M41), .B0_f (new_AGEMA_signal_10652), .B1_t (new_AGEMA_signal_10653), .B1_f (new_AGEMA_signal_10654), .Z0_t (SubBytesIns_Inst_Sbox_7_M45), .Z0_f (new_AGEMA_signal_11372), .Z1_t (new_AGEMA_signal_11373), .Z1_f (new_AGEMA_signal_11374) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M44), .A0_f (new_AGEMA_signal_10661), .A1_t (new_AGEMA_signal_10662), .A1_f (new_AGEMA_signal_10663), .B0_t (SubBytesIns_Inst_Sbox_7_T6), .B0_f (new_AGEMA_signal_7096), .B1_t (new_AGEMA_signal_7097), .B1_f (new_AGEMA_signal_7098), .Z0_t (SubBytesIns_Inst_Sbox_7_M46), .Z0_f (new_AGEMA_signal_11375), .Z1_t (new_AGEMA_signal_11376), .Z1_f (new_AGEMA_signal_11377) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M40), .A0_f (new_AGEMA_signal_10157), .A1_t (new_AGEMA_signal_10158), .A1_f (new_AGEMA_signal_10159), .B0_t (SubBytesIns_Inst_Sbox_7_T8), .B0_f (new_AGEMA_signal_7745), .B1_t (new_AGEMA_signal_7746), .B1_f (new_AGEMA_signal_7747), .Z0_t (SubBytesIns_Inst_Sbox_7_M47), .Z0_f (new_AGEMA_signal_10664), .Z1_t (new_AGEMA_signal_10665), .Z1_f (new_AGEMA_signal_10666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M39), .A0_f (new_AGEMA_signal_10154), .A1_t (new_AGEMA_signal_10155), .A1_f (new_AGEMA_signal_10156), .B0_t (ciphertext_s0_t[56]), .B0_f (ciphertext_s0_f[56]), .B1_t (ciphertext_s1_t[56]), .B1_f (ciphertext_s1_f[56]), .Z0_t (SubBytesIns_Inst_Sbox_7_M48), .Z0_f (new_AGEMA_signal_10667), .Z1_t (new_AGEMA_signal_10668), .Z1_f (new_AGEMA_signal_10669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M43), .A0_f (new_AGEMA_signal_10658), .A1_t (new_AGEMA_signal_10659), .A1_f (new_AGEMA_signal_10660), .B0_t (SubBytesIns_Inst_Sbox_7_T16), .B0_f (new_AGEMA_signal_7108), .B1_t (new_AGEMA_signal_7109), .B1_f (new_AGEMA_signal_7110), .Z0_t (SubBytesIns_Inst_Sbox_7_M49), .Z0_f (new_AGEMA_signal_11378), .Z1_t (new_AGEMA_signal_11379), .Z1_f (new_AGEMA_signal_11380) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M38), .A0_f (new_AGEMA_signal_10151), .A1_t (new_AGEMA_signal_10152), .A1_f (new_AGEMA_signal_10153), .B0_t (SubBytesIns_Inst_Sbox_7_T9), .B0_f (new_AGEMA_signal_7099), .B1_t (new_AGEMA_signal_7100), .B1_f (new_AGEMA_signal_7101), .Z0_t (SubBytesIns_Inst_Sbox_7_M50), .Z0_f (new_AGEMA_signal_10670), .Z1_t (new_AGEMA_signal_10671), .Z1_f (new_AGEMA_signal_10672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M37), .A0_f (new_AGEMA_signal_10148), .A1_t (new_AGEMA_signal_10149), .A1_f (new_AGEMA_signal_10150), .B0_t (SubBytesIns_Inst_Sbox_7_T17), .B0_f (new_AGEMA_signal_7754), .B1_t (new_AGEMA_signal_7755), .B1_f (new_AGEMA_signal_7756), .Z0_t (SubBytesIns_Inst_Sbox_7_M51), .Z0_f (new_AGEMA_signal_10673), .Z1_t (new_AGEMA_signal_10674), .Z1_f (new_AGEMA_signal_10675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M42), .A0_f (new_AGEMA_signal_10655), .A1_t (new_AGEMA_signal_10656), .A1_f (new_AGEMA_signal_10657), .B0_t (SubBytesIns_Inst_Sbox_7_T15), .B0_f (new_AGEMA_signal_7105), .B1_t (new_AGEMA_signal_7106), .B1_f (new_AGEMA_signal_7107), .Z0_t (SubBytesIns_Inst_Sbox_7_M52), .Z0_f (new_AGEMA_signal_11381), .Z1_t (new_AGEMA_signal_11382), .Z1_f (new_AGEMA_signal_11383) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M45), .A0_f (new_AGEMA_signal_11372), .A1_t (new_AGEMA_signal_11373), .A1_f (new_AGEMA_signal_11374), .B0_t (SubBytesIns_Inst_Sbox_7_T27), .B0_f (new_AGEMA_signal_7117), .B1_t (new_AGEMA_signal_7118), .B1_f (new_AGEMA_signal_7119), .Z0_t (SubBytesIns_Inst_Sbox_7_M53), .Z0_f (new_AGEMA_signal_12026), .Z1_t (new_AGEMA_signal_12027), .Z1_f (new_AGEMA_signal_12028) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M41), .A0_f (new_AGEMA_signal_10652), .A1_t (new_AGEMA_signal_10653), .A1_f (new_AGEMA_signal_10654), .B0_t (SubBytesIns_Inst_Sbox_7_T10), .B0_f (new_AGEMA_signal_7748), .B1_t (new_AGEMA_signal_7749), .B1_f (new_AGEMA_signal_7750), .Z0_t (SubBytesIns_Inst_Sbox_7_M54), .Z0_f (new_AGEMA_signal_11384), .Z1_t (new_AGEMA_signal_11385), .Z1_f (new_AGEMA_signal_11386) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M44), .A0_f (new_AGEMA_signal_10661), .A1_t (new_AGEMA_signal_10662), .A1_f (new_AGEMA_signal_10663), .B0_t (SubBytesIns_Inst_Sbox_7_T13), .B0_f (new_AGEMA_signal_7102), .B1_t (new_AGEMA_signal_7103), .B1_f (new_AGEMA_signal_7104), .Z0_t (SubBytesIns_Inst_Sbox_7_M55), .Z0_f (new_AGEMA_signal_11387), .Z1_t (new_AGEMA_signal_11388), .Z1_f (new_AGEMA_signal_11389) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M40), .A0_f (new_AGEMA_signal_10157), .A1_t (new_AGEMA_signal_10158), .A1_f (new_AGEMA_signal_10159), .B0_t (SubBytesIns_Inst_Sbox_7_T23), .B0_f (new_AGEMA_signal_7760), .B1_t (new_AGEMA_signal_7761), .B1_f (new_AGEMA_signal_7762), .Z0_t (SubBytesIns_Inst_Sbox_7_M56), .Z0_f (new_AGEMA_signal_10676), .Z1_t (new_AGEMA_signal_10677), .Z1_f (new_AGEMA_signal_10678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M39), .A0_f (new_AGEMA_signal_10154), .A1_t (new_AGEMA_signal_10155), .A1_f (new_AGEMA_signal_10156), .B0_t (SubBytesIns_Inst_Sbox_7_T19), .B0_f (new_AGEMA_signal_7111), .B1_t (new_AGEMA_signal_7112), .B1_f (new_AGEMA_signal_7113), .Z0_t (SubBytesIns_Inst_Sbox_7_M57), .Z0_f (new_AGEMA_signal_10679), .Z1_t (new_AGEMA_signal_10680), .Z1_f (new_AGEMA_signal_10681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M43), .A0_f (new_AGEMA_signal_10658), .A1_t (new_AGEMA_signal_10659), .A1_f (new_AGEMA_signal_10660), .B0_t (SubBytesIns_Inst_Sbox_7_T3), .B0_f (new_AGEMA_signal_6562), .B1_t (new_AGEMA_signal_6563), .B1_f (new_AGEMA_signal_6564), .Z0_t (SubBytesIns_Inst_Sbox_7_M58), .Z0_f (new_AGEMA_signal_11390), .Z1_t (new_AGEMA_signal_11391), .Z1_f (new_AGEMA_signal_11392) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M38), .A0_f (new_AGEMA_signal_10151), .A1_t (new_AGEMA_signal_10152), .A1_f (new_AGEMA_signal_10153), .B0_t (SubBytesIns_Inst_Sbox_7_T22), .B0_f (new_AGEMA_signal_7114), .B1_t (new_AGEMA_signal_7115), .B1_f (new_AGEMA_signal_7116), .Z0_t (SubBytesIns_Inst_Sbox_7_M59), .Z0_f (new_AGEMA_signal_10682), .Z1_t (new_AGEMA_signal_10683), .Z1_f (new_AGEMA_signal_10684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M37), .A0_f (new_AGEMA_signal_10148), .A1_t (new_AGEMA_signal_10149), .A1_f (new_AGEMA_signal_10150), .B0_t (SubBytesIns_Inst_Sbox_7_T20), .B0_f (new_AGEMA_signal_7757), .B1_t (new_AGEMA_signal_7758), .B1_f (new_AGEMA_signal_7759), .Z0_t (SubBytesIns_Inst_Sbox_7_M60), .Z0_f (new_AGEMA_signal_10685), .Z1_t (new_AGEMA_signal_10686), .Z1_f (new_AGEMA_signal_10687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M42), .A0_f (new_AGEMA_signal_10655), .A1_t (new_AGEMA_signal_10656), .A1_f (new_AGEMA_signal_10657), .B0_t (SubBytesIns_Inst_Sbox_7_T1), .B0_f (new_AGEMA_signal_6556), .B1_t (new_AGEMA_signal_6557), .B1_f (new_AGEMA_signal_6558), .Z0_t (SubBytesIns_Inst_Sbox_7_M61), .Z0_f (new_AGEMA_signal_11393), .Z1_t (new_AGEMA_signal_11394), .Z1_f (new_AGEMA_signal_11395) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M45), .A0_f (new_AGEMA_signal_11372), .A1_t (new_AGEMA_signal_11373), .A1_f (new_AGEMA_signal_11374), .B0_t (SubBytesIns_Inst_Sbox_7_T4), .B0_f (new_AGEMA_signal_6565), .B1_t (new_AGEMA_signal_6566), .B1_f (new_AGEMA_signal_6567), .Z0_t (SubBytesIns_Inst_Sbox_7_M62), .Z0_f (new_AGEMA_signal_12029), .Z1_t (new_AGEMA_signal_12030), .Z1_f (new_AGEMA_signal_12031) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M41), .A0_f (new_AGEMA_signal_10652), .A1_t (new_AGEMA_signal_10653), .A1_f (new_AGEMA_signal_10654), .B0_t (SubBytesIns_Inst_Sbox_7_T2), .B0_f (new_AGEMA_signal_6559), .B1_t (new_AGEMA_signal_6560), .B1_f (new_AGEMA_signal_6561), .Z0_t (SubBytesIns_Inst_Sbox_7_M63), .Z0_f (new_AGEMA_signal_11396), .Z1_t (new_AGEMA_signal_11397), .Z1_f (new_AGEMA_signal_11398) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M61), .A0_f (new_AGEMA_signal_11393), .A1_t (new_AGEMA_signal_11394), .A1_f (new_AGEMA_signal_11395), .B0_t (SubBytesIns_Inst_Sbox_7_M62), .B0_f (new_AGEMA_signal_12029), .B1_t (new_AGEMA_signal_12030), .B1_f (new_AGEMA_signal_12031), .Z0_t (SubBytesIns_Inst_Sbox_7_L0), .Z0_f (new_AGEMA_signal_12593), .Z1_t (new_AGEMA_signal_12594), .Z1_f (new_AGEMA_signal_12595) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M50), .A0_f (new_AGEMA_signal_10670), .A1_t (new_AGEMA_signal_10671), .A1_f (new_AGEMA_signal_10672), .B0_t (SubBytesIns_Inst_Sbox_7_M56), .B0_f (new_AGEMA_signal_10676), .B1_t (new_AGEMA_signal_10677), .B1_f (new_AGEMA_signal_10678), .Z0_t (SubBytesIns_Inst_Sbox_7_L1), .Z0_f (new_AGEMA_signal_11399), .Z1_t (new_AGEMA_signal_11400), .Z1_f (new_AGEMA_signal_11401) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M46), .A0_f (new_AGEMA_signal_11375), .A1_t (new_AGEMA_signal_11376), .A1_f (new_AGEMA_signal_11377), .B0_t (SubBytesIns_Inst_Sbox_7_M48), .B0_f (new_AGEMA_signal_10667), .B1_t (new_AGEMA_signal_10668), .B1_f (new_AGEMA_signal_10669), .Z0_t (SubBytesIns_Inst_Sbox_7_L2), .Z0_f (new_AGEMA_signal_12032), .Z1_t (new_AGEMA_signal_12033), .Z1_f (new_AGEMA_signal_12034) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M47), .A0_f (new_AGEMA_signal_10664), .A1_t (new_AGEMA_signal_10665), .A1_f (new_AGEMA_signal_10666), .B0_t (SubBytesIns_Inst_Sbox_7_M55), .B0_f (new_AGEMA_signal_11387), .B1_t (new_AGEMA_signal_11388), .B1_f (new_AGEMA_signal_11389), .Z0_t (SubBytesIns_Inst_Sbox_7_L3), .Z0_f (new_AGEMA_signal_12035), .Z1_t (new_AGEMA_signal_12036), .Z1_f (new_AGEMA_signal_12037) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M54), .A0_f (new_AGEMA_signal_11384), .A1_t (new_AGEMA_signal_11385), .A1_f (new_AGEMA_signal_11386), .B0_t (SubBytesIns_Inst_Sbox_7_M58), .B0_f (new_AGEMA_signal_11390), .B1_t (new_AGEMA_signal_11391), .B1_f (new_AGEMA_signal_11392), .Z0_t (SubBytesIns_Inst_Sbox_7_L4), .Z0_f (new_AGEMA_signal_12038), .Z1_t (new_AGEMA_signal_12039), .Z1_f (new_AGEMA_signal_12040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M49), .A0_f (new_AGEMA_signal_11378), .A1_t (new_AGEMA_signal_11379), .A1_f (new_AGEMA_signal_11380), .B0_t (SubBytesIns_Inst_Sbox_7_M61), .B0_f (new_AGEMA_signal_11393), .B1_t (new_AGEMA_signal_11394), .B1_f (new_AGEMA_signal_11395), .Z0_t (SubBytesIns_Inst_Sbox_7_L5), .Z0_f (new_AGEMA_signal_12041), .Z1_t (new_AGEMA_signal_12042), .Z1_f (new_AGEMA_signal_12043) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M62), .A0_f (new_AGEMA_signal_12029), .A1_t (new_AGEMA_signal_12030), .A1_f (new_AGEMA_signal_12031), .B0_t (SubBytesIns_Inst_Sbox_7_L5), .B0_f (new_AGEMA_signal_12041), .B1_t (new_AGEMA_signal_12042), .B1_f (new_AGEMA_signal_12043), .Z0_t (SubBytesIns_Inst_Sbox_7_L6), .Z0_f (new_AGEMA_signal_12596), .Z1_t (new_AGEMA_signal_12597), .Z1_f (new_AGEMA_signal_12598) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M46), .A0_f (new_AGEMA_signal_11375), .A1_t (new_AGEMA_signal_11376), .A1_f (new_AGEMA_signal_11377), .B0_t (SubBytesIns_Inst_Sbox_7_L3), .B0_f (new_AGEMA_signal_12035), .B1_t (new_AGEMA_signal_12036), .B1_f (new_AGEMA_signal_12037), .Z0_t (SubBytesIns_Inst_Sbox_7_L7), .Z0_f (new_AGEMA_signal_12599), .Z1_t (new_AGEMA_signal_12600), .Z1_f (new_AGEMA_signal_12601) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M51), .A0_f (new_AGEMA_signal_10673), .A1_t (new_AGEMA_signal_10674), .A1_f (new_AGEMA_signal_10675), .B0_t (SubBytesIns_Inst_Sbox_7_M59), .B0_f (new_AGEMA_signal_10682), .B1_t (new_AGEMA_signal_10683), .B1_f (new_AGEMA_signal_10684), .Z0_t (SubBytesIns_Inst_Sbox_7_L8), .Z0_f (new_AGEMA_signal_11402), .Z1_t (new_AGEMA_signal_11403), .Z1_f (new_AGEMA_signal_11404) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M52), .A0_f (new_AGEMA_signal_11381), .A1_t (new_AGEMA_signal_11382), .A1_f (new_AGEMA_signal_11383), .B0_t (SubBytesIns_Inst_Sbox_7_M53), .B0_f (new_AGEMA_signal_12026), .B1_t (new_AGEMA_signal_12027), .B1_f (new_AGEMA_signal_12028), .Z0_t (SubBytesIns_Inst_Sbox_7_L9), .Z0_f (new_AGEMA_signal_12602), .Z1_t (new_AGEMA_signal_12603), .Z1_f (new_AGEMA_signal_12604) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M53), .A0_f (new_AGEMA_signal_12026), .A1_t (new_AGEMA_signal_12027), .A1_f (new_AGEMA_signal_12028), .B0_t (SubBytesIns_Inst_Sbox_7_L4), .B0_f (new_AGEMA_signal_12038), .B1_t (new_AGEMA_signal_12039), .B1_f (new_AGEMA_signal_12040), .Z0_t (SubBytesIns_Inst_Sbox_7_L10), .Z0_f (new_AGEMA_signal_12605), .Z1_t (new_AGEMA_signal_12606), .Z1_f (new_AGEMA_signal_12607) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M60), .A0_f (new_AGEMA_signal_10685), .A1_t (new_AGEMA_signal_10686), .A1_f (new_AGEMA_signal_10687), .B0_t (SubBytesIns_Inst_Sbox_7_L2), .B0_f (new_AGEMA_signal_12032), .B1_t (new_AGEMA_signal_12033), .B1_f (new_AGEMA_signal_12034), .Z0_t (SubBytesIns_Inst_Sbox_7_L11), .Z0_f (new_AGEMA_signal_12608), .Z1_t (new_AGEMA_signal_12609), .Z1_f (new_AGEMA_signal_12610) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M48), .A0_f (new_AGEMA_signal_10667), .A1_t (new_AGEMA_signal_10668), .A1_f (new_AGEMA_signal_10669), .B0_t (SubBytesIns_Inst_Sbox_7_M51), .B0_f (new_AGEMA_signal_10673), .B1_t (new_AGEMA_signal_10674), .B1_f (new_AGEMA_signal_10675), .Z0_t (SubBytesIns_Inst_Sbox_7_L12), .Z0_f (new_AGEMA_signal_11405), .Z1_t (new_AGEMA_signal_11406), .Z1_f (new_AGEMA_signal_11407) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M50), .A0_f (new_AGEMA_signal_10670), .A1_t (new_AGEMA_signal_10671), .A1_f (new_AGEMA_signal_10672), .B0_t (SubBytesIns_Inst_Sbox_7_L0), .B0_f (new_AGEMA_signal_12593), .B1_t (new_AGEMA_signal_12594), .B1_f (new_AGEMA_signal_12595), .Z0_t (SubBytesIns_Inst_Sbox_7_L13), .Z0_f (new_AGEMA_signal_13199), .Z1_t (new_AGEMA_signal_13200), .Z1_f (new_AGEMA_signal_13201) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M52), .A0_f (new_AGEMA_signal_11381), .A1_t (new_AGEMA_signal_11382), .A1_f (new_AGEMA_signal_11383), .B0_t (SubBytesIns_Inst_Sbox_7_M61), .B0_f (new_AGEMA_signal_11393), .B1_t (new_AGEMA_signal_11394), .B1_f (new_AGEMA_signal_11395), .Z0_t (SubBytesIns_Inst_Sbox_7_L14), .Z0_f (new_AGEMA_signal_12044), .Z1_t (new_AGEMA_signal_12045), .Z1_f (new_AGEMA_signal_12046) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M55), .A0_f (new_AGEMA_signal_11387), .A1_t (new_AGEMA_signal_11388), .A1_f (new_AGEMA_signal_11389), .B0_t (SubBytesIns_Inst_Sbox_7_L1), .B0_f (new_AGEMA_signal_11399), .B1_t (new_AGEMA_signal_11400), .B1_f (new_AGEMA_signal_11401), .Z0_t (SubBytesIns_Inst_Sbox_7_L15), .Z0_f (new_AGEMA_signal_12047), .Z1_t (new_AGEMA_signal_12048), .Z1_f (new_AGEMA_signal_12049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M56), .A0_f (new_AGEMA_signal_10676), .A1_t (new_AGEMA_signal_10677), .A1_f (new_AGEMA_signal_10678), .B0_t (SubBytesIns_Inst_Sbox_7_L0), .B0_f (new_AGEMA_signal_12593), .B1_t (new_AGEMA_signal_12594), .B1_f (new_AGEMA_signal_12595), .Z0_t (SubBytesIns_Inst_Sbox_7_L16), .Z0_f (new_AGEMA_signal_13202), .Z1_t (new_AGEMA_signal_13203), .Z1_f (new_AGEMA_signal_13204) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M57), .A0_f (new_AGEMA_signal_10679), .A1_t (new_AGEMA_signal_10680), .A1_f (new_AGEMA_signal_10681), .B0_t (SubBytesIns_Inst_Sbox_7_L1), .B0_f (new_AGEMA_signal_11399), .B1_t (new_AGEMA_signal_11400), .B1_f (new_AGEMA_signal_11401), .Z0_t (SubBytesIns_Inst_Sbox_7_L17), .Z0_f (new_AGEMA_signal_12050), .Z1_t (new_AGEMA_signal_12051), .Z1_f (new_AGEMA_signal_12052) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M58), .A0_f (new_AGEMA_signal_11390), .A1_t (new_AGEMA_signal_11391), .A1_f (new_AGEMA_signal_11392), .B0_t (SubBytesIns_Inst_Sbox_7_L8), .B0_f (new_AGEMA_signal_11402), .B1_t (new_AGEMA_signal_11403), .B1_f (new_AGEMA_signal_11404), .Z0_t (SubBytesIns_Inst_Sbox_7_L18), .Z0_f (new_AGEMA_signal_12053), .Z1_t (new_AGEMA_signal_12054), .Z1_f (new_AGEMA_signal_12055) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M63), .A0_f (new_AGEMA_signal_11396), .A1_t (new_AGEMA_signal_11397), .A1_f (new_AGEMA_signal_11398), .B0_t (SubBytesIns_Inst_Sbox_7_L4), .B0_f (new_AGEMA_signal_12038), .B1_t (new_AGEMA_signal_12039), .B1_f (new_AGEMA_signal_12040), .Z0_t (SubBytesIns_Inst_Sbox_7_L19), .Z0_f (new_AGEMA_signal_12611), .Z1_t (new_AGEMA_signal_12612), .Z1_f (new_AGEMA_signal_12613) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L0), .A0_f (new_AGEMA_signal_12593), .A1_t (new_AGEMA_signal_12594), .A1_f (new_AGEMA_signal_12595), .B0_t (SubBytesIns_Inst_Sbox_7_L1), .B0_f (new_AGEMA_signal_11399), .B1_t (new_AGEMA_signal_11400), .B1_f (new_AGEMA_signal_11401), .Z0_t (SubBytesIns_Inst_Sbox_7_L20), .Z0_f (new_AGEMA_signal_13205), .Z1_t (new_AGEMA_signal_13206), .Z1_f (new_AGEMA_signal_13207) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L1), .A0_f (new_AGEMA_signal_11399), .A1_t (new_AGEMA_signal_11400), .A1_f (new_AGEMA_signal_11401), .B0_t (SubBytesIns_Inst_Sbox_7_L7), .B0_f (new_AGEMA_signal_12599), .B1_t (new_AGEMA_signal_12600), .B1_f (new_AGEMA_signal_12601), .Z0_t (SubBytesIns_Inst_Sbox_7_L21), .Z0_f (new_AGEMA_signal_13208), .Z1_t (new_AGEMA_signal_13209), .Z1_f (new_AGEMA_signal_13210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L3), .A0_f (new_AGEMA_signal_12035), .A1_t (new_AGEMA_signal_12036), .A1_f (new_AGEMA_signal_12037), .B0_t (SubBytesIns_Inst_Sbox_7_L12), .B0_f (new_AGEMA_signal_11405), .B1_t (new_AGEMA_signal_11406), .B1_f (new_AGEMA_signal_11407), .Z0_t (SubBytesIns_Inst_Sbox_7_L22), .Z0_f (new_AGEMA_signal_12614), .Z1_t (new_AGEMA_signal_12615), .Z1_f (new_AGEMA_signal_12616) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L18), .A0_f (new_AGEMA_signal_12053), .A1_t (new_AGEMA_signal_12054), .A1_f (new_AGEMA_signal_12055), .B0_t (SubBytesIns_Inst_Sbox_7_L2), .B0_f (new_AGEMA_signal_12032), .B1_t (new_AGEMA_signal_12033), .B1_f (new_AGEMA_signal_12034), .Z0_t (SubBytesIns_Inst_Sbox_7_L23), .Z0_f (new_AGEMA_signal_12617), .Z1_t (new_AGEMA_signal_12618), .Z1_f (new_AGEMA_signal_12619) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L15), .A0_f (new_AGEMA_signal_12047), .A1_t (new_AGEMA_signal_12048), .A1_f (new_AGEMA_signal_12049), .B0_t (SubBytesIns_Inst_Sbox_7_L9), .B0_f (new_AGEMA_signal_12602), .B1_t (new_AGEMA_signal_12603), .B1_f (new_AGEMA_signal_12604), .Z0_t (SubBytesIns_Inst_Sbox_7_L24), .Z0_f (new_AGEMA_signal_13211), .Z1_t (new_AGEMA_signal_13212), .Z1_f (new_AGEMA_signal_13213) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L6), .A0_f (new_AGEMA_signal_12596), .A1_t (new_AGEMA_signal_12597), .A1_f (new_AGEMA_signal_12598), .B0_t (SubBytesIns_Inst_Sbox_7_L10), .B0_f (new_AGEMA_signal_12605), .B1_t (new_AGEMA_signal_12606), .B1_f (new_AGEMA_signal_12607), .Z0_t (SubBytesIns_Inst_Sbox_7_L25), .Z0_f (new_AGEMA_signal_13214), .Z1_t (new_AGEMA_signal_13215), .Z1_f (new_AGEMA_signal_13216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L7), .A0_f (new_AGEMA_signal_12599), .A1_t (new_AGEMA_signal_12600), .A1_f (new_AGEMA_signal_12601), .B0_t (SubBytesIns_Inst_Sbox_7_L9), .B0_f (new_AGEMA_signal_12602), .B1_t (new_AGEMA_signal_12603), .B1_f (new_AGEMA_signal_12604), .Z0_t (SubBytesIns_Inst_Sbox_7_L26), .Z0_f (new_AGEMA_signal_13217), .Z1_t (new_AGEMA_signal_13218), .Z1_f (new_AGEMA_signal_13219) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L8), .A0_f (new_AGEMA_signal_11402), .A1_t (new_AGEMA_signal_11403), .A1_f (new_AGEMA_signal_11404), .B0_t (SubBytesIns_Inst_Sbox_7_L10), .B0_f (new_AGEMA_signal_12605), .B1_t (new_AGEMA_signal_12606), .B1_f (new_AGEMA_signal_12607), .Z0_t (SubBytesIns_Inst_Sbox_7_L27), .Z0_f (new_AGEMA_signal_13220), .Z1_t (new_AGEMA_signal_13221), .Z1_f (new_AGEMA_signal_13222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L11), .A0_f (new_AGEMA_signal_12608), .A1_t (new_AGEMA_signal_12609), .A1_f (new_AGEMA_signal_12610), .B0_t (SubBytesIns_Inst_Sbox_7_L14), .B0_f (new_AGEMA_signal_12044), .B1_t (new_AGEMA_signal_12045), .B1_f (new_AGEMA_signal_12046), .Z0_t (SubBytesIns_Inst_Sbox_7_L28), .Z0_f (new_AGEMA_signal_13223), .Z1_t (new_AGEMA_signal_13224), .Z1_f (new_AGEMA_signal_13225) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L11), .A0_f (new_AGEMA_signal_12608), .A1_t (new_AGEMA_signal_12609), .A1_f (new_AGEMA_signal_12610), .B0_t (SubBytesIns_Inst_Sbox_7_L17), .B0_f (new_AGEMA_signal_12050), .B1_t (new_AGEMA_signal_12051), .B1_f (new_AGEMA_signal_12052), .Z0_t (SubBytesIns_Inst_Sbox_7_L29), .Z0_f (new_AGEMA_signal_13226), .Z1_t (new_AGEMA_signal_13227), .Z1_f (new_AGEMA_signal_13228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L6), .A0_f (new_AGEMA_signal_12596), .A1_t (new_AGEMA_signal_12597), .A1_f (new_AGEMA_signal_12598), .B0_t (SubBytesIns_Inst_Sbox_7_L24), .B0_f (new_AGEMA_signal_13211), .B1_t (new_AGEMA_signal_13212), .B1_f (new_AGEMA_signal_13213), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .Z0_f (new_AGEMA_signal_13787), .Z1_t (new_AGEMA_signal_13788), .Z1_f (new_AGEMA_signal_13789) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L16), .A0_f (new_AGEMA_signal_13202), .A1_t (new_AGEMA_signal_13203), .A1_f (new_AGEMA_signal_13204), .B0_t (SubBytesIns_Inst_Sbox_7_L26), .B0_f (new_AGEMA_signal_13217), .B1_t (new_AGEMA_signal_13218), .B1_f (new_AGEMA_signal_13219), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .Z0_f (new_AGEMA_signal_13790), .Z1_t (new_AGEMA_signal_13791), .Z1_f (new_AGEMA_signal_13792) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L19), .A0_f (new_AGEMA_signal_12611), .A1_t (new_AGEMA_signal_12612), .A1_f (new_AGEMA_signal_12613), .B0_t (SubBytesIns_Inst_Sbox_7_L28), .B0_f (new_AGEMA_signal_13223), .B1_t (new_AGEMA_signal_13224), .B1_f (new_AGEMA_signal_13225), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .Z0_f (new_AGEMA_signal_13793), .Z1_t (new_AGEMA_signal_13794), .Z1_f (new_AGEMA_signal_13795) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L6), .A0_f (new_AGEMA_signal_12596), .A1_t (new_AGEMA_signal_12597), .A1_f (new_AGEMA_signal_12598), .B0_t (SubBytesIns_Inst_Sbox_7_L21), .B0_f (new_AGEMA_signal_13208), .B1_t (new_AGEMA_signal_13209), .B1_f (new_AGEMA_signal_13210), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .Z0_f (new_AGEMA_signal_13796), .Z1_t (new_AGEMA_signal_13797), .Z1_f (new_AGEMA_signal_13798) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L20), .A0_f (new_AGEMA_signal_13205), .A1_t (new_AGEMA_signal_13206), .A1_f (new_AGEMA_signal_13207), .B0_t (SubBytesIns_Inst_Sbox_7_L22), .B0_f (new_AGEMA_signal_12614), .B1_t (new_AGEMA_signal_12615), .B1_f (new_AGEMA_signal_12616), .Z0_t (MixColumnsInput[59]), .Z0_f (new_AGEMA_signal_13799), .Z1_t (new_AGEMA_signal_13800), .Z1_f (new_AGEMA_signal_13801) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L25), .A0_f (new_AGEMA_signal_13214), .A1_t (new_AGEMA_signal_13215), .A1_f (new_AGEMA_signal_13216), .B0_t (SubBytesIns_Inst_Sbox_7_L29), .B0_f (new_AGEMA_signal_13226), .B1_t (new_AGEMA_signal_13227), .B1_f (new_AGEMA_signal_13228), .Z0_t (MixColumnsInput[58]), .Z0_f (new_AGEMA_signal_13802), .Z1_t (new_AGEMA_signal_13803), .Z1_f (new_AGEMA_signal_13804) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L13), .A0_f (new_AGEMA_signal_13199), .A1_t (new_AGEMA_signal_13200), .A1_f (new_AGEMA_signal_13201), .B0_t (SubBytesIns_Inst_Sbox_7_L27), .B0_f (new_AGEMA_signal_13220), .B1_t (new_AGEMA_signal_13221), .B1_f (new_AGEMA_signal_13222), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .Z0_f (new_AGEMA_signal_13805), .Z1_t (new_AGEMA_signal_13806), .Z1_f (new_AGEMA_signal_13807) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L6), .A0_f (new_AGEMA_signal_12596), .A1_t (new_AGEMA_signal_12597), .A1_f (new_AGEMA_signal_12598), .B0_t (SubBytesIns_Inst_Sbox_7_L23), .B0_f (new_AGEMA_signal_12617), .B1_t (new_AGEMA_signal_12618), .B1_f (new_AGEMA_signal_12619), .Z0_t (MixColumnsInput[56]), .Z0_f (new_AGEMA_signal_13229), .Z1_t (new_AGEMA_signal_13230), .Z1_f (new_AGEMA_signal_13231) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[71]), .A0_f (ciphertext_s0_f[71]), .A1_t (ciphertext_s1_t[71]), .A1_f (ciphertext_s1_f[71]), .B0_t (ciphertext_s0_t[68]), .B0_f (ciphertext_s0_f[68]), .B1_t (ciphertext_s1_t[68]), .B1_f (ciphertext_s1_f[68]), .Z0_t (SubBytesIns_Inst_Sbox_8_T1), .Z0_f (new_AGEMA_signal_6586), .Z1_t (new_AGEMA_signal_6587), .Z1_f (new_AGEMA_signal_6588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[71]), .A0_f (ciphertext_s0_f[71]), .A1_t (ciphertext_s1_t[71]), .A1_f (ciphertext_s1_f[71]), .B0_t (ciphertext_s0_t[66]), .B0_f (ciphertext_s0_f[66]), .B1_t (ciphertext_s1_t[66]), .B1_f (ciphertext_s1_f[66]), .Z0_t (SubBytesIns_Inst_Sbox_8_T2), .Z0_f (new_AGEMA_signal_6589), .Z1_t (new_AGEMA_signal_6590), .Z1_f (new_AGEMA_signal_6591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[71]), .A0_f (ciphertext_s0_f[71]), .A1_t (ciphertext_s1_t[71]), .A1_f (ciphertext_s1_f[71]), .B0_t (ciphertext_s0_t[65]), .B0_f (ciphertext_s0_f[65]), .B1_t (ciphertext_s1_t[65]), .B1_f (ciphertext_s1_f[65]), .Z0_t (SubBytesIns_Inst_Sbox_8_T3), .Z0_f (new_AGEMA_signal_6592), .Z1_t (new_AGEMA_signal_6593), .Z1_f (new_AGEMA_signal_6594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[68]), .A0_f (ciphertext_s0_f[68]), .A1_t (ciphertext_s1_t[68]), .A1_f (ciphertext_s1_f[68]), .B0_t (ciphertext_s0_t[66]), .B0_f (ciphertext_s0_f[66]), .B1_t (ciphertext_s1_t[66]), .B1_f (ciphertext_s1_f[66]), .Z0_t (SubBytesIns_Inst_Sbox_8_T4), .Z0_f (new_AGEMA_signal_6595), .Z1_t (new_AGEMA_signal_6596), .Z1_f (new_AGEMA_signal_6597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[67]), .A0_f (ciphertext_s0_f[67]), .A1_t (ciphertext_s1_t[67]), .A1_f (ciphertext_s1_f[67]), .B0_t (ciphertext_s0_t[65]), .B0_f (ciphertext_s0_f[65]), .B1_t (ciphertext_s1_t[65]), .B1_f (ciphertext_s1_f[65]), .Z0_t (SubBytesIns_Inst_Sbox_8_T5), .Z0_f (new_AGEMA_signal_6598), .Z1_t (new_AGEMA_signal_6599), .Z1_f (new_AGEMA_signal_6600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T1), .A0_f (new_AGEMA_signal_6586), .A1_t (new_AGEMA_signal_6587), .A1_f (new_AGEMA_signal_6588), .B0_t (SubBytesIns_Inst_Sbox_8_T5), .B0_f (new_AGEMA_signal_6598), .B1_t (new_AGEMA_signal_6599), .B1_f (new_AGEMA_signal_6600), .Z0_t (SubBytesIns_Inst_Sbox_8_T6), .Z0_f (new_AGEMA_signal_7120), .Z1_t (new_AGEMA_signal_7121), .Z1_f (new_AGEMA_signal_7122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[70]), .A0_f (ciphertext_s0_f[70]), .A1_t (ciphertext_s1_t[70]), .A1_f (ciphertext_s1_f[70]), .B0_t (ciphertext_s0_t[69]), .B0_f (ciphertext_s0_f[69]), .B1_t (ciphertext_s1_t[69]), .B1_f (ciphertext_s1_f[69]), .Z0_t (SubBytesIns_Inst_Sbox_8_T7), .Z0_f (new_AGEMA_signal_6601), .Z1_t (new_AGEMA_signal_6602), .Z1_f (new_AGEMA_signal_6603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[64]), .A0_f (ciphertext_s0_f[64]), .A1_t (ciphertext_s1_t[64]), .A1_f (ciphertext_s1_f[64]), .B0_t (SubBytesIns_Inst_Sbox_8_T6), .B0_f (new_AGEMA_signal_7120), .B1_t (new_AGEMA_signal_7121), .B1_f (new_AGEMA_signal_7122), .Z0_t (SubBytesIns_Inst_Sbox_8_T8), .Z0_f (new_AGEMA_signal_7784), .Z1_t (new_AGEMA_signal_7785), .Z1_f (new_AGEMA_signal_7786) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[64]), .A0_f (ciphertext_s0_f[64]), .A1_t (ciphertext_s1_t[64]), .A1_f (ciphertext_s1_f[64]), .B0_t (SubBytesIns_Inst_Sbox_8_T7), .B0_f (new_AGEMA_signal_6601), .B1_t (new_AGEMA_signal_6602), .B1_f (new_AGEMA_signal_6603), .Z0_t (SubBytesIns_Inst_Sbox_8_T9), .Z0_f (new_AGEMA_signal_7123), .Z1_t (new_AGEMA_signal_7124), .Z1_f (new_AGEMA_signal_7125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T6), .A0_f (new_AGEMA_signal_7120), .A1_t (new_AGEMA_signal_7121), .A1_f (new_AGEMA_signal_7122), .B0_t (SubBytesIns_Inst_Sbox_8_T7), .B0_f (new_AGEMA_signal_6601), .B1_t (new_AGEMA_signal_6602), .B1_f (new_AGEMA_signal_6603), .Z0_t (SubBytesIns_Inst_Sbox_8_T10), .Z0_f (new_AGEMA_signal_7787), .Z1_t (new_AGEMA_signal_7788), .Z1_f (new_AGEMA_signal_7789) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[70]), .A0_f (ciphertext_s0_f[70]), .A1_t (ciphertext_s1_t[70]), .A1_f (ciphertext_s1_f[70]), .B0_t (ciphertext_s0_t[66]), .B0_f (ciphertext_s0_f[66]), .B1_t (ciphertext_s1_t[66]), .B1_f (ciphertext_s1_f[66]), .Z0_t (SubBytesIns_Inst_Sbox_8_T11), .Z0_f (new_AGEMA_signal_6604), .Z1_t (new_AGEMA_signal_6605), .Z1_f (new_AGEMA_signal_6606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[69]), .A0_f (ciphertext_s0_f[69]), .A1_t (ciphertext_s1_t[69]), .A1_f (ciphertext_s1_f[69]), .B0_t (ciphertext_s0_t[66]), .B0_f (ciphertext_s0_f[66]), .B1_t (ciphertext_s1_t[66]), .B1_f (ciphertext_s1_f[66]), .Z0_t (SubBytesIns_Inst_Sbox_8_T12), .Z0_f (new_AGEMA_signal_6607), .Z1_t (new_AGEMA_signal_6608), .Z1_f (new_AGEMA_signal_6609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T3), .A0_f (new_AGEMA_signal_6592), .A1_t (new_AGEMA_signal_6593), .A1_f (new_AGEMA_signal_6594), .B0_t (SubBytesIns_Inst_Sbox_8_T4), .B0_f (new_AGEMA_signal_6595), .B1_t (new_AGEMA_signal_6596), .B1_f (new_AGEMA_signal_6597), .Z0_t (SubBytesIns_Inst_Sbox_8_T13), .Z0_f (new_AGEMA_signal_7126), .Z1_t (new_AGEMA_signal_7127), .Z1_f (new_AGEMA_signal_7128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T6), .A0_f (new_AGEMA_signal_7120), .A1_t (new_AGEMA_signal_7121), .A1_f (new_AGEMA_signal_7122), .B0_t (SubBytesIns_Inst_Sbox_8_T11), .B0_f (new_AGEMA_signal_6604), .B1_t (new_AGEMA_signal_6605), .B1_f (new_AGEMA_signal_6606), .Z0_t (SubBytesIns_Inst_Sbox_8_T14), .Z0_f (new_AGEMA_signal_7790), .Z1_t (new_AGEMA_signal_7791), .Z1_f (new_AGEMA_signal_7792) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T5), .A0_f (new_AGEMA_signal_6598), .A1_t (new_AGEMA_signal_6599), .A1_f (new_AGEMA_signal_6600), .B0_t (SubBytesIns_Inst_Sbox_8_T11), .B0_f (new_AGEMA_signal_6604), .B1_t (new_AGEMA_signal_6605), .B1_f (new_AGEMA_signal_6606), .Z0_t (SubBytesIns_Inst_Sbox_8_T15), .Z0_f (new_AGEMA_signal_7129), .Z1_t (new_AGEMA_signal_7130), .Z1_f (new_AGEMA_signal_7131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T5), .A0_f (new_AGEMA_signal_6598), .A1_t (new_AGEMA_signal_6599), .A1_f (new_AGEMA_signal_6600), .B0_t (SubBytesIns_Inst_Sbox_8_T12), .B0_f (new_AGEMA_signal_6607), .B1_t (new_AGEMA_signal_6608), .B1_f (new_AGEMA_signal_6609), .Z0_t (SubBytesIns_Inst_Sbox_8_T16), .Z0_f (new_AGEMA_signal_7132), .Z1_t (new_AGEMA_signal_7133), .Z1_f (new_AGEMA_signal_7134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T9), .A0_f (new_AGEMA_signal_7123), .A1_t (new_AGEMA_signal_7124), .A1_f (new_AGEMA_signal_7125), .B0_t (SubBytesIns_Inst_Sbox_8_T16), .B0_f (new_AGEMA_signal_7132), .B1_t (new_AGEMA_signal_7133), .B1_f (new_AGEMA_signal_7134), .Z0_t (SubBytesIns_Inst_Sbox_8_T17), .Z0_f (new_AGEMA_signal_7793), .Z1_t (new_AGEMA_signal_7794), .Z1_f (new_AGEMA_signal_7795) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[68]), .A0_f (ciphertext_s0_f[68]), .A1_t (ciphertext_s1_t[68]), .A1_f (ciphertext_s1_f[68]), .B0_t (ciphertext_s0_t[64]), .B0_f (ciphertext_s0_f[64]), .B1_t (ciphertext_s1_t[64]), .B1_f (ciphertext_s1_f[64]), .Z0_t (SubBytesIns_Inst_Sbox_8_T18), .Z0_f (new_AGEMA_signal_6610), .Z1_t (new_AGEMA_signal_6611), .Z1_f (new_AGEMA_signal_6612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T7), .A0_f (new_AGEMA_signal_6601), .A1_t (new_AGEMA_signal_6602), .A1_f (new_AGEMA_signal_6603), .B0_t (SubBytesIns_Inst_Sbox_8_T18), .B0_f (new_AGEMA_signal_6610), .B1_t (new_AGEMA_signal_6611), .B1_f (new_AGEMA_signal_6612), .Z0_t (SubBytesIns_Inst_Sbox_8_T19), .Z0_f (new_AGEMA_signal_7135), .Z1_t (new_AGEMA_signal_7136), .Z1_f (new_AGEMA_signal_7137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T1), .A0_f (new_AGEMA_signal_6586), .A1_t (new_AGEMA_signal_6587), .A1_f (new_AGEMA_signal_6588), .B0_t (SubBytesIns_Inst_Sbox_8_T19), .B0_f (new_AGEMA_signal_7135), .B1_t (new_AGEMA_signal_7136), .B1_f (new_AGEMA_signal_7137), .Z0_t (SubBytesIns_Inst_Sbox_8_T20), .Z0_f (new_AGEMA_signal_7796), .Z1_t (new_AGEMA_signal_7797), .Z1_f (new_AGEMA_signal_7798) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[65]), .A0_f (ciphertext_s0_f[65]), .A1_t (ciphertext_s1_t[65]), .A1_f (ciphertext_s1_f[65]), .B0_t (ciphertext_s0_t[64]), .B0_f (ciphertext_s0_f[64]), .B1_t (ciphertext_s1_t[64]), .B1_f (ciphertext_s1_f[64]), .Z0_t (SubBytesIns_Inst_Sbox_8_T21), .Z0_f (new_AGEMA_signal_6613), .Z1_t (new_AGEMA_signal_6614), .Z1_f (new_AGEMA_signal_6615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T7), .A0_f (new_AGEMA_signal_6601), .A1_t (new_AGEMA_signal_6602), .A1_f (new_AGEMA_signal_6603), .B0_t (SubBytesIns_Inst_Sbox_8_T21), .B0_f (new_AGEMA_signal_6613), .B1_t (new_AGEMA_signal_6614), .B1_f (new_AGEMA_signal_6615), .Z0_t (SubBytesIns_Inst_Sbox_8_T22), .Z0_f (new_AGEMA_signal_7138), .Z1_t (new_AGEMA_signal_7139), .Z1_f (new_AGEMA_signal_7140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T2), .A0_f (new_AGEMA_signal_6589), .A1_t (new_AGEMA_signal_6590), .A1_f (new_AGEMA_signal_6591), .B0_t (SubBytesIns_Inst_Sbox_8_T22), .B0_f (new_AGEMA_signal_7138), .B1_t (new_AGEMA_signal_7139), .B1_f (new_AGEMA_signal_7140), .Z0_t (SubBytesIns_Inst_Sbox_8_T23), .Z0_f (new_AGEMA_signal_7799), .Z1_t (new_AGEMA_signal_7800), .Z1_f (new_AGEMA_signal_7801) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T2), .A0_f (new_AGEMA_signal_6589), .A1_t (new_AGEMA_signal_6590), .A1_f (new_AGEMA_signal_6591), .B0_t (SubBytesIns_Inst_Sbox_8_T10), .B0_f (new_AGEMA_signal_7787), .B1_t (new_AGEMA_signal_7788), .B1_f (new_AGEMA_signal_7789), .Z0_t (SubBytesIns_Inst_Sbox_8_T24), .Z0_f (new_AGEMA_signal_8420), .Z1_t (new_AGEMA_signal_8421), .Z1_f (new_AGEMA_signal_8422) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T20), .A0_f (new_AGEMA_signal_7796), .A1_t (new_AGEMA_signal_7797), .A1_f (new_AGEMA_signal_7798), .B0_t (SubBytesIns_Inst_Sbox_8_T17), .B0_f (new_AGEMA_signal_7793), .B1_t (new_AGEMA_signal_7794), .B1_f (new_AGEMA_signal_7795), .Z0_t (SubBytesIns_Inst_Sbox_8_T25), .Z0_f (new_AGEMA_signal_8423), .Z1_t (new_AGEMA_signal_8424), .Z1_f (new_AGEMA_signal_8425) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T3), .A0_f (new_AGEMA_signal_6592), .A1_t (new_AGEMA_signal_6593), .A1_f (new_AGEMA_signal_6594), .B0_t (SubBytesIns_Inst_Sbox_8_T16), .B0_f (new_AGEMA_signal_7132), .B1_t (new_AGEMA_signal_7133), .B1_f (new_AGEMA_signal_7134), .Z0_t (SubBytesIns_Inst_Sbox_8_T26), .Z0_f (new_AGEMA_signal_7802), .Z1_t (new_AGEMA_signal_7803), .Z1_f (new_AGEMA_signal_7804) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T1), .A0_f (new_AGEMA_signal_6586), .A1_t (new_AGEMA_signal_6587), .A1_f (new_AGEMA_signal_6588), .B0_t (SubBytesIns_Inst_Sbox_8_T12), .B0_f (new_AGEMA_signal_6607), .B1_t (new_AGEMA_signal_6608), .B1_f (new_AGEMA_signal_6609), .Z0_t (SubBytesIns_Inst_Sbox_8_T27), .Z0_f (new_AGEMA_signal_7141), .Z1_t (new_AGEMA_signal_7142), .Z1_f (new_AGEMA_signal_7143) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T13), .A0_f (new_AGEMA_signal_7126), .A1_t (new_AGEMA_signal_7127), .A1_f (new_AGEMA_signal_7128), .B0_t (SubBytesIns_Inst_Sbox_8_T6), .B0_f (new_AGEMA_signal_7120), .B1_t (new_AGEMA_signal_7121), .B1_f (new_AGEMA_signal_7122), .Z0_t (SubBytesIns_Inst_Sbox_8_M1), .Z0_f (new_AGEMA_signal_7805), .Z1_t (new_AGEMA_signal_7806), .Z1_f (new_AGEMA_signal_7807) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T23), .A0_f (new_AGEMA_signal_7799), .A1_t (new_AGEMA_signal_7800), .A1_f (new_AGEMA_signal_7801), .B0_t (SubBytesIns_Inst_Sbox_8_T8), .B0_f (new_AGEMA_signal_7784), .B1_t (new_AGEMA_signal_7785), .B1_f (new_AGEMA_signal_7786), .Z0_t (SubBytesIns_Inst_Sbox_8_M2), .Z0_f (new_AGEMA_signal_8426), .Z1_t (new_AGEMA_signal_8427), .Z1_f (new_AGEMA_signal_8428) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T14), .A0_f (new_AGEMA_signal_7790), .A1_t (new_AGEMA_signal_7791), .A1_f (new_AGEMA_signal_7792), .B0_t (SubBytesIns_Inst_Sbox_8_M1), .B0_f (new_AGEMA_signal_7805), .B1_t (new_AGEMA_signal_7806), .B1_f (new_AGEMA_signal_7807), .Z0_t (SubBytesIns_Inst_Sbox_8_M3), .Z0_f (new_AGEMA_signal_8429), .Z1_t (new_AGEMA_signal_8430), .Z1_f (new_AGEMA_signal_8431) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T19), .A0_f (new_AGEMA_signal_7135), .A1_t (new_AGEMA_signal_7136), .A1_f (new_AGEMA_signal_7137), .B0_t (ciphertext_s0_t[64]), .B0_f (ciphertext_s0_f[64]), .B1_t (ciphertext_s1_t[64]), .B1_f (ciphertext_s1_f[64]), .Z0_t (SubBytesIns_Inst_Sbox_8_M4), .Z0_f (new_AGEMA_signal_7808), .Z1_t (new_AGEMA_signal_7809), .Z1_f (new_AGEMA_signal_7810) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M4), .A0_f (new_AGEMA_signal_7808), .A1_t (new_AGEMA_signal_7809), .A1_f (new_AGEMA_signal_7810), .B0_t (SubBytesIns_Inst_Sbox_8_M1), .B0_f (new_AGEMA_signal_7805), .B1_t (new_AGEMA_signal_7806), .B1_f (new_AGEMA_signal_7807), .Z0_t (SubBytesIns_Inst_Sbox_8_M5), .Z0_f (new_AGEMA_signal_8432), .Z1_t (new_AGEMA_signal_8433), .Z1_f (new_AGEMA_signal_8434) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T3), .A0_f (new_AGEMA_signal_6592), .A1_t (new_AGEMA_signal_6593), .A1_f (new_AGEMA_signal_6594), .B0_t (SubBytesIns_Inst_Sbox_8_T16), .B0_f (new_AGEMA_signal_7132), .B1_t (new_AGEMA_signal_7133), .B1_f (new_AGEMA_signal_7134), .Z0_t (SubBytesIns_Inst_Sbox_8_M6), .Z0_f (new_AGEMA_signal_7811), .Z1_t (new_AGEMA_signal_7812), .Z1_f (new_AGEMA_signal_7813) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T22), .A0_f (new_AGEMA_signal_7138), .A1_t (new_AGEMA_signal_7139), .A1_f (new_AGEMA_signal_7140), .B0_t (SubBytesIns_Inst_Sbox_8_T9), .B0_f (new_AGEMA_signal_7123), .B1_t (new_AGEMA_signal_7124), .B1_f (new_AGEMA_signal_7125), .Z0_t (SubBytesIns_Inst_Sbox_8_M7), .Z0_f (new_AGEMA_signal_7814), .Z1_t (new_AGEMA_signal_7815), .Z1_f (new_AGEMA_signal_7816) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T26), .A0_f (new_AGEMA_signal_7802), .A1_t (new_AGEMA_signal_7803), .A1_f (new_AGEMA_signal_7804), .B0_t (SubBytesIns_Inst_Sbox_8_M6), .B0_f (new_AGEMA_signal_7811), .B1_t (new_AGEMA_signal_7812), .B1_f (new_AGEMA_signal_7813), .Z0_t (SubBytesIns_Inst_Sbox_8_M8), .Z0_f (new_AGEMA_signal_8435), .Z1_t (new_AGEMA_signal_8436), .Z1_f (new_AGEMA_signal_8437) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T20), .A0_f (new_AGEMA_signal_7796), .A1_t (new_AGEMA_signal_7797), .A1_f (new_AGEMA_signal_7798), .B0_t (SubBytesIns_Inst_Sbox_8_T17), .B0_f (new_AGEMA_signal_7793), .B1_t (new_AGEMA_signal_7794), .B1_f (new_AGEMA_signal_7795), .Z0_t (SubBytesIns_Inst_Sbox_8_M9), .Z0_f (new_AGEMA_signal_8438), .Z1_t (new_AGEMA_signal_8439), .Z1_f (new_AGEMA_signal_8440) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M9), .A0_f (new_AGEMA_signal_8438), .A1_t (new_AGEMA_signal_8439), .A1_f (new_AGEMA_signal_8440), .B0_t (SubBytesIns_Inst_Sbox_8_M6), .B0_f (new_AGEMA_signal_7811), .B1_t (new_AGEMA_signal_7812), .B1_f (new_AGEMA_signal_7813), .Z0_t (SubBytesIns_Inst_Sbox_8_M10), .Z0_f (new_AGEMA_signal_8816), .Z1_t (new_AGEMA_signal_8817), .Z1_f (new_AGEMA_signal_8818) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T1), .A0_f (new_AGEMA_signal_6586), .A1_t (new_AGEMA_signal_6587), .A1_f (new_AGEMA_signal_6588), .B0_t (SubBytesIns_Inst_Sbox_8_T15), .B0_f (new_AGEMA_signal_7129), .B1_t (new_AGEMA_signal_7130), .B1_f (new_AGEMA_signal_7131), .Z0_t (SubBytesIns_Inst_Sbox_8_M11), .Z0_f (new_AGEMA_signal_7817), .Z1_t (new_AGEMA_signal_7818), .Z1_f (new_AGEMA_signal_7819) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T4), .A0_f (new_AGEMA_signal_6595), .A1_t (new_AGEMA_signal_6596), .A1_f (new_AGEMA_signal_6597), .B0_t (SubBytesIns_Inst_Sbox_8_T27), .B0_f (new_AGEMA_signal_7141), .B1_t (new_AGEMA_signal_7142), .B1_f (new_AGEMA_signal_7143), .Z0_t (SubBytesIns_Inst_Sbox_8_M12), .Z0_f (new_AGEMA_signal_7820), .Z1_t (new_AGEMA_signal_7821), .Z1_f (new_AGEMA_signal_7822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M12), .A0_f (new_AGEMA_signal_7820), .A1_t (new_AGEMA_signal_7821), .A1_f (new_AGEMA_signal_7822), .B0_t (SubBytesIns_Inst_Sbox_8_M11), .B0_f (new_AGEMA_signal_7817), .B1_t (new_AGEMA_signal_7818), .B1_f (new_AGEMA_signal_7819), .Z0_t (SubBytesIns_Inst_Sbox_8_M13), .Z0_f (new_AGEMA_signal_8441), .Z1_t (new_AGEMA_signal_8442), .Z1_f (new_AGEMA_signal_8443) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T2), .A0_f (new_AGEMA_signal_6589), .A1_t (new_AGEMA_signal_6590), .A1_f (new_AGEMA_signal_6591), .B0_t (SubBytesIns_Inst_Sbox_8_T10), .B0_f (new_AGEMA_signal_7787), .B1_t (new_AGEMA_signal_7788), .B1_f (new_AGEMA_signal_7789), .Z0_t (SubBytesIns_Inst_Sbox_8_M14), .Z0_f (new_AGEMA_signal_8444), .Z1_t (new_AGEMA_signal_8445), .Z1_f (new_AGEMA_signal_8446) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M14), .A0_f (new_AGEMA_signal_8444), .A1_t (new_AGEMA_signal_8445), .A1_f (new_AGEMA_signal_8446), .B0_t (SubBytesIns_Inst_Sbox_8_M11), .B0_f (new_AGEMA_signal_7817), .B1_t (new_AGEMA_signal_7818), .B1_f (new_AGEMA_signal_7819), .Z0_t (SubBytesIns_Inst_Sbox_8_M15), .Z0_f (new_AGEMA_signal_8819), .Z1_t (new_AGEMA_signal_8820), .Z1_f (new_AGEMA_signal_8821) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M3), .A0_f (new_AGEMA_signal_8429), .A1_t (new_AGEMA_signal_8430), .A1_f (new_AGEMA_signal_8431), .B0_t (SubBytesIns_Inst_Sbox_8_M2), .B0_f (new_AGEMA_signal_8426), .B1_t (new_AGEMA_signal_8427), .B1_f (new_AGEMA_signal_8428), .Z0_t (SubBytesIns_Inst_Sbox_8_M16), .Z0_f (new_AGEMA_signal_8822), .Z1_t (new_AGEMA_signal_8823), .Z1_f (new_AGEMA_signal_8824) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M5), .A0_f (new_AGEMA_signal_8432), .A1_t (new_AGEMA_signal_8433), .A1_f (new_AGEMA_signal_8434), .B0_t (SubBytesIns_Inst_Sbox_8_T24), .B0_f (new_AGEMA_signal_8420), .B1_t (new_AGEMA_signal_8421), .B1_f (new_AGEMA_signal_8422), .Z0_t (SubBytesIns_Inst_Sbox_8_M17), .Z0_f (new_AGEMA_signal_8825), .Z1_t (new_AGEMA_signal_8826), .Z1_f (new_AGEMA_signal_8827) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M8), .A0_f (new_AGEMA_signal_8435), .A1_t (new_AGEMA_signal_8436), .A1_f (new_AGEMA_signal_8437), .B0_t (SubBytesIns_Inst_Sbox_8_M7), .B0_f (new_AGEMA_signal_7814), .B1_t (new_AGEMA_signal_7815), .B1_f (new_AGEMA_signal_7816), .Z0_t (SubBytesIns_Inst_Sbox_8_M18), .Z0_f (new_AGEMA_signal_8828), .Z1_t (new_AGEMA_signal_8829), .Z1_f (new_AGEMA_signal_8830) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M10), .A0_f (new_AGEMA_signal_8816), .A1_t (new_AGEMA_signal_8817), .A1_f (new_AGEMA_signal_8818), .B0_t (SubBytesIns_Inst_Sbox_8_M15), .B0_f (new_AGEMA_signal_8819), .B1_t (new_AGEMA_signal_8820), .B1_f (new_AGEMA_signal_8821), .Z0_t (SubBytesIns_Inst_Sbox_8_M19), .Z0_f (new_AGEMA_signal_9080), .Z1_t (new_AGEMA_signal_9081), .Z1_f (new_AGEMA_signal_9082) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M16), .A0_f (new_AGEMA_signal_8822), .A1_t (new_AGEMA_signal_8823), .A1_f (new_AGEMA_signal_8824), .B0_t (SubBytesIns_Inst_Sbox_8_M13), .B0_f (new_AGEMA_signal_8441), .B1_t (new_AGEMA_signal_8442), .B1_f (new_AGEMA_signal_8443), .Z0_t (SubBytesIns_Inst_Sbox_8_M20), .Z0_f (new_AGEMA_signal_9083), .Z1_t (new_AGEMA_signal_9084), .Z1_f (new_AGEMA_signal_9085) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M17), .A0_f (new_AGEMA_signal_8825), .A1_t (new_AGEMA_signal_8826), .A1_f (new_AGEMA_signal_8827), .B0_t (SubBytesIns_Inst_Sbox_8_M15), .B0_f (new_AGEMA_signal_8819), .B1_t (new_AGEMA_signal_8820), .B1_f (new_AGEMA_signal_8821), .Z0_t (SubBytesIns_Inst_Sbox_8_M21), .Z0_f (new_AGEMA_signal_9086), .Z1_t (new_AGEMA_signal_9087), .Z1_f (new_AGEMA_signal_9088) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M18), .A0_f (new_AGEMA_signal_8828), .A1_t (new_AGEMA_signal_8829), .A1_f (new_AGEMA_signal_8830), .B0_t (SubBytesIns_Inst_Sbox_8_M13), .B0_f (new_AGEMA_signal_8441), .B1_t (new_AGEMA_signal_8442), .B1_f (new_AGEMA_signal_8443), .Z0_t (SubBytesIns_Inst_Sbox_8_M22), .Z0_f (new_AGEMA_signal_9089), .Z1_t (new_AGEMA_signal_9090), .Z1_f (new_AGEMA_signal_9091) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M19), .A0_f (new_AGEMA_signal_9080), .A1_t (new_AGEMA_signal_9081), .A1_f (new_AGEMA_signal_9082), .B0_t (SubBytesIns_Inst_Sbox_8_T25), .B0_f (new_AGEMA_signal_8423), .B1_t (new_AGEMA_signal_8424), .B1_f (new_AGEMA_signal_8425), .Z0_t (SubBytesIns_Inst_Sbox_8_M23), .Z0_f (new_AGEMA_signal_9320), .Z1_t (new_AGEMA_signal_9321), .Z1_f (new_AGEMA_signal_9322) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M22), .A0_f (new_AGEMA_signal_9089), .A1_t (new_AGEMA_signal_9090), .A1_f (new_AGEMA_signal_9091), .B0_t (SubBytesIns_Inst_Sbox_8_M23), .B0_f (new_AGEMA_signal_9320), .B1_t (new_AGEMA_signal_9321), .B1_f (new_AGEMA_signal_9322), .Z0_t (SubBytesIns_Inst_Sbox_8_M24), .Z0_f (new_AGEMA_signal_9596), .Z1_t (new_AGEMA_signal_9597), .Z1_f (new_AGEMA_signal_9598) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M22), .A0_f (new_AGEMA_signal_9089), .A1_t (new_AGEMA_signal_9090), .A1_f (new_AGEMA_signal_9091), .B0_t (SubBytesIns_Inst_Sbox_8_M20), .B0_f (new_AGEMA_signal_9083), .B1_t (new_AGEMA_signal_9084), .B1_f (new_AGEMA_signal_9085), .Z0_t (SubBytesIns_Inst_Sbox_8_M25), .Z0_f (new_AGEMA_signal_9323), .Z1_t (new_AGEMA_signal_9324), .Z1_f (new_AGEMA_signal_9325) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M21), .A0_f (new_AGEMA_signal_9086), .A1_t (new_AGEMA_signal_9087), .A1_f (new_AGEMA_signal_9088), .B0_t (SubBytesIns_Inst_Sbox_8_M25), .B0_f (new_AGEMA_signal_9323), .B1_t (new_AGEMA_signal_9324), .B1_f (new_AGEMA_signal_9325), .Z0_t (SubBytesIns_Inst_Sbox_8_M26), .Z0_f (new_AGEMA_signal_9599), .Z1_t (new_AGEMA_signal_9600), .Z1_f (new_AGEMA_signal_9601) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M20), .A0_f (new_AGEMA_signal_9083), .A1_t (new_AGEMA_signal_9084), .A1_f (new_AGEMA_signal_9085), .B0_t (SubBytesIns_Inst_Sbox_8_M21), .B0_f (new_AGEMA_signal_9086), .B1_t (new_AGEMA_signal_9087), .B1_f (new_AGEMA_signal_9088), .Z0_t (SubBytesIns_Inst_Sbox_8_M27), .Z0_f (new_AGEMA_signal_9326), .Z1_t (new_AGEMA_signal_9327), .Z1_f (new_AGEMA_signal_9328) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M23), .A0_f (new_AGEMA_signal_9320), .A1_t (new_AGEMA_signal_9321), .A1_f (new_AGEMA_signal_9322), .B0_t (SubBytesIns_Inst_Sbox_8_M25), .B0_f (new_AGEMA_signal_9323), .B1_t (new_AGEMA_signal_9324), .B1_f (new_AGEMA_signal_9325), .Z0_t (SubBytesIns_Inst_Sbox_8_M28), .Z0_f (new_AGEMA_signal_9602), .Z1_t (new_AGEMA_signal_9603), .Z1_f (new_AGEMA_signal_9604) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M28), .A0_f (new_AGEMA_signal_9602), .A1_t (new_AGEMA_signal_9603), .A1_f (new_AGEMA_signal_9604), .B0_t (SubBytesIns_Inst_Sbox_8_M27), .B0_f (new_AGEMA_signal_9326), .B1_t (new_AGEMA_signal_9327), .B1_f (new_AGEMA_signal_9328), .Z0_t (SubBytesIns_Inst_Sbox_8_M29), .Z0_f (new_AGEMA_signal_9896), .Z1_t (new_AGEMA_signal_9897), .Z1_f (new_AGEMA_signal_9898) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M26), .A0_f (new_AGEMA_signal_9599), .A1_t (new_AGEMA_signal_9600), .A1_f (new_AGEMA_signal_9601), .B0_t (SubBytesIns_Inst_Sbox_8_M24), .B0_f (new_AGEMA_signal_9596), .B1_t (new_AGEMA_signal_9597), .B1_f (new_AGEMA_signal_9598), .Z0_t (SubBytesIns_Inst_Sbox_8_M30), .Z0_f (new_AGEMA_signal_9899), .Z1_t (new_AGEMA_signal_9900), .Z1_f (new_AGEMA_signal_9901) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M20), .A0_f (new_AGEMA_signal_9083), .A1_t (new_AGEMA_signal_9084), .A1_f (new_AGEMA_signal_9085), .B0_t (SubBytesIns_Inst_Sbox_8_M23), .B0_f (new_AGEMA_signal_9320), .B1_t (new_AGEMA_signal_9321), .B1_f (new_AGEMA_signal_9322), .Z0_t (SubBytesIns_Inst_Sbox_8_M31), .Z0_f (new_AGEMA_signal_9605), .Z1_t (new_AGEMA_signal_9606), .Z1_f (new_AGEMA_signal_9607) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M27), .A0_f (new_AGEMA_signal_9326), .A1_t (new_AGEMA_signal_9327), .A1_f (new_AGEMA_signal_9328), .B0_t (SubBytesIns_Inst_Sbox_8_M31), .B0_f (new_AGEMA_signal_9605), .B1_t (new_AGEMA_signal_9606), .B1_f (new_AGEMA_signal_9607), .Z0_t (SubBytesIns_Inst_Sbox_8_M32), .Z0_f (new_AGEMA_signal_9902), .Z1_t (new_AGEMA_signal_9903), .Z1_f (new_AGEMA_signal_9904) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M27), .A0_f (new_AGEMA_signal_9326), .A1_t (new_AGEMA_signal_9327), .A1_f (new_AGEMA_signal_9328), .B0_t (SubBytesIns_Inst_Sbox_8_M25), .B0_f (new_AGEMA_signal_9323), .B1_t (new_AGEMA_signal_9324), .B1_f (new_AGEMA_signal_9325), .Z0_t (SubBytesIns_Inst_Sbox_8_M33), .Z0_f (new_AGEMA_signal_9608), .Z1_t (new_AGEMA_signal_9609), .Z1_f (new_AGEMA_signal_9610) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M21), .A0_f (new_AGEMA_signal_9086), .A1_t (new_AGEMA_signal_9087), .A1_f (new_AGEMA_signal_9088), .B0_t (SubBytesIns_Inst_Sbox_8_M22), .B0_f (new_AGEMA_signal_9089), .B1_t (new_AGEMA_signal_9090), .B1_f (new_AGEMA_signal_9091), .Z0_t (SubBytesIns_Inst_Sbox_8_M34), .Z0_f (new_AGEMA_signal_9329), .Z1_t (new_AGEMA_signal_9330), .Z1_f (new_AGEMA_signal_9331) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M24), .A0_f (new_AGEMA_signal_9596), .A1_t (new_AGEMA_signal_9597), .A1_f (new_AGEMA_signal_9598), .B0_t (SubBytesIns_Inst_Sbox_8_M34), .B0_f (new_AGEMA_signal_9329), .B1_t (new_AGEMA_signal_9330), .B1_f (new_AGEMA_signal_9331), .Z0_t (SubBytesIns_Inst_Sbox_8_M35), .Z0_f (new_AGEMA_signal_9905), .Z1_t (new_AGEMA_signal_9906), .Z1_f (new_AGEMA_signal_9907) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M24), .A0_f (new_AGEMA_signal_9596), .A1_t (new_AGEMA_signal_9597), .A1_f (new_AGEMA_signal_9598), .B0_t (SubBytesIns_Inst_Sbox_8_M25), .B0_f (new_AGEMA_signal_9323), .B1_t (new_AGEMA_signal_9324), .B1_f (new_AGEMA_signal_9325), .Z0_t (SubBytesIns_Inst_Sbox_8_M36), .Z0_f (new_AGEMA_signal_9908), .Z1_t (new_AGEMA_signal_9909), .Z1_f (new_AGEMA_signal_9910) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M21), .A0_f (new_AGEMA_signal_9086), .A1_t (new_AGEMA_signal_9087), .A1_f (new_AGEMA_signal_9088), .B0_t (SubBytesIns_Inst_Sbox_8_M29), .B0_f (new_AGEMA_signal_9896), .B1_t (new_AGEMA_signal_9897), .B1_f (new_AGEMA_signal_9898), .Z0_t (SubBytesIns_Inst_Sbox_8_M37), .Z0_f (new_AGEMA_signal_10160), .Z1_t (new_AGEMA_signal_10161), .Z1_f (new_AGEMA_signal_10162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M32), .A0_f (new_AGEMA_signal_9902), .A1_t (new_AGEMA_signal_9903), .A1_f (new_AGEMA_signal_9904), .B0_t (SubBytesIns_Inst_Sbox_8_M33), .B0_f (new_AGEMA_signal_9608), .B1_t (new_AGEMA_signal_9609), .B1_f (new_AGEMA_signal_9610), .Z0_t (SubBytesIns_Inst_Sbox_8_M38), .Z0_f (new_AGEMA_signal_10163), .Z1_t (new_AGEMA_signal_10164), .Z1_f (new_AGEMA_signal_10165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M23), .A0_f (new_AGEMA_signal_9320), .A1_t (new_AGEMA_signal_9321), .A1_f (new_AGEMA_signal_9322), .B0_t (SubBytesIns_Inst_Sbox_8_M30), .B0_f (new_AGEMA_signal_9899), .B1_t (new_AGEMA_signal_9900), .B1_f (new_AGEMA_signal_9901), .Z0_t (SubBytesIns_Inst_Sbox_8_M39), .Z0_f (new_AGEMA_signal_10166), .Z1_t (new_AGEMA_signal_10167), .Z1_f (new_AGEMA_signal_10168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M35), .A0_f (new_AGEMA_signal_9905), .A1_t (new_AGEMA_signal_9906), .A1_f (new_AGEMA_signal_9907), .B0_t (SubBytesIns_Inst_Sbox_8_M36), .B0_f (new_AGEMA_signal_9908), .B1_t (new_AGEMA_signal_9909), .B1_f (new_AGEMA_signal_9910), .Z0_t (SubBytesIns_Inst_Sbox_8_M40), .Z0_f (new_AGEMA_signal_10169), .Z1_t (new_AGEMA_signal_10170), .Z1_f (new_AGEMA_signal_10171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M38), .A0_f (new_AGEMA_signal_10163), .A1_t (new_AGEMA_signal_10164), .A1_f (new_AGEMA_signal_10165), .B0_t (SubBytesIns_Inst_Sbox_8_M40), .B0_f (new_AGEMA_signal_10169), .B1_t (new_AGEMA_signal_10170), .B1_f (new_AGEMA_signal_10171), .Z0_t (SubBytesIns_Inst_Sbox_8_M41), .Z0_f (new_AGEMA_signal_10688), .Z1_t (new_AGEMA_signal_10689), .Z1_f (new_AGEMA_signal_10690) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M37), .A0_f (new_AGEMA_signal_10160), .A1_t (new_AGEMA_signal_10161), .A1_f (new_AGEMA_signal_10162), .B0_t (SubBytesIns_Inst_Sbox_8_M39), .B0_f (new_AGEMA_signal_10166), .B1_t (new_AGEMA_signal_10167), .B1_f (new_AGEMA_signal_10168), .Z0_t (SubBytesIns_Inst_Sbox_8_M42), .Z0_f (new_AGEMA_signal_10691), .Z1_t (new_AGEMA_signal_10692), .Z1_f (new_AGEMA_signal_10693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M37), .A0_f (new_AGEMA_signal_10160), .A1_t (new_AGEMA_signal_10161), .A1_f (new_AGEMA_signal_10162), .B0_t (SubBytesIns_Inst_Sbox_8_M38), .B0_f (new_AGEMA_signal_10163), .B1_t (new_AGEMA_signal_10164), .B1_f (new_AGEMA_signal_10165), .Z0_t (SubBytesIns_Inst_Sbox_8_M43), .Z0_f (new_AGEMA_signal_10694), .Z1_t (new_AGEMA_signal_10695), .Z1_f (new_AGEMA_signal_10696) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M39), .A0_f (new_AGEMA_signal_10166), .A1_t (new_AGEMA_signal_10167), .A1_f (new_AGEMA_signal_10168), .B0_t (SubBytesIns_Inst_Sbox_8_M40), .B0_f (new_AGEMA_signal_10169), .B1_t (new_AGEMA_signal_10170), .B1_f (new_AGEMA_signal_10171), .Z0_t (SubBytesIns_Inst_Sbox_8_M44), .Z0_f (new_AGEMA_signal_10697), .Z1_t (new_AGEMA_signal_10698), .Z1_f (new_AGEMA_signal_10699) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M42), .A0_f (new_AGEMA_signal_10691), .A1_t (new_AGEMA_signal_10692), .A1_f (new_AGEMA_signal_10693), .B0_t (SubBytesIns_Inst_Sbox_8_M41), .B0_f (new_AGEMA_signal_10688), .B1_t (new_AGEMA_signal_10689), .B1_f (new_AGEMA_signal_10690), .Z0_t (SubBytesIns_Inst_Sbox_8_M45), .Z0_f (new_AGEMA_signal_11408), .Z1_t (new_AGEMA_signal_11409), .Z1_f (new_AGEMA_signal_11410) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M44), .A0_f (new_AGEMA_signal_10697), .A1_t (new_AGEMA_signal_10698), .A1_f (new_AGEMA_signal_10699), .B0_t (SubBytesIns_Inst_Sbox_8_T6), .B0_f (new_AGEMA_signal_7120), .B1_t (new_AGEMA_signal_7121), .B1_f (new_AGEMA_signal_7122), .Z0_t (SubBytesIns_Inst_Sbox_8_M46), .Z0_f (new_AGEMA_signal_11411), .Z1_t (new_AGEMA_signal_11412), .Z1_f (new_AGEMA_signal_11413) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M40), .A0_f (new_AGEMA_signal_10169), .A1_t (new_AGEMA_signal_10170), .A1_f (new_AGEMA_signal_10171), .B0_t (SubBytesIns_Inst_Sbox_8_T8), .B0_f (new_AGEMA_signal_7784), .B1_t (new_AGEMA_signal_7785), .B1_f (new_AGEMA_signal_7786), .Z0_t (SubBytesIns_Inst_Sbox_8_M47), .Z0_f (new_AGEMA_signal_10700), .Z1_t (new_AGEMA_signal_10701), .Z1_f (new_AGEMA_signal_10702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M39), .A0_f (new_AGEMA_signal_10166), .A1_t (new_AGEMA_signal_10167), .A1_f (new_AGEMA_signal_10168), .B0_t (ciphertext_s0_t[64]), .B0_f (ciphertext_s0_f[64]), .B1_t (ciphertext_s1_t[64]), .B1_f (ciphertext_s1_f[64]), .Z0_t (SubBytesIns_Inst_Sbox_8_M48), .Z0_f (new_AGEMA_signal_10703), .Z1_t (new_AGEMA_signal_10704), .Z1_f (new_AGEMA_signal_10705) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M43), .A0_f (new_AGEMA_signal_10694), .A1_t (new_AGEMA_signal_10695), .A1_f (new_AGEMA_signal_10696), .B0_t (SubBytesIns_Inst_Sbox_8_T16), .B0_f (new_AGEMA_signal_7132), .B1_t (new_AGEMA_signal_7133), .B1_f (new_AGEMA_signal_7134), .Z0_t (SubBytesIns_Inst_Sbox_8_M49), .Z0_f (new_AGEMA_signal_11414), .Z1_t (new_AGEMA_signal_11415), .Z1_f (new_AGEMA_signal_11416) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M38), .A0_f (new_AGEMA_signal_10163), .A1_t (new_AGEMA_signal_10164), .A1_f (new_AGEMA_signal_10165), .B0_t (SubBytesIns_Inst_Sbox_8_T9), .B0_f (new_AGEMA_signal_7123), .B1_t (new_AGEMA_signal_7124), .B1_f (new_AGEMA_signal_7125), .Z0_t (SubBytesIns_Inst_Sbox_8_M50), .Z0_f (new_AGEMA_signal_10706), .Z1_t (new_AGEMA_signal_10707), .Z1_f (new_AGEMA_signal_10708) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M37), .A0_f (new_AGEMA_signal_10160), .A1_t (new_AGEMA_signal_10161), .A1_f (new_AGEMA_signal_10162), .B0_t (SubBytesIns_Inst_Sbox_8_T17), .B0_f (new_AGEMA_signal_7793), .B1_t (new_AGEMA_signal_7794), .B1_f (new_AGEMA_signal_7795), .Z0_t (SubBytesIns_Inst_Sbox_8_M51), .Z0_f (new_AGEMA_signal_10709), .Z1_t (new_AGEMA_signal_10710), .Z1_f (new_AGEMA_signal_10711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M42), .A0_f (new_AGEMA_signal_10691), .A1_t (new_AGEMA_signal_10692), .A1_f (new_AGEMA_signal_10693), .B0_t (SubBytesIns_Inst_Sbox_8_T15), .B0_f (new_AGEMA_signal_7129), .B1_t (new_AGEMA_signal_7130), .B1_f (new_AGEMA_signal_7131), .Z0_t (SubBytesIns_Inst_Sbox_8_M52), .Z0_f (new_AGEMA_signal_11417), .Z1_t (new_AGEMA_signal_11418), .Z1_f (new_AGEMA_signal_11419) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M45), .A0_f (new_AGEMA_signal_11408), .A1_t (new_AGEMA_signal_11409), .A1_f (new_AGEMA_signal_11410), .B0_t (SubBytesIns_Inst_Sbox_8_T27), .B0_f (new_AGEMA_signal_7141), .B1_t (new_AGEMA_signal_7142), .B1_f (new_AGEMA_signal_7143), .Z0_t (SubBytesIns_Inst_Sbox_8_M53), .Z0_f (new_AGEMA_signal_12056), .Z1_t (new_AGEMA_signal_12057), .Z1_f (new_AGEMA_signal_12058) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M41), .A0_f (new_AGEMA_signal_10688), .A1_t (new_AGEMA_signal_10689), .A1_f (new_AGEMA_signal_10690), .B0_t (SubBytesIns_Inst_Sbox_8_T10), .B0_f (new_AGEMA_signal_7787), .B1_t (new_AGEMA_signal_7788), .B1_f (new_AGEMA_signal_7789), .Z0_t (SubBytesIns_Inst_Sbox_8_M54), .Z0_f (new_AGEMA_signal_11420), .Z1_t (new_AGEMA_signal_11421), .Z1_f (new_AGEMA_signal_11422) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M44), .A0_f (new_AGEMA_signal_10697), .A1_t (new_AGEMA_signal_10698), .A1_f (new_AGEMA_signal_10699), .B0_t (SubBytesIns_Inst_Sbox_8_T13), .B0_f (new_AGEMA_signal_7126), .B1_t (new_AGEMA_signal_7127), .B1_f (new_AGEMA_signal_7128), .Z0_t (SubBytesIns_Inst_Sbox_8_M55), .Z0_f (new_AGEMA_signal_11423), .Z1_t (new_AGEMA_signal_11424), .Z1_f (new_AGEMA_signal_11425) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M40), .A0_f (new_AGEMA_signal_10169), .A1_t (new_AGEMA_signal_10170), .A1_f (new_AGEMA_signal_10171), .B0_t (SubBytesIns_Inst_Sbox_8_T23), .B0_f (new_AGEMA_signal_7799), .B1_t (new_AGEMA_signal_7800), .B1_f (new_AGEMA_signal_7801), .Z0_t (SubBytesIns_Inst_Sbox_8_M56), .Z0_f (new_AGEMA_signal_10712), .Z1_t (new_AGEMA_signal_10713), .Z1_f (new_AGEMA_signal_10714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M39), .A0_f (new_AGEMA_signal_10166), .A1_t (new_AGEMA_signal_10167), .A1_f (new_AGEMA_signal_10168), .B0_t (SubBytesIns_Inst_Sbox_8_T19), .B0_f (new_AGEMA_signal_7135), .B1_t (new_AGEMA_signal_7136), .B1_f (new_AGEMA_signal_7137), .Z0_t (SubBytesIns_Inst_Sbox_8_M57), .Z0_f (new_AGEMA_signal_10715), .Z1_t (new_AGEMA_signal_10716), .Z1_f (new_AGEMA_signal_10717) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M43), .A0_f (new_AGEMA_signal_10694), .A1_t (new_AGEMA_signal_10695), .A1_f (new_AGEMA_signal_10696), .B0_t (SubBytesIns_Inst_Sbox_8_T3), .B0_f (new_AGEMA_signal_6592), .B1_t (new_AGEMA_signal_6593), .B1_f (new_AGEMA_signal_6594), .Z0_t (SubBytesIns_Inst_Sbox_8_M58), .Z0_f (new_AGEMA_signal_11426), .Z1_t (new_AGEMA_signal_11427), .Z1_f (new_AGEMA_signal_11428) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M38), .A0_f (new_AGEMA_signal_10163), .A1_t (new_AGEMA_signal_10164), .A1_f (new_AGEMA_signal_10165), .B0_t (SubBytesIns_Inst_Sbox_8_T22), .B0_f (new_AGEMA_signal_7138), .B1_t (new_AGEMA_signal_7139), .B1_f (new_AGEMA_signal_7140), .Z0_t (SubBytesIns_Inst_Sbox_8_M59), .Z0_f (new_AGEMA_signal_10718), .Z1_t (new_AGEMA_signal_10719), .Z1_f (new_AGEMA_signal_10720) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M37), .A0_f (new_AGEMA_signal_10160), .A1_t (new_AGEMA_signal_10161), .A1_f (new_AGEMA_signal_10162), .B0_t (SubBytesIns_Inst_Sbox_8_T20), .B0_f (new_AGEMA_signal_7796), .B1_t (new_AGEMA_signal_7797), .B1_f (new_AGEMA_signal_7798), .Z0_t (SubBytesIns_Inst_Sbox_8_M60), .Z0_f (new_AGEMA_signal_10721), .Z1_t (new_AGEMA_signal_10722), .Z1_f (new_AGEMA_signal_10723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M42), .A0_f (new_AGEMA_signal_10691), .A1_t (new_AGEMA_signal_10692), .A1_f (new_AGEMA_signal_10693), .B0_t (SubBytesIns_Inst_Sbox_8_T1), .B0_f (new_AGEMA_signal_6586), .B1_t (new_AGEMA_signal_6587), .B1_f (new_AGEMA_signal_6588), .Z0_t (SubBytesIns_Inst_Sbox_8_M61), .Z0_f (new_AGEMA_signal_11429), .Z1_t (new_AGEMA_signal_11430), .Z1_f (new_AGEMA_signal_11431) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M45), .A0_f (new_AGEMA_signal_11408), .A1_t (new_AGEMA_signal_11409), .A1_f (new_AGEMA_signal_11410), .B0_t (SubBytesIns_Inst_Sbox_8_T4), .B0_f (new_AGEMA_signal_6595), .B1_t (new_AGEMA_signal_6596), .B1_f (new_AGEMA_signal_6597), .Z0_t (SubBytesIns_Inst_Sbox_8_M62), .Z0_f (new_AGEMA_signal_12059), .Z1_t (new_AGEMA_signal_12060), .Z1_f (new_AGEMA_signal_12061) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M41), .A0_f (new_AGEMA_signal_10688), .A1_t (new_AGEMA_signal_10689), .A1_f (new_AGEMA_signal_10690), .B0_t (SubBytesIns_Inst_Sbox_8_T2), .B0_f (new_AGEMA_signal_6589), .B1_t (new_AGEMA_signal_6590), .B1_f (new_AGEMA_signal_6591), .Z0_t (SubBytesIns_Inst_Sbox_8_M63), .Z0_f (new_AGEMA_signal_11432), .Z1_t (new_AGEMA_signal_11433), .Z1_f (new_AGEMA_signal_11434) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M61), .A0_f (new_AGEMA_signal_11429), .A1_t (new_AGEMA_signal_11430), .A1_f (new_AGEMA_signal_11431), .B0_t (SubBytesIns_Inst_Sbox_8_M62), .B0_f (new_AGEMA_signal_12059), .B1_t (new_AGEMA_signal_12060), .B1_f (new_AGEMA_signal_12061), .Z0_t (SubBytesIns_Inst_Sbox_8_L0), .Z0_f (new_AGEMA_signal_12620), .Z1_t (new_AGEMA_signal_12621), .Z1_f (new_AGEMA_signal_12622) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M50), .A0_f (new_AGEMA_signal_10706), .A1_t (new_AGEMA_signal_10707), .A1_f (new_AGEMA_signal_10708), .B0_t (SubBytesIns_Inst_Sbox_8_M56), .B0_f (new_AGEMA_signal_10712), .B1_t (new_AGEMA_signal_10713), .B1_f (new_AGEMA_signal_10714), .Z0_t (SubBytesIns_Inst_Sbox_8_L1), .Z0_f (new_AGEMA_signal_11435), .Z1_t (new_AGEMA_signal_11436), .Z1_f (new_AGEMA_signal_11437) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M46), .A0_f (new_AGEMA_signal_11411), .A1_t (new_AGEMA_signal_11412), .A1_f (new_AGEMA_signal_11413), .B0_t (SubBytesIns_Inst_Sbox_8_M48), .B0_f (new_AGEMA_signal_10703), .B1_t (new_AGEMA_signal_10704), .B1_f (new_AGEMA_signal_10705), .Z0_t (SubBytesIns_Inst_Sbox_8_L2), .Z0_f (new_AGEMA_signal_12062), .Z1_t (new_AGEMA_signal_12063), .Z1_f (new_AGEMA_signal_12064) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M47), .A0_f (new_AGEMA_signal_10700), .A1_t (new_AGEMA_signal_10701), .A1_f (new_AGEMA_signal_10702), .B0_t (SubBytesIns_Inst_Sbox_8_M55), .B0_f (new_AGEMA_signal_11423), .B1_t (new_AGEMA_signal_11424), .B1_f (new_AGEMA_signal_11425), .Z0_t (SubBytesIns_Inst_Sbox_8_L3), .Z0_f (new_AGEMA_signal_12065), .Z1_t (new_AGEMA_signal_12066), .Z1_f (new_AGEMA_signal_12067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M54), .A0_f (new_AGEMA_signal_11420), .A1_t (new_AGEMA_signal_11421), .A1_f (new_AGEMA_signal_11422), .B0_t (SubBytesIns_Inst_Sbox_8_M58), .B0_f (new_AGEMA_signal_11426), .B1_t (new_AGEMA_signal_11427), .B1_f (new_AGEMA_signal_11428), .Z0_t (SubBytesIns_Inst_Sbox_8_L4), .Z0_f (new_AGEMA_signal_12068), .Z1_t (new_AGEMA_signal_12069), .Z1_f (new_AGEMA_signal_12070) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M49), .A0_f (new_AGEMA_signal_11414), .A1_t (new_AGEMA_signal_11415), .A1_f (new_AGEMA_signal_11416), .B0_t (SubBytesIns_Inst_Sbox_8_M61), .B0_f (new_AGEMA_signal_11429), .B1_t (new_AGEMA_signal_11430), .B1_f (new_AGEMA_signal_11431), .Z0_t (SubBytesIns_Inst_Sbox_8_L5), .Z0_f (new_AGEMA_signal_12071), .Z1_t (new_AGEMA_signal_12072), .Z1_f (new_AGEMA_signal_12073) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M62), .A0_f (new_AGEMA_signal_12059), .A1_t (new_AGEMA_signal_12060), .A1_f (new_AGEMA_signal_12061), .B0_t (SubBytesIns_Inst_Sbox_8_L5), .B0_f (new_AGEMA_signal_12071), .B1_t (new_AGEMA_signal_12072), .B1_f (new_AGEMA_signal_12073), .Z0_t (SubBytesIns_Inst_Sbox_8_L6), .Z0_f (new_AGEMA_signal_12623), .Z1_t (new_AGEMA_signal_12624), .Z1_f (new_AGEMA_signal_12625) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M46), .A0_f (new_AGEMA_signal_11411), .A1_t (new_AGEMA_signal_11412), .A1_f (new_AGEMA_signal_11413), .B0_t (SubBytesIns_Inst_Sbox_8_L3), .B0_f (new_AGEMA_signal_12065), .B1_t (new_AGEMA_signal_12066), .B1_f (new_AGEMA_signal_12067), .Z0_t (SubBytesIns_Inst_Sbox_8_L7), .Z0_f (new_AGEMA_signal_12626), .Z1_t (new_AGEMA_signal_12627), .Z1_f (new_AGEMA_signal_12628) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M51), .A0_f (new_AGEMA_signal_10709), .A1_t (new_AGEMA_signal_10710), .A1_f (new_AGEMA_signal_10711), .B0_t (SubBytesIns_Inst_Sbox_8_M59), .B0_f (new_AGEMA_signal_10718), .B1_t (new_AGEMA_signal_10719), .B1_f (new_AGEMA_signal_10720), .Z0_t (SubBytesIns_Inst_Sbox_8_L8), .Z0_f (new_AGEMA_signal_11438), .Z1_t (new_AGEMA_signal_11439), .Z1_f (new_AGEMA_signal_11440) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M52), .A0_f (new_AGEMA_signal_11417), .A1_t (new_AGEMA_signal_11418), .A1_f (new_AGEMA_signal_11419), .B0_t (SubBytesIns_Inst_Sbox_8_M53), .B0_f (new_AGEMA_signal_12056), .B1_t (new_AGEMA_signal_12057), .B1_f (new_AGEMA_signal_12058), .Z0_t (SubBytesIns_Inst_Sbox_8_L9), .Z0_f (new_AGEMA_signal_12629), .Z1_t (new_AGEMA_signal_12630), .Z1_f (new_AGEMA_signal_12631) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M53), .A0_f (new_AGEMA_signal_12056), .A1_t (new_AGEMA_signal_12057), .A1_f (new_AGEMA_signal_12058), .B0_t (SubBytesIns_Inst_Sbox_8_L4), .B0_f (new_AGEMA_signal_12068), .B1_t (new_AGEMA_signal_12069), .B1_f (new_AGEMA_signal_12070), .Z0_t (SubBytesIns_Inst_Sbox_8_L10), .Z0_f (new_AGEMA_signal_12632), .Z1_t (new_AGEMA_signal_12633), .Z1_f (new_AGEMA_signal_12634) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M60), .A0_f (new_AGEMA_signal_10721), .A1_t (new_AGEMA_signal_10722), .A1_f (new_AGEMA_signal_10723), .B0_t (SubBytesIns_Inst_Sbox_8_L2), .B0_f (new_AGEMA_signal_12062), .B1_t (new_AGEMA_signal_12063), .B1_f (new_AGEMA_signal_12064), .Z0_t (SubBytesIns_Inst_Sbox_8_L11), .Z0_f (new_AGEMA_signal_12635), .Z1_t (new_AGEMA_signal_12636), .Z1_f (new_AGEMA_signal_12637) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M48), .A0_f (new_AGEMA_signal_10703), .A1_t (new_AGEMA_signal_10704), .A1_f (new_AGEMA_signal_10705), .B0_t (SubBytesIns_Inst_Sbox_8_M51), .B0_f (new_AGEMA_signal_10709), .B1_t (new_AGEMA_signal_10710), .B1_f (new_AGEMA_signal_10711), .Z0_t (SubBytesIns_Inst_Sbox_8_L12), .Z0_f (new_AGEMA_signal_11441), .Z1_t (new_AGEMA_signal_11442), .Z1_f (new_AGEMA_signal_11443) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M50), .A0_f (new_AGEMA_signal_10706), .A1_t (new_AGEMA_signal_10707), .A1_f (new_AGEMA_signal_10708), .B0_t (SubBytesIns_Inst_Sbox_8_L0), .B0_f (new_AGEMA_signal_12620), .B1_t (new_AGEMA_signal_12621), .B1_f (new_AGEMA_signal_12622), .Z0_t (SubBytesIns_Inst_Sbox_8_L13), .Z0_f (new_AGEMA_signal_13232), .Z1_t (new_AGEMA_signal_13233), .Z1_f (new_AGEMA_signal_13234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M52), .A0_f (new_AGEMA_signal_11417), .A1_t (new_AGEMA_signal_11418), .A1_f (new_AGEMA_signal_11419), .B0_t (SubBytesIns_Inst_Sbox_8_M61), .B0_f (new_AGEMA_signal_11429), .B1_t (new_AGEMA_signal_11430), .B1_f (new_AGEMA_signal_11431), .Z0_t (SubBytesIns_Inst_Sbox_8_L14), .Z0_f (new_AGEMA_signal_12074), .Z1_t (new_AGEMA_signal_12075), .Z1_f (new_AGEMA_signal_12076) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M55), .A0_f (new_AGEMA_signal_11423), .A1_t (new_AGEMA_signal_11424), .A1_f (new_AGEMA_signal_11425), .B0_t (SubBytesIns_Inst_Sbox_8_L1), .B0_f (new_AGEMA_signal_11435), .B1_t (new_AGEMA_signal_11436), .B1_f (new_AGEMA_signal_11437), .Z0_t (SubBytesIns_Inst_Sbox_8_L15), .Z0_f (new_AGEMA_signal_12077), .Z1_t (new_AGEMA_signal_12078), .Z1_f (new_AGEMA_signal_12079) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M56), .A0_f (new_AGEMA_signal_10712), .A1_t (new_AGEMA_signal_10713), .A1_f (new_AGEMA_signal_10714), .B0_t (SubBytesIns_Inst_Sbox_8_L0), .B0_f (new_AGEMA_signal_12620), .B1_t (new_AGEMA_signal_12621), .B1_f (new_AGEMA_signal_12622), .Z0_t (SubBytesIns_Inst_Sbox_8_L16), .Z0_f (new_AGEMA_signal_13235), .Z1_t (new_AGEMA_signal_13236), .Z1_f (new_AGEMA_signal_13237) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M57), .A0_f (new_AGEMA_signal_10715), .A1_t (new_AGEMA_signal_10716), .A1_f (new_AGEMA_signal_10717), .B0_t (SubBytesIns_Inst_Sbox_8_L1), .B0_f (new_AGEMA_signal_11435), .B1_t (new_AGEMA_signal_11436), .B1_f (new_AGEMA_signal_11437), .Z0_t (SubBytesIns_Inst_Sbox_8_L17), .Z0_f (new_AGEMA_signal_12080), .Z1_t (new_AGEMA_signal_12081), .Z1_f (new_AGEMA_signal_12082) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M58), .A0_f (new_AGEMA_signal_11426), .A1_t (new_AGEMA_signal_11427), .A1_f (new_AGEMA_signal_11428), .B0_t (SubBytesIns_Inst_Sbox_8_L8), .B0_f (new_AGEMA_signal_11438), .B1_t (new_AGEMA_signal_11439), .B1_f (new_AGEMA_signal_11440), .Z0_t (SubBytesIns_Inst_Sbox_8_L18), .Z0_f (new_AGEMA_signal_12083), .Z1_t (new_AGEMA_signal_12084), .Z1_f (new_AGEMA_signal_12085) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M63), .A0_f (new_AGEMA_signal_11432), .A1_t (new_AGEMA_signal_11433), .A1_f (new_AGEMA_signal_11434), .B0_t (SubBytesIns_Inst_Sbox_8_L4), .B0_f (new_AGEMA_signal_12068), .B1_t (new_AGEMA_signal_12069), .B1_f (new_AGEMA_signal_12070), .Z0_t (SubBytesIns_Inst_Sbox_8_L19), .Z0_f (new_AGEMA_signal_12638), .Z1_t (new_AGEMA_signal_12639), .Z1_f (new_AGEMA_signal_12640) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L0), .A0_f (new_AGEMA_signal_12620), .A1_t (new_AGEMA_signal_12621), .A1_f (new_AGEMA_signal_12622), .B0_t (SubBytesIns_Inst_Sbox_8_L1), .B0_f (new_AGEMA_signal_11435), .B1_t (new_AGEMA_signal_11436), .B1_f (new_AGEMA_signal_11437), .Z0_t (SubBytesIns_Inst_Sbox_8_L20), .Z0_f (new_AGEMA_signal_13238), .Z1_t (new_AGEMA_signal_13239), .Z1_f (new_AGEMA_signal_13240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L1), .A0_f (new_AGEMA_signal_11435), .A1_t (new_AGEMA_signal_11436), .A1_f (new_AGEMA_signal_11437), .B0_t (SubBytesIns_Inst_Sbox_8_L7), .B0_f (new_AGEMA_signal_12626), .B1_t (new_AGEMA_signal_12627), .B1_f (new_AGEMA_signal_12628), .Z0_t (SubBytesIns_Inst_Sbox_8_L21), .Z0_f (new_AGEMA_signal_13241), .Z1_t (new_AGEMA_signal_13242), .Z1_f (new_AGEMA_signal_13243) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L3), .A0_f (new_AGEMA_signal_12065), .A1_t (new_AGEMA_signal_12066), .A1_f (new_AGEMA_signal_12067), .B0_t (SubBytesIns_Inst_Sbox_8_L12), .B0_f (new_AGEMA_signal_11441), .B1_t (new_AGEMA_signal_11442), .B1_f (new_AGEMA_signal_11443), .Z0_t (SubBytesIns_Inst_Sbox_8_L22), .Z0_f (new_AGEMA_signal_12641), .Z1_t (new_AGEMA_signal_12642), .Z1_f (new_AGEMA_signal_12643) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L18), .A0_f (new_AGEMA_signal_12083), .A1_t (new_AGEMA_signal_12084), .A1_f (new_AGEMA_signal_12085), .B0_t (SubBytesIns_Inst_Sbox_8_L2), .B0_f (new_AGEMA_signal_12062), .B1_t (new_AGEMA_signal_12063), .B1_f (new_AGEMA_signal_12064), .Z0_t (SubBytesIns_Inst_Sbox_8_L23), .Z0_f (new_AGEMA_signal_12644), .Z1_t (new_AGEMA_signal_12645), .Z1_f (new_AGEMA_signal_12646) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L15), .A0_f (new_AGEMA_signal_12077), .A1_t (new_AGEMA_signal_12078), .A1_f (new_AGEMA_signal_12079), .B0_t (SubBytesIns_Inst_Sbox_8_L9), .B0_f (new_AGEMA_signal_12629), .B1_t (new_AGEMA_signal_12630), .B1_f (new_AGEMA_signal_12631), .Z0_t (SubBytesIns_Inst_Sbox_8_L24), .Z0_f (new_AGEMA_signal_13244), .Z1_t (new_AGEMA_signal_13245), .Z1_f (new_AGEMA_signal_13246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L6), .A0_f (new_AGEMA_signal_12623), .A1_t (new_AGEMA_signal_12624), .A1_f (new_AGEMA_signal_12625), .B0_t (SubBytesIns_Inst_Sbox_8_L10), .B0_f (new_AGEMA_signal_12632), .B1_t (new_AGEMA_signal_12633), .B1_f (new_AGEMA_signal_12634), .Z0_t (SubBytesIns_Inst_Sbox_8_L25), .Z0_f (new_AGEMA_signal_13247), .Z1_t (new_AGEMA_signal_13248), .Z1_f (new_AGEMA_signal_13249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L7), .A0_f (new_AGEMA_signal_12626), .A1_t (new_AGEMA_signal_12627), .A1_f (new_AGEMA_signal_12628), .B0_t (SubBytesIns_Inst_Sbox_8_L9), .B0_f (new_AGEMA_signal_12629), .B1_t (new_AGEMA_signal_12630), .B1_f (new_AGEMA_signal_12631), .Z0_t (SubBytesIns_Inst_Sbox_8_L26), .Z0_f (new_AGEMA_signal_13250), .Z1_t (new_AGEMA_signal_13251), .Z1_f (new_AGEMA_signal_13252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L8), .A0_f (new_AGEMA_signal_11438), .A1_t (new_AGEMA_signal_11439), .A1_f (new_AGEMA_signal_11440), .B0_t (SubBytesIns_Inst_Sbox_8_L10), .B0_f (new_AGEMA_signal_12632), .B1_t (new_AGEMA_signal_12633), .B1_f (new_AGEMA_signal_12634), .Z0_t (SubBytesIns_Inst_Sbox_8_L27), .Z0_f (new_AGEMA_signal_13253), .Z1_t (new_AGEMA_signal_13254), .Z1_f (new_AGEMA_signal_13255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L11), .A0_f (new_AGEMA_signal_12635), .A1_t (new_AGEMA_signal_12636), .A1_f (new_AGEMA_signal_12637), .B0_t (SubBytesIns_Inst_Sbox_8_L14), .B0_f (new_AGEMA_signal_12074), .B1_t (new_AGEMA_signal_12075), .B1_f (new_AGEMA_signal_12076), .Z0_t (SubBytesIns_Inst_Sbox_8_L28), .Z0_f (new_AGEMA_signal_13256), .Z1_t (new_AGEMA_signal_13257), .Z1_f (new_AGEMA_signal_13258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L11), .A0_f (new_AGEMA_signal_12635), .A1_t (new_AGEMA_signal_12636), .A1_f (new_AGEMA_signal_12637), .B0_t (SubBytesIns_Inst_Sbox_8_L17), .B0_f (new_AGEMA_signal_12080), .B1_t (new_AGEMA_signal_12081), .B1_f (new_AGEMA_signal_12082), .Z0_t (SubBytesIns_Inst_Sbox_8_L29), .Z0_f (new_AGEMA_signal_13259), .Z1_t (new_AGEMA_signal_13260), .Z1_f (new_AGEMA_signal_13261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L6), .A0_f (new_AGEMA_signal_12623), .A1_t (new_AGEMA_signal_12624), .A1_f (new_AGEMA_signal_12625), .B0_t (SubBytesIns_Inst_Sbox_8_L24), .B0_f (new_AGEMA_signal_13244), .B1_t (new_AGEMA_signal_13245), .B1_f (new_AGEMA_signal_13246), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .Z0_f (new_AGEMA_signal_13808), .Z1_t (new_AGEMA_signal_13809), .Z1_f (new_AGEMA_signal_13810) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L16), .A0_f (new_AGEMA_signal_13235), .A1_t (new_AGEMA_signal_13236), .A1_f (new_AGEMA_signal_13237), .B0_t (SubBytesIns_Inst_Sbox_8_L26), .B0_f (new_AGEMA_signal_13250), .B1_t (new_AGEMA_signal_13251), .B1_f (new_AGEMA_signal_13252), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .Z0_f (new_AGEMA_signal_13811), .Z1_t (new_AGEMA_signal_13812), .Z1_f (new_AGEMA_signal_13813) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L19), .A0_f (new_AGEMA_signal_12638), .A1_t (new_AGEMA_signal_12639), .A1_f (new_AGEMA_signal_12640), .B0_t (SubBytesIns_Inst_Sbox_8_L28), .B0_f (new_AGEMA_signal_13256), .B1_t (new_AGEMA_signal_13257), .B1_f (new_AGEMA_signal_13258), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .Z0_f (new_AGEMA_signal_13814), .Z1_t (new_AGEMA_signal_13815), .Z1_f (new_AGEMA_signal_13816) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L6), .A0_f (new_AGEMA_signal_12623), .A1_t (new_AGEMA_signal_12624), .A1_f (new_AGEMA_signal_12625), .B0_t (SubBytesIns_Inst_Sbox_8_L21), .B0_f (new_AGEMA_signal_13241), .B1_t (new_AGEMA_signal_13242), .B1_f (new_AGEMA_signal_13243), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .Z0_f (new_AGEMA_signal_13817), .Z1_t (new_AGEMA_signal_13818), .Z1_f (new_AGEMA_signal_13819) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L20), .A0_f (new_AGEMA_signal_13238), .A1_t (new_AGEMA_signal_13239), .A1_f (new_AGEMA_signal_13240), .B0_t (SubBytesIns_Inst_Sbox_8_L22), .B0_f (new_AGEMA_signal_12641), .B1_t (new_AGEMA_signal_12642), .B1_f (new_AGEMA_signal_12643), .Z0_t (MixColumnsInput[35]), .Z0_f (new_AGEMA_signal_13820), .Z1_t (new_AGEMA_signal_13821), .Z1_f (new_AGEMA_signal_13822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L25), .A0_f (new_AGEMA_signal_13247), .A1_t (new_AGEMA_signal_13248), .A1_f (new_AGEMA_signal_13249), .B0_t (SubBytesIns_Inst_Sbox_8_L29), .B0_f (new_AGEMA_signal_13259), .B1_t (new_AGEMA_signal_13260), .B1_f (new_AGEMA_signal_13261), .Z0_t (MixColumnsInput[34]), .Z0_f (new_AGEMA_signal_13823), .Z1_t (new_AGEMA_signal_13824), .Z1_f (new_AGEMA_signal_13825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L13), .A0_f (new_AGEMA_signal_13232), .A1_t (new_AGEMA_signal_13233), .A1_f (new_AGEMA_signal_13234), .B0_t (SubBytesIns_Inst_Sbox_8_L27), .B0_f (new_AGEMA_signal_13253), .B1_t (new_AGEMA_signal_13254), .B1_f (new_AGEMA_signal_13255), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .Z0_f (new_AGEMA_signal_13826), .Z1_t (new_AGEMA_signal_13827), .Z1_f (new_AGEMA_signal_13828) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L6), .A0_f (new_AGEMA_signal_12623), .A1_t (new_AGEMA_signal_12624), .A1_f (new_AGEMA_signal_12625), .B0_t (SubBytesIns_Inst_Sbox_8_L23), .B0_f (new_AGEMA_signal_12644), .B1_t (new_AGEMA_signal_12645), .B1_f (new_AGEMA_signal_12646), .Z0_t (MixColumnsInput[32]), .Z0_f (new_AGEMA_signal_13262), .Z1_t (new_AGEMA_signal_13263), .Z1_f (new_AGEMA_signal_13264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[79]), .A0_f (ciphertext_s0_f[79]), .A1_t (ciphertext_s1_t[79]), .A1_f (ciphertext_s1_f[79]), .B0_t (ciphertext_s0_t[76]), .B0_f (ciphertext_s0_f[76]), .B1_t (ciphertext_s1_t[76]), .B1_f (ciphertext_s1_f[76]), .Z0_t (SubBytesIns_Inst_Sbox_9_T1), .Z0_f (new_AGEMA_signal_6616), .Z1_t (new_AGEMA_signal_6617), .Z1_f (new_AGEMA_signal_6618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[79]), .A0_f (ciphertext_s0_f[79]), .A1_t (ciphertext_s1_t[79]), .A1_f (ciphertext_s1_f[79]), .B0_t (ciphertext_s0_t[74]), .B0_f (ciphertext_s0_f[74]), .B1_t (ciphertext_s1_t[74]), .B1_f (ciphertext_s1_f[74]), .Z0_t (SubBytesIns_Inst_Sbox_9_T2), .Z0_f (new_AGEMA_signal_6619), .Z1_t (new_AGEMA_signal_6620), .Z1_f (new_AGEMA_signal_6621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[79]), .A0_f (ciphertext_s0_f[79]), .A1_t (ciphertext_s1_t[79]), .A1_f (ciphertext_s1_f[79]), .B0_t (ciphertext_s0_t[73]), .B0_f (ciphertext_s0_f[73]), .B1_t (ciphertext_s1_t[73]), .B1_f (ciphertext_s1_f[73]), .Z0_t (SubBytesIns_Inst_Sbox_9_T3), .Z0_f (new_AGEMA_signal_6622), .Z1_t (new_AGEMA_signal_6623), .Z1_f (new_AGEMA_signal_6624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[76]), .A0_f (ciphertext_s0_f[76]), .A1_t (ciphertext_s1_t[76]), .A1_f (ciphertext_s1_f[76]), .B0_t (ciphertext_s0_t[74]), .B0_f (ciphertext_s0_f[74]), .B1_t (ciphertext_s1_t[74]), .B1_f (ciphertext_s1_f[74]), .Z0_t (SubBytesIns_Inst_Sbox_9_T4), .Z0_f (new_AGEMA_signal_6625), .Z1_t (new_AGEMA_signal_6626), .Z1_f (new_AGEMA_signal_6627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[75]), .A0_f (ciphertext_s0_f[75]), .A1_t (ciphertext_s1_t[75]), .A1_f (ciphertext_s1_f[75]), .B0_t (ciphertext_s0_t[73]), .B0_f (ciphertext_s0_f[73]), .B1_t (ciphertext_s1_t[73]), .B1_f (ciphertext_s1_f[73]), .Z0_t (SubBytesIns_Inst_Sbox_9_T5), .Z0_f (new_AGEMA_signal_6628), .Z1_t (new_AGEMA_signal_6629), .Z1_f (new_AGEMA_signal_6630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T1), .A0_f (new_AGEMA_signal_6616), .A1_t (new_AGEMA_signal_6617), .A1_f (new_AGEMA_signal_6618), .B0_t (SubBytesIns_Inst_Sbox_9_T5), .B0_f (new_AGEMA_signal_6628), .B1_t (new_AGEMA_signal_6629), .B1_f (new_AGEMA_signal_6630), .Z0_t (SubBytesIns_Inst_Sbox_9_T6), .Z0_f (new_AGEMA_signal_7144), .Z1_t (new_AGEMA_signal_7145), .Z1_f (new_AGEMA_signal_7146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[78]), .A0_f (ciphertext_s0_f[78]), .A1_t (ciphertext_s1_t[78]), .A1_f (ciphertext_s1_f[78]), .B0_t (ciphertext_s0_t[77]), .B0_f (ciphertext_s0_f[77]), .B1_t (ciphertext_s1_t[77]), .B1_f (ciphertext_s1_f[77]), .Z0_t (SubBytesIns_Inst_Sbox_9_T7), .Z0_f (new_AGEMA_signal_6631), .Z1_t (new_AGEMA_signal_6632), .Z1_f (new_AGEMA_signal_6633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[72]), .A0_f (ciphertext_s0_f[72]), .A1_t (ciphertext_s1_t[72]), .A1_f (ciphertext_s1_f[72]), .B0_t (SubBytesIns_Inst_Sbox_9_T6), .B0_f (new_AGEMA_signal_7144), .B1_t (new_AGEMA_signal_7145), .B1_f (new_AGEMA_signal_7146), .Z0_t (SubBytesIns_Inst_Sbox_9_T8), .Z0_f (new_AGEMA_signal_7823), .Z1_t (new_AGEMA_signal_7824), .Z1_f (new_AGEMA_signal_7825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[72]), .A0_f (ciphertext_s0_f[72]), .A1_t (ciphertext_s1_t[72]), .A1_f (ciphertext_s1_f[72]), .B0_t (SubBytesIns_Inst_Sbox_9_T7), .B0_f (new_AGEMA_signal_6631), .B1_t (new_AGEMA_signal_6632), .B1_f (new_AGEMA_signal_6633), .Z0_t (SubBytesIns_Inst_Sbox_9_T9), .Z0_f (new_AGEMA_signal_7147), .Z1_t (new_AGEMA_signal_7148), .Z1_f (new_AGEMA_signal_7149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T6), .A0_f (new_AGEMA_signal_7144), .A1_t (new_AGEMA_signal_7145), .A1_f (new_AGEMA_signal_7146), .B0_t (SubBytesIns_Inst_Sbox_9_T7), .B0_f (new_AGEMA_signal_6631), .B1_t (new_AGEMA_signal_6632), .B1_f (new_AGEMA_signal_6633), .Z0_t (SubBytesIns_Inst_Sbox_9_T10), .Z0_f (new_AGEMA_signal_7826), .Z1_t (new_AGEMA_signal_7827), .Z1_f (new_AGEMA_signal_7828) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[78]), .A0_f (ciphertext_s0_f[78]), .A1_t (ciphertext_s1_t[78]), .A1_f (ciphertext_s1_f[78]), .B0_t (ciphertext_s0_t[74]), .B0_f (ciphertext_s0_f[74]), .B1_t (ciphertext_s1_t[74]), .B1_f (ciphertext_s1_f[74]), .Z0_t (SubBytesIns_Inst_Sbox_9_T11), .Z0_f (new_AGEMA_signal_6634), .Z1_t (new_AGEMA_signal_6635), .Z1_f (new_AGEMA_signal_6636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[77]), .A0_f (ciphertext_s0_f[77]), .A1_t (ciphertext_s1_t[77]), .A1_f (ciphertext_s1_f[77]), .B0_t (ciphertext_s0_t[74]), .B0_f (ciphertext_s0_f[74]), .B1_t (ciphertext_s1_t[74]), .B1_f (ciphertext_s1_f[74]), .Z0_t (SubBytesIns_Inst_Sbox_9_T12), .Z0_f (new_AGEMA_signal_6637), .Z1_t (new_AGEMA_signal_6638), .Z1_f (new_AGEMA_signal_6639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T3), .A0_f (new_AGEMA_signal_6622), .A1_t (new_AGEMA_signal_6623), .A1_f (new_AGEMA_signal_6624), .B0_t (SubBytesIns_Inst_Sbox_9_T4), .B0_f (new_AGEMA_signal_6625), .B1_t (new_AGEMA_signal_6626), .B1_f (new_AGEMA_signal_6627), .Z0_t (SubBytesIns_Inst_Sbox_9_T13), .Z0_f (new_AGEMA_signal_7150), .Z1_t (new_AGEMA_signal_7151), .Z1_f (new_AGEMA_signal_7152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T6), .A0_f (new_AGEMA_signal_7144), .A1_t (new_AGEMA_signal_7145), .A1_f (new_AGEMA_signal_7146), .B0_t (SubBytesIns_Inst_Sbox_9_T11), .B0_f (new_AGEMA_signal_6634), .B1_t (new_AGEMA_signal_6635), .B1_f (new_AGEMA_signal_6636), .Z0_t (SubBytesIns_Inst_Sbox_9_T14), .Z0_f (new_AGEMA_signal_7829), .Z1_t (new_AGEMA_signal_7830), .Z1_f (new_AGEMA_signal_7831) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T5), .A0_f (new_AGEMA_signal_6628), .A1_t (new_AGEMA_signal_6629), .A1_f (new_AGEMA_signal_6630), .B0_t (SubBytesIns_Inst_Sbox_9_T11), .B0_f (new_AGEMA_signal_6634), .B1_t (new_AGEMA_signal_6635), .B1_f (new_AGEMA_signal_6636), .Z0_t (SubBytesIns_Inst_Sbox_9_T15), .Z0_f (new_AGEMA_signal_7153), .Z1_t (new_AGEMA_signal_7154), .Z1_f (new_AGEMA_signal_7155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T5), .A0_f (new_AGEMA_signal_6628), .A1_t (new_AGEMA_signal_6629), .A1_f (new_AGEMA_signal_6630), .B0_t (SubBytesIns_Inst_Sbox_9_T12), .B0_f (new_AGEMA_signal_6637), .B1_t (new_AGEMA_signal_6638), .B1_f (new_AGEMA_signal_6639), .Z0_t (SubBytesIns_Inst_Sbox_9_T16), .Z0_f (new_AGEMA_signal_7156), .Z1_t (new_AGEMA_signal_7157), .Z1_f (new_AGEMA_signal_7158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T9), .A0_f (new_AGEMA_signal_7147), .A1_t (new_AGEMA_signal_7148), .A1_f (new_AGEMA_signal_7149), .B0_t (SubBytesIns_Inst_Sbox_9_T16), .B0_f (new_AGEMA_signal_7156), .B1_t (new_AGEMA_signal_7157), .B1_f (new_AGEMA_signal_7158), .Z0_t (SubBytesIns_Inst_Sbox_9_T17), .Z0_f (new_AGEMA_signal_7832), .Z1_t (new_AGEMA_signal_7833), .Z1_f (new_AGEMA_signal_7834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[76]), .A0_f (ciphertext_s0_f[76]), .A1_t (ciphertext_s1_t[76]), .A1_f (ciphertext_s1_f[76]), .B0_t (ciphertext_s0_t[72]), .B0_f (ciphertext_s0_f[72]), .B1_t (ciphertext_s1_t[72]), .B1_f (ciphertext_s1_f[72]), .Z0_t (SubBytesIns_Inst_Sbox_9_T18), .Z0_f (new_AGEMA_signal_6640), .Z1_t (new_AGEMA_signal_6641), .Z1_f (new_AGEMA_signal_6642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T7), .A0_f (new_AGEMA_signal_6631), .A1_t (new_AGEMA_signal_6632), .A1_f (new_AGEMA_signal_6633), .B0_t (SubBytesIns_Inst_Sbox_9_T18), .B0_f (new_AGEMA_signal_6640), .B1_t (new_AGEMA_signal_6641), .B1_f (new_AGEMA_signal_6642), .Z0_t (SubBytesIns_Inst_Sbox_9_T19), .Z0_f (new_AGEMA_signal_7159), .Z1_t (new_AGEMA_signal_7160), .Z1_f (new_AGEMA_signal_7161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T1), .A0_f (new_AGEMA_signal_6616), .A1_t (new_AGEMA_signal_6617), .A1_f (new_AGEMA_signal_6618), .B0_t (SubBytesIns_Inst_Sbox_9_T19), .B0_f (new_AGEMA_signal_7159), .B1_t (new_AGEMA_signal_7160), .B1_f (new_AGEMA_signal_7161), .Z0_t (SubBytesIns_Inst_Sbox_9_T20), .Z0_f (new_AGEMA_signal_7835), .Z1_t (new_AGEMA_signal_7836), .Z1_f (new_AGEMA_signal_7837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[73]), .A0_f (ciphertext_s0_f[73]), .A1_t (ciphertext_s1_t[73]), .A1_f (ciphertext_s1_f[73]), .B0_t (ciphertext_s0_t[72]), .B0_f (ciphertext_s0_f[72]), .B1_t (ciphertext_s1_t[72]), .B1_f (ciphertext_s1_f[72]), .Z0_t (SubBytesIns_Inst_Sbox_9_T21), .Z0_f (new_AGEMA_signal_6643), .Z1_t (new_AGEMA_signal_6644), .Z1_f (new_AGEMA_signal_6645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T7), .A0_f (new_AGEMA_signal_6631), .A1_t (new_AGEMA_signal_6632), .A1_f (new_AGEMA_signal_6633), .B0_t (SubBytesIns_Inst_Sbox_9_T21), .B0_f (new_AGEMA_signal_6643), .B1_t (new_AGEMA_signal_6644), .B1_f (new_AGEMA_signal_6645), .Z0_t (SubBytesIns_Inst_Sbox_9_T22), .Z0_f (new_AGEMA_signal_7162), .Z1_t (new_AGEMA_signal_7163), .Z1_f (new_AGEMA_signal_7164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T2), .A0_f (new_AGEMA_signal_6619), .A1_t (new_AGEMA_signal_6620), .A1_f (new_AGEMA_signal_6621), .B0_t (SubBytesIns_Inst_Sbox_9_T22), .B0_f (new_AGEMA_signal_7162), .B1_t (new_AGEMA_signal_7163), .B1_f (new_AGEMA_signal_7164), .Z0_t (SubBytesIns_Inst_Sbox_9_T23), .Z0_f (new_AGEMA_signal_7838), .Z1_t (new_AGEMA_signal_7839), .Z1_f (new_AGEMA_signal_7840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T2), .A0_f (new_AGEMA_signal_6619), .A1_t (new_AGEMA_signal_6620), .A1_f (new_AGEMA_signal_6621), .B0_t (SubBytesIns_Inst_Sbox_9_T10), .B0_f (new_AGEMA_signal_7826), .B1_t (new_AGEMA_signal_7827), .B1_f (new_AGEMA_signal_7828), .Z0_t (SubBytesIns_Inst_Sbox_9_T24), .Z0_f (new_AGEMA_signal_8447), .Z1_t (new_AGEMA_signal_8448), .Z1_f (new_AGEMA_signal_8449) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T20), .A0_f (new_AGEMA_signal_7835), .A1_t (new_AGEMA_signal_7836), .A1_f (new_AGEMA_signal_7837), .B0_t (SubBytesIns_Inst_Sbox_9_T17), .B0_f (new_AGEMA_signal_7832), .B1_t (new_AGEMA_signal_7833), .B1_f (new_AGEMA_signal_7834), .Z0_t (SubBytesIns_Inst_Sbox_9_T25), .Z0_f (new_AGEMA_signal_8450), .Z1_t (new_AGEMA_signal_8451), .Z1_f (new_AGEMA_signal_8452) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T3), .A0_f (new_AGEMA_signal_6622), .A1_t (new_AGEMA_signal_6623), .A1_f (new_AGEMA_signal_6624), .B0_t (SubBytesIns_Inst_Sbox_9_T16), .B0_f (new_AGEMA_signal_7156), .B1_t (new_AGEMA_signal_7157), .B1_f (new_AGEMA_signal_7158), .Z0_t (SubBytesIns_Inst_Sbox_9_T26), .Z0_f (new_AGEMA_signal_7841), .Z1_t (new_AGEMA_signal_7842), .Z1_f (new_AGEMA_signal_7843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T1), .A0_f (new_AGEMA_signal_6616), .A1_t (new_AGEMA_signal_6617), .A1_f (new_AGEMA_signal_6618), .B0_t (SubBytesIns_Inst_Sbox_9_T12), .B0_f (new_AGEMA_signal_6637), .B1_t (new_AGEMA_signal_6638), .B1_f (new_AGEMA_signal_6639), .Z0_t (SubBytesIns_Inst_Sbox_9_T27), .Z0_f (new_AGEMA_signal_7165), .Z1_t (new_AGEMA_signal_7166), .Z1_f (new_AGEMA_signal_7167) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T13), .A0_f (new_AGEMA_signal_7150), .A1_t (new_AGEMA_signal_7151), .A1_f (new_AGEMA_signal_7152), .B0_t (SubBytesIns_Inst_Sbox_9_T6), .B0_f (new_AGEMA_signal_7144), .B1_t (new_AGEMA_signal_7145), .B1_f (new_AGEMA_signal_7146), .Z0_t (SubBytesIns_Inst_Sbox_9_M1), .Z0_f (new_AGEMA_signal_7844), .Z1_t (new_AGEMA_signal_7845), .Z1_f (new_AGEMA_signal_7846) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T23), .A0_f (new_AGEMA_signal_7838), .A1_t (new_AGEMA_signal_7839), .A1_f (new_AGEMA_signal_7840), .B0_t (SubBytesIns_Inst_Sbox_9_T8), .B0_f (new_AGEMA_signal_7823), .B1_t (new_AGEMA_signal_7824), .B1_f (new_AGEMA_signal_7825), .Z0_t (SubBytesIns_Inst_Sbox_9_M2), .Z0_f (new_AGEMA_signal_8453), .Z1_t (new_AGEMA_signal_8454), .Z1_f (new_AGEMA_signal_8455) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T14), .A0_f (new_AGEMA_signal_7829), .A1_t (new_AGEMA_signal_7830), .A1_f (new_AGEMA_signal_7831), .B0_t (SubBytesIns_Inst_Sbox_9_M1), .B0_f (new_AGEMA_signal_7844), .B1_t (new_AGEMA_signal_7845), .B1_f (new_AGEMA_signal_7846), .Z0_t (SubBytesIns_Inst_Sbox_9_M3), .Z0_f (new_AGEMA_signal_8456), .Z1_t (new_AGEMA_signal_8457), .Z1_f (new_AGEMA_signal_8458) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T19), .A0_f (new_AGEMA_signal_7159), .A1_t (new_AGEMA_signal_7160), .A1_f (new_AGEMA_signal_7161), .B0_t (ciphertext_s0_t[72]), .B0_f (ciphertext_s0_f[72]), .B1_t (ciphertext_s1_t[72]), .B1_f (ciphertext_s1_f[72]), .Z0_t (SubBytesIns_Inst_Sbox_9_M4), .Z0_f (new_AGEMA_signal_7847), .Z1_t (new_AGEMA_signal_7848), .Z1_f (new_AGEMA_signal_7849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M4), .A0_f (new_AGEMA_signal_7847), .A1_t (new_AGEMA_signal_7848), .A1_f (new_AGEMA_signal_7849), .B0_t (SubBytesIns_Inst_Sbox_9_M1), .B0_f (new_AGEMA_signal_7844), .B1_t (new_AGEMA_signal_7845), .B1_f (new_AGEMA_signal_7846), .Z0_t (SubBytesIns_Inst_Sbox_9_M5), .Z0_f (new_AGEMA_signal_8459), .Z1_t (new_AGEMA_signal_8460), .Z1_f (new_AGEMA_signal_8461) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T3), .A0_f (new_AGEMA_signal_6622), .A1_t (new_AGEMA_signal_6623), .A1_f (new_AGEMA_signal_6624), .B0_t (SubBytesIns_Inst_Sbox_9_T16), .B0_f (new_AGEMA_signal_7156), .B1_t (new_AGEMA_signal_7157), .B1_f (new_AGEMA_signal_7158), .Z0_t (SubBytesIns_Inst_Sbox_9_M6), .Z0_f (new_AGEMA_signal_7850), .Z1_t (new_AGEMA_signal_7851), .Z1_f (new_AGEMA_signal_7852) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T22), .A0_f (new_AGEMA_signal_7162), .A1_t (new_AGEMA_signal_7163), .A1_f (new_AGEMA_signal_7164), .B0_t (SubBytesIns_Inst_Sbox_9_T9), .B0_f (new_AGEMA_signal_7147), .B1_t (new_AGEMA_signal_7148), .B1_f (new_AGEMA_signal_7149), .Z0_t (SubBytesIns_Inst_Sbox_9_M7), .Z0_f (new_AGEMA_signal_7853), .Z1_t (new_AGEMA_signal_7854), .Z1_f (new_AGEMA_signal_7855) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T26), .A0_f (new_AGEMA_signal_7841), .A1_t (new_AGEMA_signal_7842), .A1_f (new_AGEMA_signal_7843), .B0_t (SubBytesIns_Inst_Sbox_9_M6), .B0_f (new_AGEMA_signal_7850), .B1_t (new_AGEMA_signal_7851), .B1_f (new_AGEMA_signal_7852), .Z0_t (SubBytesIns_Inst_Sbox_9_M8), .Z0_f (new_AGEMA_signal_8462), .Z1_t (new_AGEMA_signal_8463), .Z1_f (new_AGEMA_signal_8464) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T20), .A0_f (new_AGEMA_signal_7835), .A1_t (new_AGEMA_signal_7836), .A1_f (new_AGEMA_signal_7837), .B0_t (SubBytesIns_Inst_Sbox_9_T17), .B0_f (new_AGEMA_signal_7832), .B1_t (new_AGEMA_signal_7833), .B1_f (new_AGEMA_signal_7834), .Z0_t (SubBytesIns_Inst_Sbox_9_M9), .Z0_f (new_AGEMA_signal_8465), .Z1_t (new_AGEMA_signal_8466), .Z1_f (new_AGEMA_signal_8467) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M9), .A0_f (new_AGEMA_signal_8465), .A1_t (new_AGEMA_signal_8466), .A1_f (new_AGEMA_signal_8467), .B0_t (SubBytesIns_Inst_Sbox_9_M6), .B0_f (new_AGEMA_signal_7850), .B1_t (new_AGEMA_signal_7851), .B1_f (new_AGEMA_signal_7852), .Z0_t (SubBytesIns_Inst_Sbox_9_M10), .Z0_f (new_AGEMA_signal_8831), .Z1_t (new_AGEMA_signal_8832), .Z1_f (new_AGEMA_signal_8833) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T1), .A0_f (new_AGEMA_signal_6616), .A1_t (new_AGEMA_signal_6617), .A1_f (new_AGEMA_signal_6618), .B0_t (SubBytesIns_Inst_Sbox_9_T15), .B0_f (new_AGEMA_signal_7153), .B1_t (new_AGEMA_signal_7154), .B1_f (new_AGEMA_signal_7155), .Z0_t (SubBytesIns_Inst_Sbox_9_M11), .Z0_f (new_AGEMA_signal_7856), .Z1_t (new_AGEMA_signal_7857), .Z1_f (new_AGEMA_signal_7858) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T4), .A0_f (new_AGEMA_signal_6625), .A1_t (new_AGEMA_signal_6626), .A1_f (new_AGEMA_signal_6627), .B0_t (SubBytesIns_Inst_Sbox_9_T27), .B0_f (new_AGEMA_signal_7165), .B1_t (new_AGEMA_signal_7166), .B1_f (new_AGEMA_signal_7167), .Z0_t (SubBytesIns_Inst_Sbox_9_M12), .Z0_f (new_AGEMA_signal_7859), .Z1_t (new_AGEMA_signal_7860), .Z1_f (new_AGEMA_signal_7861) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M12), .A0_f (new_AGEMA_signal_7859), .A1_t (new_AGEMA_signal_7860), .A1_f (new_AGEMA_signal_7861), .B0_t (SubBytesIns_Inst_Sbox_9_M11), .B0_f (new_AGEMA_signal_7856), .B1_t (new_AGEMA_signal_7857), .B1_f (new_AGEMA_signal_7858), .Z0_t (SubBytesIns_Inst_Sbox_9_M13), .Z0_f (new_AGEMA_signal_8468), .Z1_t (new_AGEMA_signal_8469), .Z1_f (new_AGEMA_signal_8470) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T2), .A0_f (new_AGEMA_signal_6619), .A1_t (new_AGEMA_signal_6620), .A1_f (new_AGEMA_signal_6621), .B0_t (SubBytesIns_Inst_Sbox_9_T10), .B0_f (new_AGEMA_signal_7826), .B1_t (new_AGEMA_signal_7827), .B1_f (new_AGEMA_signal_7828), .Z0_t (SubBytesIns_Inst_Sbox_9_M14), .Z0_f (new_AGEMA_signal_8471), .Z1_t (new_AGEMA_signal_8472), .Z1_f (new_AGEMA_signal_8473) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M14), .A0_f (new_AGEMA_signal_8471), .A1_t (new_AGEMA_signal_8472), .A1_f (new_AGEMA_signal_8473), .B0_t (SubBytesIns_Inst_Sbox_9_M11), .B0_f (new_AGEMA_signal_7856), .B1_t (new_AGEMA_signal_7857), .B1_f (new_AGEMA_signal_7858), .Z0_t (SubBytesIns_Inst_Sbox_9_M15), .Z0_f (new_AGEMA_signal_8834), .Z1_t (new_AGEMA_signal_8835), .Z1_f (new_AGEMA_signal_8836) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M3), .A0_f (new_AGEMA_signal_8456), .A1_t (new_AGEMA_signal_8457), .A1_f (new_AGEMA_signal_8458), .B0_t (SubBytesIns_Inst_Sbox_9_M2), .B0_f (new_AGEMA_signal_8453), .B1_t (new_AGEMA_signal_8454), .B1_f (new_AGEMA_signal_8455), .Z0_t (SubBytesIns_Inst_Sbox_9_M16), .Z0_f (new_AGEMA_signal_8837), .Z1_t (new_AGEMA_signal_8838), .Z1_f (new_AGEMA_signal_8839) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M5), .A0_f (new_AGEMA_signal_8459), .A1_t (new_AGEMA_signal_8460), .A1_f (new_AGEMA_signal_8461), .B0_t (SubBytesIns_Inst_Sbox_9_T24), .B0_f (new_AGEMA_signal_8447), .B1_t (new_AGEMA_signal_8448), .B1_f (new_AGEMA_signal_8449), .Z0_t (SubBytesIns_Inst_Sbox_9_M17), .Z0_f (new_AGEMA_signal_8840), .Z1_t (new_AGEMA_signal_8841), .Z1_f (new_AGEMA_signal_8842) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M8), .A0_f (new_AGEMA_signal_8462), .A1_t (new_AGEMA_signal_8463), .A1_f (new_AGEMA_signal_8464), .B0_t (SubBytesIns_Inst_Sbox_9_M7), .B0_f (new_AGEMA_signal_7853), .B1_t (new_AGEMA_signal_7854), .B1_f (new_AGEMA_signal_7855), .Z0_t (SubBytesIns_Inst_Sbox_9_M18), .Z0_f (new_AGEMA_signal_8843), .Z1_t (new_AGEMA_signal_8844), .Z1_f (new_AGEMA_signal_8845) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M10), .A0_f (new_AGEMA_signal_8831), .A1_t (new_AGEMA_signal_8832), .A1_f (new_AGEMA_signal_8833), .B0_t (SubBytesIns_Inst_Sbox_9_M15), .B0_f (new_AGEMA_signal_8834), .B1_t (new_AGEMA_signal_8835), .B1_f (new_AGEMA_signal_8836), .Z0_t (SubBytesIns_Inst_Sbox_9_M19), .Z0_f (new_AGEMA_signal_9092), .Z1_t (new_AGEMA_signal_9093), .Z1_f (new_AGEMA_signal_9094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M16), .A0_f (new_AGEMA_signal_8837), .A1_t (new_AGEMA_signal_8838), .A1_f (new_AGEMA_signal_8839), .B0_t (SubBytesIns_Inst_Sbox_9_M13), .B0_f (new_AGEMA_signal_8468), .B1_t (new_AGEMA_signal_8469), .B1_f (new_AGEMA_signal_8470), .Z0_t (SubBytesIns_Inst_Sbox_9_M20), .Z0_f (new_AGEMA_signal_9095), .Z1_t (new_AGEMA_signal_9096), .Z1_f (new_AGEMA_signal_9097) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M17), .A0_f (new_AGEMA_signal_8840), .A1_t (new_AGEMA_signal_8841), .A1_f (new_AGEMA_signal_8842), .B0_t (SubBytesIns_Inst_Sbox_9_M15), .B0_f (new_AGEMA_signal_8834), .B1_t (new_AGEMA_signal_8835), .B1_f (new_AGEMA_signal_8836), .Z0_t (SubBytesIns_Inst_Sbox_9_M21), .Z0_f (new_AGEMA_signal_9098), .Z1_t (new_AGEMA_signal_9099), .Z1_f (new_AGEMA_signal_9100) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M18), .A0_f (new_AGEMA_signal_8843), .A1_t (new_AGEMA_signal_8844), .A1_f (new_AGEMA_signal_8845), .B0_t (SubBytesIns_Inst_Sbox_9_M13), .B0_f (new_AGEMA_signal_8468), .B1_t (new_AGEMA_signal_8469), .B1_f (new_AGEMA_signal_8470), .Z0_t (SubBytesIns_Inst_Sbox_9_M22), .Z0_f (new_AGEMA_signal_9101), .Z1_t (new_AGEMA_signal_9102), .Z1_f (new_AGEMA_signal_9103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M19), .A0_f (new_AGEMA_signal_9092), .A1_t (new_AGEMA_signal_9093), .A1_f (new_AGEMA_signal_9094), .B0_t (SubBytesIns_Inst_Sbox_9_T25), .B0_f (new_AGEMA_signal_8450), .B1_t (new_AGEMA_signal_8451), .B1_f (new_AGEMA_signal_8452), .Z0_t (SubBytesIns_Inst_Sbox_9_M23), .Z0_f (new_AGEMA_signal_9332), .Z1_t (new_AGEMA_signal_9333), .Z1_f (new_AGEMA_signal_9334) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M22), .A0_f (new_AGEMA_signal_9101), .A1_t (new_AGEMA_signal_9102), .A1_f (new_AGEMA_signal_9103), .B0_t (SubBytesIns_Inst_Sbox_9_M23), .B0_f (new_AGEMA_signal_9332), .B1_t (new_AGEMA_signal_9333), .B1_f (new_AGEMA_signal_9334), .Z0_t (SubBytesIns_Inst_Sbox_9_M24), .Z0_f (new_AGEMA_signal_9611), .Z1_t (new_AGEMA_signal_9612), .Z1_f (new_AGEMA_signal_9613) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M22), .A0_f (new_AGEMA_signal_9101), .A1_t (new_AGEMA_signal_9102), .A1_f (new_AGEMA_signal_9103), .B0_t (SubBytesIns_Inst_Sbox_9_M20), .B0_f (new_AGEMA_signal_9095), .B1_t (new_AGEMA_signal_9096), .B1_f (new_AGEMA_signal_9097), .Z0_t (SubBytesIns_Inst_Sbox_9_M25), .Z0_f (new_AGEMA_signal_9335), .Z1_t (new_AGEMA_signal_9336), .Z1_f (new_AGEMA_signal_9337) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M21), .A0_f (new_AGEMA_signal_9098), .A1_t (new_AGEMA_signal_9099), .A1_f (new_AGEMA_signal_9100), .B0_t (SubBytesIns_Inst_Sbox_9_M25), .B0_f (new_AGEMA_signal_9335), .B1_t (new_AGEMA_signal_9336), .B1_f (new_AGEMA_signal_9337), .Z0_t (SubBytesIns_Inst_Sbox_9_M26), .Z0_f (new_AGEMA_signal_9614), .Z1_t (new_AGEMA_signal_9615), .Z1_f (new_AGEMA_signal_9616) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M20), .A0_f (new_AGEMA_signal_9095), .A1_t (new_AGEMA_signal_9096), .A1_f (new_AGEMA_signal_9097), .B0_t (SubBytesIns_Inst_Sbox_9_M21), .B0_f (new_AGEMA_signal_9098), .B1_t (new_AGEMA_signal_9099), .B1_f (new_AGEMA_signal_9100), .Z0_t (SubBytesIns_Inst_Sbox_9_M27), .Z0_f (new_AGEMA_signal_9338), .Z1_t (new_AGEMA_signal_9339), .Z1_f (new_AGEMA_signal_9340) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M23), .A0_f (new_AGEMA_signal_9332), .A1_t (new_AGEMA_signal_9333), .A1_f (new_AGEMA_signal_9334), .B0_t (SubBytesIns_Inst_Sbox_9_M25), .B0_f (new_AGEMA_signal_9335), .B1_t (new_AGEMA_signal_9336), .B1_f (new_AGEMA_signal_9337), .Z0_t (SubBytesIns_Inst_Sbox_9_M28), .Z0_f (new_AGEMA_signal_9617), .Z1_t (new_AGEMA_signal_9618), .Z1_f (new_AGEMA_signal_9619) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M28), .A0_f (new_AGEMA_signal_9617), .A1_t (new_AGEMA_signal_9618), .A1_f (new_AGEMA_signal_9619), .B0_t (SubBytesIns_Inst_Sbox_9_M27), .B0_f (new_AGEMA_signal_9338), .B1_t (new_AGEMA_signal_9339), .B1_f (new_AGEMA_signal_9340), .Z0_t (SubBytesIns_Inst_Sbox_9_M29), .Z0_f (new_AGEMA_signal_9911), .Z1_t (new_AGEMA_signal_9912), .Z1_f (new_AGEMA_signal_9913) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M26), .A0_f (new_AGEMA_signal_9614), .A1_t (new_AGEMA_signal_9615), .A1_f (new_AGEMA_signal_9616), .B0_t (SubBytesIns_Inst_Sbox_9_M24), .B0_f (new_AGEMA_signal_9611), .B1_t (new_AGEMA_signal_9612), .B1_f (new_AGEMA_signal_9613), .Z0_t (SubBytesIns_Inst_Sbox_9_M30), .Z0_f (new_AGEMA_signal_9914), .Z1_t (new_AGEMA_signal_9915), .Z1_f (new_AGEMA_signal_9916) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M20), .A0_f (new_AGEMA_signal_9095), .A1_t (new_AGEMA_signal_9096), .A1_f (new_AGEMA_signal_9097), .B0_t (SubBytesIns_Inst_Sbox_9_M23), .B0_f (new_AGEMA_signal_9332), .B1_t (new_AGEMA_signal_9333), .B1_f (new_AGEMA_signal_9334), .Z0_t (SubBytesIns_Inst_Sbox_9_M31), .Z0_f (new_AGEMA_signal_9620), .Z1_t (new_AGEMA_signal_9621), .Z1_f (new_AGEMA_signal_9622) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M27), .A0_f (new_AGEMA_signal_9338), .A1_t (new_AGEMA_signal_9339), .A1_f (new_AGEMA_signal_9340), .B0_t (SubBytesIns_Inst_Sbox_9_M31), .B0_f (new_AGEMA_signal_9620), .B1_t (new_AGEMA_signal_9621), .B1_f (new_AGEMA_signal_9622), .Z0_t (SubBytesIns_Inst_Sbox_9_M32), .Z0_f (new_AGEMA_signal_9917), .Z1_t (new_AGEMA_signal_9918), .Z1_f (new_AGEMA_signal_9919) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M27), .A0_f (new_AGEMA_signal_9338), .A1_t (new_AGEMA_signal_9339), .A1_f (new_AGEMA_signal_9340), .B0_t (SubBytesIns_Inst_Sbox_9_M25), .B0_f (new_AGEMA_signal_9335), .B1_t (new_AGEMA_signal_9336), .B1_f (new_AGEMA_signal_9337), .Z0_t (SubBytesIns_Inst_Sbox_9_M33), .Z0_f (new_AGEMA_signal_9623), .Z1_t (new_AGEMA_signal_9624), .Z1_f (new_AGEMA_signal_9625) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M21), .A0_f (new_AGEMA_signal_9098), .A1_t (new_AGEMA_signal_9099), .A1_f (new_AGEMA_signal_9100), .B0_t (SubBytesIns_Inst_Sbox_9_M22), .B0_f (new_AGEMA_signal_9101), .B1_t (new_AGEMA_signal_9102), .B1_f (new_AGEMA_signal_9103), .Z0_t (SubBytesIns_Inst_Sbox_9_M34), .Z0_f (new_AGEMA_signal_9341), .Z1_t (new_AGEMA_signal_9342), .Z1_f (new_AGEMA_signal_9343) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M24), .A0_f (new_AGEMA_signal_9611), .A1_t (new_AGEMA_signal_9612), .A1_f (new_AGEMA_signal_9613), .B0_t (SubBytesIns_Inst_Sbox_9_M34), .B0_f (new_AGEMA_signal_9341), .B1_t (new_AGEMA_signal_9342), .B1_f (new_AGEMA_signal_9343), .Z0_t (SubBytesIns_Inst_Sbox_9_M35), .Z0_f (new_AGEMA_signal_9920), .Z1_t (new_AGEMA_signal_9921), .Z1_f (new_AGEMA_signal_9922) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M24), .A0_f (new_AGEMA_signal_9611), .A1_t (new_AGEMA_signal_9612), .A1_f (new_AGEMA_signal_9613), .B0_t (SubBytesIns_Inst_Sbox_9_M25), .B0_f (new_AGEMA_signal_9335), .B1_t (new_AGEMA_signal_9336), .B1_f (new_AGEMA_signal_9337), .Z0_t (SubBytesIns_Inst_Sbox_9_M36), .Z0_f (new_AGEMA_signal_9923), .Z1_t (new_AGEMA_signal_9924), .Z1_f (new_AGEMA_signal_9925) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M21), .A0_f (new_AGEMA_signal_9098), .A1_t (new_AGEMA_signal_9099), .A1_f (new_AGEMA_signal_9100), .B0_t (SubBytesIns_Inst_Sbox_9_M29), .B0_f (new_AGEMA_signal_9911), .B1_t (new_AGEMA_signal_9912), .B1_f (new_AGEMA_signal_9913), .Z0_t (SubBytesIns_Inst_Sbox_9_M37), .Z0_f (new_AGEMA_signal_10172), .Z1_t (new_AGEMA_signal_10173), .Z1_f (new_AGEMA_signal_10174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M32), .A0_f (new_AGEMA_signal_9917), .A1_t (new_AGEMA_signal_9918), .A1_f (new_AGEMA_signal_9919), .B0_t (SubBytesIns_Inst_Sbox_9_M33), .B0_f (new_AGEMA_signal_9623), .B1_t (new_AGEMA_signal_9624), .B1_f (new_AGEMA_signal_9625), .Z0_t (SubBytesIns_Inst_Sbox_9_M38), .Z0_f (new_AGEMA_signal_10175), .Z1_t (new_AGEMA_signal_10176), .Z1_f (new_AGEMA_signal_10177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M23), .A0_f (new_AGEMA_signal_9332), .A1_t (new_AGEMA_signal_9333), .A1_f (new_AGEMA_signal_9334), .B0_t (SubBytesIns_Inst_Sbox_9_M30), .B0_f (new_AGEMA_signal_9914), .B1_t (new_AGEMA_signal_9915), .B1_f (new_AGEMA_signal_9916), .Z0_t (SubBytesIns_Inst_Sbox_9_M39), .Z0_f (new_AGEMA_signal_10178), .Z1_t (new_AGEMA_signal_10179), .Z1_f (new_AGEMA_signal_10180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M35), .A0_f (new_AGEMA_signal_9920), .A1_t (new_AGEMA_signal_9921), .A1_f (new_AGEMA_signal_9922), .B0_t (SubBytesIns_Inst_Sbox_9_M36), .B0_f (new_AGEMA_signal_9923), .B1_t (new_AGEMA_signal_9924), .B1_f (new_AGEMA_signal_9925), .Z0_t (SubBytesIns_Inst_Sbox_9_M40), .Z0_f (new_AGEMA_signal_10181), .Z1_t (new_AGEMA_signal_10182), .Z1_f (new_AGEMA_signal_10183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M38), .A0_f (new_AGEMA_signal_10175), .A1_t (new_AGEMA_signal_10176), .A1_f (new_AGEMA_signal_10177), .B0_t (SubBytesIns_Inst_Sbox_9_M40), .B0_f (new_AGEMA_signal_10181), .B1_t (new_AGEMA_signal_10182), .B1_f (new_AGEMA_signal_10183), .Z0_t (SubBytesIns_Inst_Sbox_9_M41), .Z0_f (new_AGEMA_signal_10724), .Z1_t (new_AGEMA_signal_10725), .Z1_f (new_AGEMA_signal_10726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M37), .A0_f (new_AGEMA_signal_10172), .A1_t (new_AGEMA_signal_10173), .A1_f (new_AGEMA_signal_10174), .B0_t (SubBytesIns_Inst_Sbox_9_M39), .B0_f (new_AGEMA_signal_10178), .B1_t (new_AGEMA_signal_10179), .B1_f (new_AGEMA_signal_10180), .Z0_t (SubBytesIns_Inst_Sbox_9_M42), .Z0_f (new_AGEMA_signal_10727), .Z1_t (new_AGEMA_signal_10728), .Z1_f (new_AGEMA_signal_10729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M37), .A0_f (new_AGEMA_signal_10172), .A1_t (new_AGEMA_signal_10173), .A1_f (new_AGEMA_signal_10174), .B0_t (SubBytesIns_Inst_Sbox_9_M38), .B0_f (new_AGEMA_signal_10175), .B1_t (new_AGEMA_signal_10176), .B1_f (new_AGEMA_signal_10177), .Z0_t (SubBytesIns_Inst_Sbox_9_M43), .Z0_f (new_AGEMA_signal_10730), .Z1_t (new_AGEMA_signal_10731), .Z1_f (new_AGEMA_signal_10732) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M39), .A0_f (new_AGEMA_signal_10178), .A1_t (new_AGEMA_signal_10179), .A1_f (new_AGEMA_signal_10180), .B0_t (SubBytesIns_Inst_Sbox_9_M40), .B0_f (new_AGEMA_signal_10181), .B1_t (new_AGEMA_signal_10182), .B1_f (new_AGEMA_signal_10183), .Z0_t (SubBytesIns_Inst_Sbox_9_M44), .Z0_f (new_AGEMA_signal_10733), .Z1_t (new_AGEMA_signal_10734), .Z1_f (new_AGEMA_signal_10735) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M42), .A0_f (new_AGEMA_signal_10727), .A1_t (new_AGEMA_signal_10728), .A1_f (new_AGEMA_signal_10729), .B0_t (SubBytesIns_Inst_Sbox_9_M41), .B0_f (new_AGEMA_signal_10724), .B1_t (new_AGEMA_signal_10725), .B1_f (new_AGEMA_signal_10726), .Z0_t (SubBytesIns_Inst_Sbox_9_M45), .Z0_f (new_AGEMA_signal_11444), .Z1_t (new_AGEMA_signal_11445), .Z1_f (new_AGEMA_signal_11446) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M44), .A0_f (new_AGEMA_signal_10733), .A1_t (new_AGEMA_signal_10734), .A1_f (new_AGEMA_signal_10735), .B0_t (SubBytesIns_Inst_Sbox_9_T6), .B0_f (new_AGEMA_signal_7144), .B1_t (new_AGEMA_signal_7145), .B1_f (new_AGEMA_signal_7146), .Z0_t (SubBytesIns_Inst_Sbox_9_M46), .Z0_f (new_AGEMA_signal_11447), .Z1_t (new_AGEMA_signal_11448), .Z1_f (new_AGEMA_signal_11449) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M40), .A0_f (new_AGEMA_signal_10181), .A1_t (new_AGEMA_signal_10182), .A1_f (new_AGEMA_signal_10183), .B0_t (SubBytesIns_Inst_Sbox_9_T8), .B0_f (new_AGEMA_signal_7823), .B1_t (new_AGEMA_signal_7824), .B1_f (new_AGEMA_signal_7825), .Z0_t (SubBytesIns_Inst_Sbox_9_M47), .Z0_f (new_AGEMA_signal_10736), .Z1_t (new_AGEMA_signal_10737), .Z1_f (new_AGEMA_signal_10738) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M39), .A0_f (new_AGEMA_signal_10178), .A1_t (new_AGEMA_signal_10179), .A1_f (new_AGEMA_signal_10180), .B0_t (ciphertext_s0_t[72]), .B0_f (ciphertext_s0_f[72]), .B1_t (ciphertext_s1_t[72]), .B1_f (ciphertext_s1_f[72]), .Z0_t (SubBytesIns_Inst_Sbox_9_M48), .Z0_f (new_AGEMA_signal_10739), .Z1_t (new_AGEMA_signal_10740), .Z1_f (new_AGEMA_signal_10741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M43), .A0_f (new_AGEMA_signal_10730), .A1_t (new_AGEMA_signal_10731), .A1_f (new_AGEMA_signal_10732), .B0_t (SubBytesIns_Inst_Sbox_9_T16), .B0_f (new_AGEMA_signal_7156), .B1_t (new_AGEMA_signal_7157), .B1_f (new_AGEMA_signal_7158), .Z0_t (SubBytesIns_Inst_Sbox_9_M49), .Z0_f (new_AGEMA_signal_11450), .Z1_t (new_AGEMA_signal_11451), .Z1_f (new_AGEMA_signal_11452) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M38), .A0_f (new_AGEMA_signal_10175), .A1_t (new_AGEMA_signal_10176), .A1_f (new_AGEMA_signal_10177), .B0_t (SubBytesIns_Inst_Sbox_9_T9), .B0_f (new_AGEMA_signal_7147), .B1_t (new_AGEMA_signal_7148), .B1_f (new_AGEMA_signal_7149), .Z0_t (SubBytesIns_Inst_Sbox_9_M50), .Z0_f (new_AGEMA_signal_10742), .Z1_t (new_AGEMA_signal_10743), .Z1_f (new_AGEMA_signal_10744) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M37), .A0_f (new_AGEMA_signal_10172), .A1_t (new_AGEMA_signal_10173), .A1_f (new_AGEMA_signal_10174), .B0_t (SubBytesIns_Inst_Sbox_9_T17), .B0_f (new_AGEMA_signal_7832), .B1_t (new_AGEMA_signal_7833), .B1_f (new_AGEMA_signal_7834), .Z0_t (SubBytesIns_Inst_Sbox_9_M51), .Z0_f (new_AGEMA_signal_10745), .Z1_t (new_AGEMA_signal_10746), .Z1_f (new_AGEMA_signal_10747) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M42), .A0_f (new_AGEMA_signal_10727), .A1_t (new_AGEMA_signal_10728), .A1_f (new_AGEMA_signal_10729), .B0_t (SubBytesIns_Inst_Sbox_9_T15), .B0_f (new_AGEMA_signal_7153), .B1_t (new_AGEMA_signal_7154), .B1_f (new_AGEMA_signal_7155), .Z0_t (SubBytesIns_Inst_Sbox_9_M52), .Z0_f (new_AGEMA_signal_11453), .Z1_t (new_AGEMA_signal_11454), .Z1_f (new_AGEMA_signal_11455) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M45), .A0_f (new_AGEMA_signal_11444), .A1_t (new_AGEMA_signal_11445), .A1_f (new_AGEMA_signal_11446), .B0_t (SubBytesIns_Inst_Sbox_9_T27), .B0_f (new_AGEMA_signal_7165), .B1_t (new_AGEMA_signal_7166), .B1_f (new_AGEMA_signal_7167), .Z0_t (SubBytesIns_Inst_Sbox_9_M53), .Z0_f (new_AGEMA_signal_12086), .Z1_t (new_AGEMA_signal_12087), .Z1_f (new_AGEMA_signal_12088) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M41), .A0_f (new_AGEMA_signal_10724), .A1_t (new_AGEMA_signal_10725), .A1_f (new_AGEMA_signal_10726), .B0_t (SubBytesIns_Inst_Sbox_9_T10), .B0_f (new_AGEMA_signal_7826), .B1_t (new_AGEMA_signal_7827), .B1_f (new_AGEMA_signal_7828), .Z0_t (SubBytesIns_Inst_Sbox_9_M54), .Z0_f (new_AGEMA_signal_11456), .Z1_t (new_AGEMA_signal_11457), .Z1_f (new_AGEMA_signal_11458) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M44), .A0_f (new_AGEMA_signal_10733), .A1_t (new_AGEMA_signal_10734), .A1_f (new_AGEMA_signal_10735), .B0_t (SubBytesIns_Inst_Sbox_9_T13), .B0_f (new_AGEMA_signal_7150), .B1_t (new_AGEMA_signal_7151), .B1_f (new_AGEMA_signal_7152), .Z0_t (SubBytesIns_Inst_Sbox_9_M55), .Z0_f (new_AGEMA_signal_11459), .Z1_t (new_AGEMA_signal_11460), .Z1_f (new_AGEMA_signal_11461) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M40), .A0_f (new_AGEMA_signal_10181), .A1_t (new_AGEMA_signal_10182), .A1_f (new_AGEMA_signal_10183), .B0_t (SubBytesIns_Inst_Sbox_9_T23), .B0_f (new_AGEMA_signal_7838), .B1_t (new_AGEMA_signal_7839), .B1_f (new_AGEMA_signal_7840), .Z0_t (SubBytesIns_Inst_Sbox_9_M56), .Z0_f (new_AGEMA_signal_10748), .Z1_t (new_AGEMA_signal_10749), .Z1_f (new_AGEMA_signal_10750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M39), .A0_f (new_AGEMA_signal_10178), .A1_t (new_AGEMA_signal_10179), .A1_f (new_AGEMA_signal_10180), .B0_t (SubBytesIns_Inst_Sbox_9_T19), .B0_f (new_AGEMA_signal_7159), .B1_t (new_AGEMA_signal_7160), .B1_f (new_AGEMA_signal_7161), .Z0_t (SubBytesIns_Inst_Sbox_9_M57), .Z0_f (new_AGEMA_signal_10751), .Z1_t (new_AGEMA_signal_10752), .Z1_f (new_AGEMA_signal_10753) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M43), .A0_f (new_AGEMA_signal_10730), .A1_t (new_AGEMA_signal_10731), .A1_f (new_AGEMA_signal_10732), .B0_t (SubBytesIns_Inst_Sbox_9_T3), .B0_f (new_AGEMA_signal_6622), .B1_t (new_AGEMA_signal_6623), .B1_f (new_AGEMA_signal_6624), .Z0_t (SubBytesIns_Inst_Sbox_9_M58), .Z0_f (new_AGEMA_signal_11462), .Z1_t (new_AGEMA_signal_11463), .Z1_f (new_AGEMA_signal_11464) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M38), .A0_f (new_AGEMA_signal_10175), .A1_t (new_AGEMA_signal_10176), .A1_f (new_AGEMA_signal_10177), .B0_t (SubBytesIns_Inst_Sbox_9_T22), .B0_f (new_AGEMA_signal_7162), .B1_t (new_AGEMA_signal_7163), .B1_f (new_AGEMA_signal_7164), .Z0_t (SubBytesIns_Inst_Sbox_9_M59), .Z0_f (new_AGEMA_signal_10754), .Z1_t (new_AGEMA_signal_10755), .Z1_f (new_AGEMA_signal_10756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M37), .A0_f (new_AGEMA_signal_10172), .A1_t (new_AGEMA_signal_10173), .A1_f (new_AGEMA_signal_10174), .B0_t (SubBytesIns_Inst_Sbox_9_T20), .B0_f (new_AGEMA_signal_7835), .B1_t (new_AGEMA_signal_7836), .B1_f (new_AGEMA_signal_7837), .Z0_t (SubBytesIns_Inst_Sbox_9_M60), .Z0_f (new_AGEMA_signal_10757), .Z1_t (new_AGEMA_signal_10758), .Z1_f (new_AGEMA_signal_10759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M42), .A0_f (new_AGEMA_signal_10727), .A1_t (new_AGEMA_signal_10728), .A1_f (new_AGEMA_signal_10729), .B0_t (SubBytesIns_Inst_Sbox_9_T1), .B0_f (new_AGEMA_signal_6616), .B1_t (new_AGEMA_signal_6617), .B1_f (new_AGEMA_signal_6618), .Z0_t (SubBytesIns_Inst_Sbox_9_M61), .Z0_f (new_AGEMA_signal_11465), .Z1_t (new_AGEMA_signal_11466), .Z1_f (new_AGEMA_signal_11467) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M45), .A0_f (new_AGEMA_signal_11444), .A1_t (new_AGEMA_signal_11445), .A1_f (new_AGEMA_signal_11446), .B0_t (SubBytesIns_Inst_Sbox_9_T4), .B0_f (new_AGEMA_signal_6625), .B1_t (new_AGEMA_signal_6626), .B1_f (new_AGEMA_signal_6627), .Z0_t (SubBytesIns_Inst_Sbox_9_M62), .Z0_f (new_AGEMA_signal_12089), .Z1_t (new_AGEMA_signal_12090), .Z1_f (new_AGEMA_signal_12091) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M41), .A0_f (new_AGEMA_signal_10724), .A1_t (new_AGEMA_signal_10725), .A1_f (new_AGEMA_signal_10726), .B0_t (SubBytesIns_Inst_Sbox_9_T2), .B0_f (new_AGEMA_signal_6619), .B1_t (new_AGEMA_signal_6620), .B1_f (new_AGEMA_signal_6621), .Z0_t (SubBytesIns_Inst_Sbox_9_M63), .Z0_f (new_AGEMA_signal_11468), .Z1_t (new_AGEMA_signal_11469), .Z1_f (new_AGEMA_signal_11470) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M61), .A0_f (new_AGEMA_signal_11465), .A1_t (new_AGEMA_signal_11466), .A1_f (new_AGEMA_signal_11467), .B0_t (SubBytesIns_Inst_Sbox_9_M62), .B0_f (new_AGEMA_signal_12089), .B1_t (new_AGEMA_signal_12090), .B1_f (new_AGEMA_signal_12091), .Z0_t (SubBytesIns_Inst_Sbox_9_L0), .Z0_f (new_AGEMA_signal_12647), .Z1_t (new_AGEMA_signal_12648), .Z1_f (new_AGEMA_signal_12649) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M50), .A0_f (new_AGEMA_signal_10742), .A1_t (new_AGEMA_signal_10743), .A1_f (new_AGEMA_signal_10744), .B0_t (SubBytesIns_Inst_Sbox_9_M56), .B0_f (new_AGEMA_signal_10748), .B1_t (new_AGEMA_signal_10749), .B1_f (new_AGEMA_signal_10750), .Z0_t (SubBytesIns_Inst_Sbox_9_L1), .Z0_f (new_AGEMA_signal_11471), .Z1_t (new_AGEMA_signal_11472), .Z1_f (new_AGEMA_signal_11473) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M46), .A0_f (new_AGEMA_signal_11447), .A1_t (new_AGEMA_signal_11448), .A1_f (new_AGEMA_signal_11449), .B0_t (SubBytesIns_Inst_Sbox_9_M48), .B0_f (new_AGEMA_signal_10739), .B1_t (new_AGEMA_signal_10740), .B1_f (new_AGEMA_signal_10741), .Z0_t (SubBytesIns_Inst_Sbox_9_L2), .Z0_f (new_AGEMA_signal_12092), .Z1_t (new_AGEMA_signal_12093), .Z1_f (new_AGEMA_signal_12094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M47), .A0_f (new_AGEMA_signal_10736), .A1_t (new_AGEMA_signal_10737), .A1_f (new_AGEMA_signal_10738), .B0_t (SubBytesIns_Inst_Sbox_9_M55), .B0_f (new_AGEMA_signal_11459), .B1_t (new_AGEMA_signal_11460), .B1_f (new_AGEMA_signal_11461), .Z0_t (SubBytesIns_Inst_Sbox_9_L3), .Z0_f (new_AGEMA_signal_12095), .Z1_t (new_AGEMA_signal_12096), .Z1_f (new_AGEMA_signal_12097) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M54), .A0_f (new_AGEMA_signal_11456), .A1_t (new_AGEMA_signal_11457), .A1_f (new_AGEMA_signal_11458), .B0_t (SubBytesIns_Inst_Sbox_9_M58), .B0_f (new_AGEMA_signal_11462), .B1_t (new_AGEMA_signal_11463), .B1_f (new_AGEMA_signal_11464), .Z0_t (SubBytesIns_Inst_Sbox_9_L4), .Z0_f (new_AGEMA_signal_12098), .Z1_t (new_AGEMA_signal_12099), .Z1_f (new_AGEMA_signal_12100) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M49), .A0_f (new_AGEMA_signal_11450), .A1_t (new_AGEMA_signal_11451), .A1_f (new_AGEMA_signal_11452), .B0_t (SubBytesIns_Inst_Sbox_9_M61), .B0_f (new_AGEMA_signal_11465), .B1_t (new_AGEMA_signal_11466), .B1_f (new_AGEMA_signal_11467), .Z0_t (SubBytesIns_Inst_Sbox_9_L5), .Z0_f (new_AGEMA_signal_12101), .Z1_t (new_AGEMA_signal_12102), .Z1_f (new_AGEMA_signal_12103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M62), .A0_f (new_AGEMA_signal_12089), .A1_t (new_AGEMA_signal_12090), .A1_f (new_AGEMA_signal_12091), .B0_t (SubBytesIns_Inst_Sbox_9_L5), .B0_f (new_AGEMA_signal_12101), .B1_t (new_AGEMA_signal_12102), .B1_f (new_AGEMA_signal_12103), .Z0_t (SubBytesIns_Inst_Sbox_9_L6), .Z0_f (new_AGEMA_signal_12650), .Z1_t (new_AGEMA_signal_12651), .Z1_f (new_AGEMA_signal_12652) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M46), .A0_f (new_AGEMA_signal_11447), .A1_t (new_AGEMA_signal_11448), .A1_f (new_AGEMA_signal_11449), .B0_t (SubBytesIns_Inst_Sbox_9_L3), .B0_f (new_AGEMA_signal_12095), .B1_t (new_AGEMA_signal_12096), .B1_f (new_AGEMA_signal_12097), .Z0_t (SubBytesIns_Inst_Sbox_9_L7), .Z0_f (new_AGEMA_signal_12653), .Z1_t (new_AGEMA_signal_12654), .Z1_f (new_AGEMA_signal_12655) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M51), .A0_f (new_AGEMA_signal_10745), .A1_t (new_AGEMA_signal_10746), .A1_f (new_AGEMA_signal_10747), .B0_t (SubBytesIns_Inst_Sbox_9_M59), .B0_f (new_AGEMA_signal_10754), .B1_t (new_AGEMA_signal_10755), .B1_f (new_AGEMA_signal_10756), .Z0_t (SubBytesIns_Inst_Sbox_9_L8), .Z0_f (new_AGEMA_signal_11474), .Z1_t (new_AGEMA_signal_11475), .Z1_f (new_AGEMA_signal_11476) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M52), .A0_f (new_AGEMA_signal_11453), .A1_t (new_AGEMA_signal_11454), .A1_f (new_AGEMA_signal_11455), .B0_t (SubBytesIns_Inst_Sbox_9_M53), .B0_f (new_AGEMA_signal_12086), .B1_t (new_AGEMA_signal_12087), .B1_f (new_AGEMA_signal_12088), .Z0_t (SubBytesIns_Inst_Sbox_9_L9), .Z0_f (new_AGEMA_signal_12656), .Z1_t (new_AGEMA_signal_12657), .Z1_f (new_AGEMA_signal_12658) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M53), .A0_f (new_AGEMA_signal_12086), .A1_t (new_AGEMA_signal_12087), .A1_f (new_AGEMA_signal_12088), .B0_t (SubBytesIns_Inst_Sbox_9_L4), .B0_f (new_AGEMA_signal_12098), .B1_t (new_AGEMA_signal_12099), .B1_f (new_AGEMA_signal_12100), .Z0_t (SubBytesIns_Inst_Sbox_9_L10), .Z0_f (new_AGEMA_signal_12659), .Z1_t (new_AGEMA_signal_12660), .Z1_f (new_AGEMA_signal_12661) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M60), .A0_f (new_AGEMA_signal_10757), .A1_t (new_AGEMA_signal_10758), .A1_f (new_AGEMA_signal_10759), .B0_t (SubBytesIns_Inst_Sbox_9_L2), .B0_f (new_AGEMA_signal_12092), .B1_t (new_AGEMA_signal_12093), .B1_f (new_AGEMA_signal_12094), .Z0_t (SubBytesIns_Inst_Sbox_9_L11), .Z0_f (new_AGEMA_signal_12662), .Z1_t (new_AGEMA_signal_12663), .Z1_f (new_AGEMA_signal_12664) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M48), .A0_f (new_AGEMA_signal_10739), .A1_t (new_AGEMA_signal_10740), .A1_f (new_AGEMA_signal_10741), .B0_t (SubBytesIns_Inst_Sbox_9_M51), .B0_f (new_AGEMA_signal_10745), .B1_t (new_AGEMA_signal_10746), .B1_f (new_AGEMA_signal_10747), .Z0_t (SubBytesIns_Inst_Sbox_9_L12), .Z0_f (new_AGEMA_signal_11477), .Z1_t (new_AGEMA_signal_11478), .Z1_f (new_AGEMA_signal_11479) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M50), .A0_f (new_AGEMA_signal_10742), .A1_t (new_AGEMA_signal_10743), .A1_f (new_AGEMA_signal_10744), .B0_t (SubBytesIns_Inst_Sbox_9_L0), .B0_f (new_AGEMA_signal_12647), .B1_t (new_AGEMA_signal_12648), .B1_f (new_AGEMA_signal_12649), .Z0_t (SubBytesIns_Inst_Sbox_9_L13), .Z0_f (new_AGEMA_signal_13265), .Z1_t (new_AGEMA_signal_13266), .Z1_f (new_AGEMA_signal_13267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M52), .A0_f (new_AGEMA_signal_11453), .A1_t (new_AGEMA_signal_11454), .A1_f (new_AGEMA_signal_11455), .B0_t (SubBytesIns_Inst_Sbox_9_M61), .B0_f (new_AGEMA_signal_11465), .B1_t (new_AGEMA_signal_11466), .B1_f (new_AGEMA_signal_11467), .Z0_t (SubBytesIns_Inst_Sbox_9_L14), .Z0_f (new_AGEMA_signal_12104), .Z1_t (new_AGEMA_signal_12105), .Z1_f (new_AGEMA_signal_12106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M55), .A0_f (new_AGEMA_signal_11459), .A1_t (new_AGEMA_signal_11460), .A1_f (new_AGEMA_signal_11461), .B0_t (SubBytesIns_Inst_Sbox_9_L1), .B0_f (new_AGEMA_signal_11471), .B1_t (new_AGEMA_signal_11472), .B1_f (new_AGEMA_signal_11473), .Z0_t (SubBytesIns_Inst_Sbox_9_L15), .Z0_f (new_AGEMA_signal_12107), .Z1_t (new_AGEMA_signal_12108), .Z1_f (new_AGEMA_signal_12109) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M56), .A0_f (new_AGEMA_signal_10748), .A1_t (new_AGEMA_signal_10749), .A1_f (new_AGEMA_signal_10750), .B0_t (SubBytesIns_Inst_Sbox_9_L0), .B0_f (new_AGEMA_signal_12647), .B1_t (new_AGEMA_signal_12648), .B1_f (new_AGEMA_signal_12649), .Z0_t (SubBytesIns_Inst_Sbox_9_L16), .Z0_f (new_AGEMA_signal_13268), .Z1_t (new_AGEMA_signal_13269), .Z1_f (new_AGEMA_signal_13270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M57), .A0_f (new_AGEMA_signal_10751), .A1_t (new_AGEMA_signal_10752), .A1_f (new_AGEMA_signal_10753), .B0_t (SubBytesIns_Inst_Sbox_9_L1), .B0_f (new_AGEMA_signal_11471), .B1_t (new_AGEMA_signal_11472), .B1_f (new_AGEMA_signal_11473), .Z0_t (SubBytesIns_Inst_Sbox_9_L17), .Z0_f (new_AGEMA_signal_12110), .Z1_t (new_AGEMA_signal_12111), .Z1_f (new_AGEMA_signal_12112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M58), .A0_f (new_AGEMA_signal_11462), .A1_t (new_AGEMA_signal_11463), .A1_f (new_AGEMA_signal_11464), .B0_t (SubBytesIns_Inst_Sbox_9_L8), .B0_f (new_AGEMA_signal_11474), .B1_t (new_AGEMA_signal_11475), .B1_f (new_AGEMA_signal_11476), .Z0_t (SubBytesIns_Inst_Sbox_9_L18), .Z0_f (new_AGEMA_signal_12113), .Z1_t (new_AGEMA_signal_12114), .Z1_f (new_AGEMA_signal_12115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M63), .A0_f (new_AGEMA_signal_11468), .A1_t (new_AGEMA_signal_11469), .A1_f (new_AGEMA_signal_11470), .B0_t (SubBytesIns_Inst_Sbox_9_L4), .B0_f (new_AGEMA_signal_12098), .B1_t (new_AGEMA_signal_12099), .B1_f (new_AGEMA_signal_12100), .Z0_t (SubBytesIns_Inst_Sbox_9_L19), .Z0_f (new_AGEMA_signal_12665), .Z1_t (new_AGEMA_signal_12666), .Z1_f (new_AGEMA_signal_12667) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L0), .A0_f (new_AGEMA_signal_12647), .A1_t (new_AGEMA_signal_12648), .A1_f (new_AGEMA_signal_12649), .B0_t (SubBytesIns_Inst_Sbox_9_L1), .B0_f (new_AGEMA_signal_11471), .B1_t (new_AGEMA_signal_11472), .B1_f (new_AGEMA_signal_11473), .Z0_t (SubBytesIns_Inst_Sbox_9_L20), .Z0_f (new_AGEMA_signal_13271), .Z1_t (new_AGEMA_signal_13272), .Z1_f (new_AGEMA_signal_13273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L1), .A0_f (new_AGEMA_signal_11471), .A1_t (new_AGEMA_signal_11472), .A1_f (new_AGEMA_signal_11473), .B0_t (SubBytesIns_Inst_Sbox_9_L7), .B0_f (new_AGEMA_signal_12653), .B1_t (new_AGEMA_signal_12654), .B1_f (new_AGEMA_signal_12655), .Z0_t (SubBytesIns_Inst_Sbox_9_L21), .Z0_f (new_AGEMA_signal_13274), .Z1_t (new_AGEMA_signal_13275), .Z1_f (new_AGEMA_signal_13276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L3), .A0_f (new_AGEMA_signal_12095), .A1_t (new_AGEMA_signal_12096), .A1_f (new_AGEMA_signal_12097), .B0_t (SubBytesIns_Inst_Sbox_9_L12), .B0_f (new_AGEMA_signal_11477), .B1_t (new_AGEMA_signal_11478), .B1_f (new_AGEMA_signal_11479), .Z0_t (SubBytesIns_Inst_Sbox_9_L22), .Z0_f (new_AGEMA_signal_12668), .Z1_t (new_AGEMA_signal_12669), .Z1_f (new_AGEMA_signal_12670) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L18), .A0_f (new_AGEMA_signal_12113), .A1_t (new_AGEMA_signal_12114), .A1_f (new_AGEMA_signal_12115), .B0_t (SubBytesIns_Inst_Sbox_9_L2), .B0_f (new_AGEMA_signal_12092), .B1_t (new_AGEMA_signal_12093), .B1_f (new_AGEMA_signal_12094), .Z0_t (SubBytesIns_Inst_Sbox_9_L23), .Z0_f (new_AGEMA_signal_12671), .Z1_t (new_AGEMA_signal_12672), .Z1_f (new_AGEMA_signal_12673) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L15), .A0_f (new_AGEMA_signal_12107), .A1_t (new_AGEMA_signal_12108), .A1_f (new_AGEMA_signal_12109), .B0_t (SubBytesIns_Inst_Sbox_9_L9), .B0_f (new_AGEMA_signal_12656), .B1_t (new_AGEMA_signal_12657), .B1_f (new_AGEMA_signal_12658), .Z0_t (SubBytesIns_Inst_Sbox_9_L24), .Z0_f (new_AGEMA_signal_13277), .Z1_t (new_AGEMA_signal_13278), .Z1_f (new_AGEMA_signal_13279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L6), .A0_f (new_AGEMA_signal_12650), .A1_t (new_AGEMA_signal_12651), .A1_f (new_AGEMA_signal_12652), .B0_t (SubBytesIns_Inst_Sbox_9_L10), .B0_f (new_AGEMA_signal_12659), .B1_t (new_AGEMA_signal_12660), .B1_f (new_AGEMA_signal_12661), .Z0_t (SubBytesIns_Inst_Sbox_9_L25), .Z0_f (new_AGEMA_signal_13280), .Z1_t (new_AGEMA_signal_13281), .Z1_f (new_AGEMA_signal_13282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L7), .A0_f (new_AGEMA_signal_12653), .A1_t (new_AGEMA_signal_12654), .A1_f (new_AGEMA_signal_12655), .B0_t (SubBytesIns_Inst_Sbox_9_L9), .B0_f (new_AGEMA_signal_12656), .B1_t (new_AGEMA_signal_12657), .B1_f (new_AGEMA_signal_12658), .Z0_t (SubBytesIns_Inst_Sbox_9_L26), .Z0_f (new_AGEMA_signal_13283), .Z1_t (new_AGEMA_signal_13284), .Z1_f (new_AGEMA_signal_13285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L8), .A0_f (new_AGEMA_signal_11474), .A1_t (new_AGEMA_signal_11475), .A1_f (new_AGEMA_signal_11476), .B0_t (SubBytesIns_Inst_Sbox_9_L10), .B0_f (new_AGEMA_signal_12659), .B1_t (new_AGEMA_signal_12660), .B1_f (new_AGEMA_signal_12661), .Z0_t (SubBytesIns_Inst_Sbox_9_L27), .Z0_f (new_AGEMA_signal_13286), .Z1_t (new_AGEMA_signal_13287), .Z1_f (new_AGEMA_signal_13288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L11), .A0_f (new_AGEMA_signal_12662), .A1_t (new_AGEMA_signal_12663), .A1_f (new_AGEMA_signal_12664), .B0_t (SubBytesIns_Inst_Sbox_9_L14), .B0_f (new_AGEMA_signal_12104), .B1_t (new_AGEMA_signal_12105), .B1_f (new_AGEMA_signal_12106), .Z0_t (SubBytesIns_Inst_Sbox_9_L28), .Z0_f (new_AGEMA_signal_13289), .Z1_t (new_AGEMA_signal_13290), .Z1_f (new_AGEMA_signal_13291) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L11), .A0_f (new_AGEMA_signal_12662), .A1_t (new_AGEMA_signal_12663), .A1_f (new_AGEMA_signal_12664), .B0_t (SubBytesIns_Inst_Sbox_9_L17), .B0_f (new_AGEMA_signal_12110), .B1_t (new_AGEMA_signal_12111), .B1_f (new_AGEMA_signal_12112), .Z0_t (SubBytesIns_Inst_Sbox_9_L29), .Z0_f (new_AGEMA_signal_13292), .Z1_t (new_AGEMA_signal_13293), .Z1_f (new_AGEMA_signal_13294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L6), .A0_f (new_AGEMA_signal_12650), .A1_t (new_AGEMA_signal_12651), .A1_f (new_AGEMA_signal_12652), .B0_t (SubBytesIns_Inst_Sbox_9_L24), .B0_f (new_AGEMA_signal_13277), .B1_t (new_AGEMA_signal_13278), .B1_f (new_AGEMA_signal_13279), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .Z0_f (new_AGEMA_signal_13829), .Z1_t (new_AGEMA_signal_13830), .Z1_f (new_AGEMA_signal_13831) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L16), .A0_f (new_AGEMA_signal_13268), .A1_t (new_AGEMA_signal_13269), .A1_f (new_AGEMA_signal_13270), .B0_t (SubBytesIns_Inst_Sbox_9_L26), .B0_f (new_AGEMA_signal_13283), .B1_t (new_AGEMA_signal_13284), .B1_f (new_AGEMA_signal_13285), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .Z0_f (new_AGEMA_signal_13832), .Z1_t (new_AGEMA_signal_13833), .Z1_f (new_AGEMA_signal_13834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L19), .A0_f (new_AGEMA_signal_12665), .A1_t (new_AGEMA_signal_12666), .A1_f (new_AGEMA_signal_12667), .B0_t (SubBytesIns_Inst_Sbox_9_L28), .B0_f (new_AGEMA_signal_13289), .B1_t (new_AGEMA_signal_13290), .B1_f (new_AGEMA_signal_13291), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .Z0_f (new_AGEMA_signal_13835), .Z1_t (new_AGEMA_signal_13836), .Z1_f (new_AGEMA_signal_13837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L6), .A0_f (new_AGEMA_signal_12650), .A1_t (new_AGEMA_signal_12651), .A1_f (new_AGEMA_signal_12652), .B0_t (SubBytesIns_Inst_Sbox_9_L21), .B0_f (new_AGEMA_signal_13274), .B1_t (new_AGEMA_signal_13275), .B1_f (new_AGEMA_signal_13276), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .Z0_f (new_AGEMA_signal_13838), .Z1_t (new_AGEMA_signal_13839), .Z1_f (new_AGEMA_signal_13840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L20), .A0_f (new_AGEMA_signal_13271), .A1_t (new_AGEMA_signal_13272), .A1_f (new_AGEMA_signal_13273), .B0_t (SubBytesIns_Inst_Sbox_9_L22), .B0_f (new_AGEMA_signal_12668), .B1_t (new_AGEMA_signal_12669), .B1_f (new_AGEMA_signal_12670), .Z0_t (MixColumnsInput[11]), .Z0_f (new_AGEMA_signal_13841), .Z1_t (new_AGEMA_signal_13842), .Z1_f (new_AGEMA_signal_13843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L25), .A0_f (new_AGEMA_signal_13280), .A1_t (new_AGEMA_signal_13281), .A1_f (new_AGEMA_signal_13282), .B0_t (SubBytesIns_Inst_Sbox_9_L29), .B0_f (new_AGEMA_signal_13292), .B1_t (new_AGEMA_signal_13293), .B1_f (new_AGEMA_signal_13294), .Z0_t (MixColumnsInput[10]), .Z0_f (new_AGEMA_signal_13844), .Z1_t (new_AGEMA_signal_13845), .Z1_f (new_AGEMA_signal_13846) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L13), .A0_f (new_AGEMA_signal_13265), .A1_t (new_AGEMA_signal_13266), .A1_f (new_AGEMA_signal_13267), .B0_t (SubBytesIns_Inst_Sbox_9_L27), .B0_f (new_AGEMA_signal_13286), .B1_t (new_AGEMA_signal_13287), .B1_f (new_AGEMA_signal_13288), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .Z0_f (new_AGEMA_signal_13847), .Z1_t (new_AGEMA_signal_13848), .Z1_f (new_AGEMA_signal_13849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L6), .A0_f (new_AGEMA_signal_12650), .A1_t (new_AGEMA_signal_12651), .A1_f (new_AGEMA_signal_12652), .B0_t (SubBytesIns_Inst_Sbox_9_L23), .B0_f (new_AGEMA_signal_12671), .B1_t (new_AGEMA_signal_12672), .B1_f (new_AGEMA_signal_12673), .Z0_t (MixColumnsInput[8]), .Z0_f (new_AGEMA_signal_13295), .Z1_t (new_AGEMA_signal_13296), .Z1_f (new_AGEMA_signal_13297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[87]), .A0_f (ciphertext_s0_f[87]), .A1_t (ciphertext_s1_t[87]), .A1_f (ciphertext_s1_f[87]), .B0_t (ciphertext_s0_t[84]), .B0_f (ciphertext_s0_f[84]), .B1_t (ciphertext_s1_t[84]), .B1_f (ciphertext_s1_f[84]), .Z0_t (SubBytesIns_Inst_Sbox_10_T1), .Z0_f (new_AGEMA_signal_6646), .Z1_t (new_AGEMA_signal_6647), .Z1_f (new_AGEMA_signal_6648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[87]), .A0_f (ciphertext_s0_f[87]), .A1_t (ciphertext_s1_t[87]), .A1_f (ciphertext_s1_f[87]), .B0_t (ciphertext_s0_t[82]), .B0_f (ciphertext_s0_f[82]), .B1_t (ciphertext_s1_t[82]), .B1_f (ciphertext_s1_f[82]), .Z0_t (SubBytesIns_Inst_Sbox_10_T2), .Z0_f (new_AGEMA_signal_6649), .Z1_t (new_AGEMA_signal_6650), .Z1_f (new_AGEMA_signal_6651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[87]), .A0_f (ciphertext_s0_f[87]), .A1_t (ciphertext_s1_t[87]), .A1_f (ciphertext_s1_f[87]), .B0_t (ciphertext_s0_t[81]), .B0_f (ciphertext_s0_f[81]), .B1_t (ciphertext_s1_t[81]), .B1_f (ciphertext_s1_f[81]), .Z0_t (SubBytesIns_Inst_Sbox_10_T3), .Z0_f (new_AGEMA_signal_6652), .Z1_t (new_AGEMA_signal_6653), .Z1_f (new_AGEMA_signal_6654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[84]), .A0_f (ciphertext_s0_f[84]), .A1_t (ciphertext_s1_t[84]), .A1_f (ciphertext_s1_f[84]), .B0_t (ciphertext_s0_t[82]), .B0_f (ciphertext_s0_f[82]), .B1_t (ciphertext_s1_t[82]), .B1_f (ciphertext_s1_f[82]), .Z0_t (SubBytesIns_Inst_Sbox_10_T4), .Z0_f (new_AGEMA_signal_6655), .Z1_t (new_AGEMA_signal_6656), .Z1_f (new_AGEMA_signal_6657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[83]), .A0_f (ciphertext_s0_f[83]), .A1_t (ciphertext_s1_t[83]), .A1_f (ciphertext_s1_f[83]), .B0_t (ciphertext_s0_t[81]), .B0_f (ciphertext_s0_f[81]), .B1_t (ciphertext_s1_t[81]), .B1_f (ciphertext_s1_f[81]), .Z0_t (SubBytesIns_Inst_Sbox_10_T5), .Z0_f (new_AGEMA_signal_6658), .Z1_t (new_AGEMA_signal_6659), .Z1_f (new_AGEMA_signal_6660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T1), .A0_f (new_AGEMA_signal_6646), .A1_t (new_AGEMA_signal_6647), .A1_f (new_AGEMA_signal_6648), .B0_t (SubBytesIns_Inst_Sbox_10_T5), .B0_f (new_AGEMA_signal_6658), .B1_t (new_AGEMA_signal_6659), .B1_f (new_AGEMA_signal_6660), .Z0_t (SubBytesIns_Inst_Sbox_10_T6), .Z0_f (new_AGEMA_signal_7168), .Z1_t (new_AGEMA_signal_7169), .Z1_f (new_AGEMA_signal_7170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[86]), .A0_f (ciphertext_s0_f[86]), .A1_t (ciphertext_s1_t[86]), .A1_f (ciphertext_s1_f[86]), .B0_t (ciphertext_s0_t[85]), .B0_f (ciphertext_s0_f[85]), .B1_t (ciphertext_s1_t[85]), .B1_f (ciphertext_s1_f[85]), .Z0_t (SubBytesIns_Inst_Sbox_10_T7), .Z0_f (new_AGEMA_signal_6661), .Z1_t (new_AGEMA_signal_6662), .Z1_f (new_AGEMA_signal_6663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[80]), .A0_f (ciphertext_s0_f[80]), .A1_t (ciphertext_s1_t[80]), .A1_f (ciphertext_s1_f[80]), .B0_t (SubBytesIns_Inst_Sbox_10_T6), .B0_f (new_AGEMA_signal_7168), .B1_t (new_AGEMA_signal_7169), .B1_f (new_AGEMA_signal_7170), .Z0_t (SubBytesIns_Inst_Sbox_10_T8), .Z0_f (new_AGEMA_signal_7862), .Z1_t (new_AGEMA_signal_7863), .Z1_f (new_AGEMA_signal_7864) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[80]), .A0_f (ciphertext_s0_f[80]), .A1_t (ciphertext_s1_t[80]), .A1_f (ciphertext_s1_f[80]), .B0_t (SubBytesIns_Inst_Sbox_10_T7), .B0_f (new_AGEMA_signal_6661), .B1_t (new_AGEMA_signal_6662), .B1_f (new_AGEMA_signal_6663), .Z0_t (SubBytesIns_Inst_Sbox_10_T9), .Z0_f (new_AGEMA_signal_7171), .Z1_t (new_AGEMA_signal_7172), .Z1_f (new_AGEMA_signal_7173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T6), .A0_f (new_AGEMA_signal_7168), .A1_t (new_AGEMA_signal_7169), .A1_f (new_AGEMA_signal_7170), .B0_t (SubBytesIns_Inst_Sbox_10_T7), .B0_f (new_AGEMA_signal_6661), .B1_t (new_AGEMA_signal_6662), .B1_f (new_AGEMA_signal_6663), .Z0_t (SubBytesIns_Inst_Sbox_10_T10), .Z0_f (new_AGEMA_signal_7865), .Z1_t (new_AGEMA_signal_7866), .Z1_f (new_AGEMA_signal_7867) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[86]), .A0_f (ciphertext_s0_f[86]), .A1_t (ciphertext_s1_t[86]), .A1_f (ciphertext_s1_f[86]), .B0_t (ciphertext_s0_t[82]), .B0_f (ciphertext_s0_f[82]), .B1_t (ciphertext_s1_t[82]), .B1_f (ciphertext_s1_f[82]), .Z0_t (SubBytesIns_Inst_Sbox_10_T11), .Z0_f (new_AGEMA_signal_6664), .Z1_t (new_AGEMA_signal_6665), .Z1_f (new_AGEMA_signal_6666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[85]), .A0_f (ciphertext_s0_f[85]), .A1_t (ciphertext_s1_t[85]), .A1_f (ciphertext_s1_f[85]), .B0_t (ciphertext_s0_t[82]), .B0_f (ciphertext_s0_f[82]), .B1_t (ciphertext_s1_t[82]), .B1_f (ciphertext_s1_f[82]), .Z0_t (SubBytesIns_Inst_Sbox_10_T12), .Z0_f (new_AGEMA_signal_6667), .Z1_t (new_AGEMA_signal_6668), .Z1_f (new_AGEMA_signal_6669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T3), .A0_f (new_AGEMA_signal_6652), .A1_t (new_AGEMA_signal_6653), .A1_f (new_AGEMA_signal_6654), .B0_t (SubBytesIns_Inst_Sbox_10_T4), .B0_f (new_AGEMA_signal_6655), .B1_t (new_AGEMA_signal_6656), .B1_f (new_AGEMA_signal_6657), .Z0_t (SubBytesIns_Inst_Sbox_10_T13), .Z0_f (new_AGEMA_signal_7174), .Z1_t (new_AGEMA_signal_7175), .Z1_f (new_AGEMA_signal_7176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T6), .A0_f (new_AGEMA_signal_7168), .A1_t (new_AGEMA_signal_7169), .A1_f (new_AGEMA_signal_7170), .B0_t (SubBytesIns_Inst_Sbox_10_T11), .B0_f (new_AGEMA_signal_6664), .B1_t (new_AGEMA_signal_6665), .B1_f (new_AGEMA_signal_6666), .Z0_t (SubBytesIns_Inst_Sbox_10_T14), .Z0_f (new_AGEMA_signal_7868), .Z1_t (new_AGEMA_signal_7869), .Z1_f (new_AGEMA_signal_7870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T5), .A0_f (new_AGEMA_signal_6658), .A1_t (new_AGEMA_signal_6659), .A1_f (new_AGEMA_signal_6660), .B0_t (SubBytesIns_Inst_Sbox_10_T11), .B0_f (new_AGEMA_signal_6664), .B1_t (new_AGEMA_signal_6665), .B1_f (new_AGEMA_signal_6666), .Z0_t (SubBytesIns_Inst_Sbox_10_T15), .Z0_f (new_AGEMA_signal_7177), .Z1_t (new_AGEMA_signal_7178), .Z1_f (new_AGEMA_signal_7179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T5), .A0_f (new_AGEMA_signal_6658), .A1_t (new_AGEMA_signal_6659), .A1_f (new_AGEMA_signal_6660), .B0_t (SubBytesIns_Inst_Sbox_10_T12), .B0_f (new_AGEMA_signal_6667), .B1_t (new_AGEMA_signal_6668), .B1_f (new_AGEMA_signal_6669), .Z0_t (SubBytesIns_Inst_Sbox_10_T16), .Z0_f (new_AGEMA_signal_7180), .Z1_t (new_AGEMA_signal_7181), .Z1_f (new_AGEMA_signal_7182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T9), .A0_f (new_AGEMA_signal_7171), .A1_t (new_AGEMA_signal_7172), .A1_f (new_AGEMA_signal_7173), .B0_t (SubBytesIns_Inst_Sbox_10_T16), .B0_f (new_AGEMA_signal_7180), .B1_t (new_AGEMA_signal_7181), .B1_f (new_AGEMA_signal_7182), .Z0_t (SubBytesIns_Inst_Sbox_10_T17), .Z0_f (new_AGEMA_signal_7871), .Z1_t (new_AGEMA_signal_7872), .Z1_f (new_AGEMA_signal_7873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[84]), .A0_f (ciphertext_s0_f[84]), .A1_t (ciphertext_s1_t[84]), .A1_f (ciphertext_s1_f[84]), .B0_t (ciphertext_s0_t[80]), .B0_f (ciphertext_s0_f[80]), .B1_t (ciphertext_s1_t[80]), .B1_f (ciphertext_s1_f[80]), .Z0_t (SubBytesIns_Inst_Sbox_10_T18), .Z0_f (new_AGEMA_signal_6670), .Z1_t (new_AGEMA_signal_6671), .Z1_f (new_AGEMA_signal_6672) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T7), .A0_f (new_AGEMA_signal_6661), .A1_t (new_AGEMA_signal_6662), .A1_f (new_AGEMA_signal_6663), .B0_t (SubBytesIns_Inst_Sbox_10_T18), .B0_f (new_AGEMA_signal_6670), .B1_t (new_AGEMA_signal_6671), .B1_f (new_AGEMA_signal_6672), .Z0_t (SubBytesIns_Inst_Sbox_10_T19), .Z0_f (new_AGEMA_signal_7183), .Z1_t (new_AGEMA_signal_7184), .Z1_f (new_AGEMA_signal_7185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T1), .A0_f (new_AGEMA_signal_6646), .A1_t (new_AGEMA_signal_6647), .A1_f (new_AGEMA_signal_6648), .B0_t (SubBytesIns_Inst_Sbox_10_T19), .B0_f (new_AGEMA_signal_7183), .B1_t (new_AGEMA_signal_7184), .B1_f (new_AGEMA_signal_7185), .Z0_t (SubBytesIns_Inst_Sbox_10_T20), .Z0_f (new_AGEMA_signal_7874), .Z1_t (new_AGEMA_signal_7875), .Z1_f (new_AGEMA_signal_7876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[81]), .A0_f (ciphertext_s0_f[81]), .A1_t (ciphertext_s1_t[81]), .A1_f (ciphertext_s1_f[81]), .B0_t (ciphertext_s0_t[80]), .B0_f (ciphertext_s0_f[80]), .B1_t (ciphertext_s1_t[80]), .B1_f (ciphertext_s1_f[80]), .Z0_t (SubBytesIns_Inst_Sbox_10_T21), .Z0_f (new_AGEMA_signal_6673), .Z1_t (new_AGEMA_signal_6674), .Z1_f (new_AGEMA_signal_6675) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T7), .A0_f (new_AGEMA_signal_6661), .A1_t (new_AGEMA_signal_6662), .A1_f (new_AGEMA_signal_6663), .B0_t (SubBytesIns_Inst_Sbox_10_T21), .B0_f (new_AGEMA_signal_6673), .B1_t (new_AGEMA_signal_6674), .B1_f (new_AGEMA_signal_6675), .Z0_t (SubBytesIns_Inst_Sbox_10_T22), .Z0_f (new_AGEMA_signal_7186), .Z1_t (new_AGEMA_signal_7187), .Z1_f (new_AGEMA_signal_7188) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T2), .A0_f (new_AGEMA_signal_6649), .A1_t (new_AGEMA_signal_6650), .A1_f (new_AGEMA_signal_6651), .B0_t (SubBytesIns_Inst_Sbox_10_T22), .B0_f (new_AGEMA_signal_7186), .B1_t (new_AGEMA_signal_7187), .B1_f (new_AGEMA_signal_7188), .Z0_t (SubBytesIns_Inst_Sbox_10_T23), .Z0_f (new_AGEMA_signal_7877), .Z1_t (new_AGEMA_signal_7878), .Z1_f (new_AGEMA_signal_7879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T2), .A0_f (new_AGEMA_signal_6649), .A1_t (new_AGEMA_signal_6650), .A1_f (new_AGEMA_signal_6651), .B0_t (SubBytesIns_Inst_Sbox_10_T10), .B0_f (new_AGEMA_signal_7865), .B1_t (new_AGEMA_signal_7866), .B1_f (new_AGEMA_signal_7867), .Z0_t (SubBytesIns_Inst_Sbox_10_T24), .Z0_f (new_AGEMA_signal_8474), .Z1_t (new_AGEMA_signal_8475), .Z1_f (new_AGEMA_signal_8476) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T20), .A0_f (new_AGEMA_signal_7874), .A1_t (new_AGEMA_signal_7875), .A1_f (new_AGEMA_signal_7876), .B0_t (SubBytesIns_Inst_Sbox_10_T17), .B0_f (new_AGEMA_signal_7871), .B1_t (new_AGEMA_signal_7872), .B1_f (new_AGEMA_signal_7873), .Z0_t (SubBytesIns_Inst_Sbox_10_T25), .Z0_f (new_AGEMA_signal_8477), .Z1_t (new_AGEMA_signal_8478), .Z1_f (new_AGEMA_signal_8479) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T3), .A0_f (new_AGEMA_signal_6652), .A1_t (new_AGEMA_signal_6653), .A1_f (new_AGEMA_signal_6654), .B0_t (SubBytesIns_Inst_Sbox_10_T16), .B0_f (new_AGEMA_signal_7180), .B1_t (new_AGEMA_signal_7181), .B1_f (new_AGEMA_signal_7182), .Z0_t (SubBytesIns_Inst_Sbox_10_T26), .Z0_f (new_AGEMA_signal_7880), .Z1_t (new_AGEMA_signal_7881), .Z1_f (new_AGEMA_signal_7882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T1), .A0_f (new_AGEMA_signal_6646), .A1_t (new_AGEMA_signal_6647), .A1_f (new_AGEMA_signal_6648), .B0_t (SubBytesIns_Inst_Sbox_10_T12), .B0_f (new_AGEMA_signal_6667), .B1_t (new_AGEMA_signal_6668), .B1_f (new_AGEMA_signal_6669), .Z0_t (SubBytesIns_Inst_Sbox_10_T27), .Z0_f (new_AGEMA_signal_7189), .Z1_t (new_AGEMA_signal_7190), .Z1_f (new_AGEMA_signal_7191) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T13), .A0_f (new_AGEMA_signal_7174), .A1_t (new_AGEMA_signal_7175), .A1_f (new_AGEMA_signal_7176), .B0_t (SubBytesIns_Inst_Sbox_10_T6), .B0_f (new_AGEMA_signal_7168), .B1_t (new_AGEMA_signal_7169), .B1_f (new_AGEMA_signal_7170), .Z0_t (SubBytesIns_Inst_Sbox_10_M1), .Z0_f (new_AGEMA_signal_7883), .Z1_t (new_AGEMA_signal_7884), .Z1_f (new_AGEMA_signal_7885) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T23), .A0_f (new_AGEMA_signal_7877), .A1_t (new_AGEMA_signal_7878), .A1_f (new_AGEMA_signal_7879), .B0_t (SubBytesIns_Inst_Sbox_10_T8), .B0_f (new_AGEMA_signal_7862), .B1_t (new_AGEMA_signal_7863), .B1_f (new_AGEMA_signal_7864), .Z0_t (SubBytesIns_Inst_Sbox_10_M2), .Z0_f (new_AGEMA_signal_8480), .Z1_t (new_AGEMA_signal_8481), .Z1_f (new_AGEMA_signal_8482) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T14), .A0_f (new_AGEMA_signal_7868), .A1_t (new_AGEMA_signal_7869), .A1_f (new_AGEMA_signal_7870), .B0_t (SubBytesIns_Inst_Sbox_10_M1), .B0_f (new_AGEMA_signal_7883), .B1_t (new_AGEMA_signal_7884), .B1_f (new_AGEMA_signal_7885), .Z0_t (SubBytesIns_Inst_Sbox_10_M3), .Z0_f (new_AGEMA_signal_8483), .Z1_t (new_AGEMA_signal_8484), .Z1_f (new_AGEMA_signal_8485) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T19), .A0_f (new_AGEMA_signal_7183), .A1_t (new_AGEMA_signal_7184), .A1_f (new_AGEMA_signal_7185), .B0_t (ciphertext_s0_t[80]), .B0_f (ciphertext_s0_f[80]), .B1_t (ciphertext_s1_t[80]), .B1_f (ciphertext_s1_f[80]), .Z0_t (SubBytesIns_Inst_Sbox_10_M4), .Z0_f (new_AGEMA_signal_7886), .Z1_t (new_AGEMA_signal_7887), .Z1_f (new_AGEMA_signal_7888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M4), .A0_f (new_AGEMA_signal_7886), .A1_t (new_AGEMA_signal_7887), .A1_f (new_AGEMA_signal_7888), .B0_t (SubBytesIns_Inst_Sbox_10_M1), .B0_f (new_AGEMA_signal_7883), .B1_t (new_AGEMA_signal_7884), .B1_f (new_AGEMA_signal_7885), .Z0_t (SubBytesIns_Inst_Sbox_10_M5), .Z0_f (new_AGEMA_signal_8486), .Z1_t (new_AGEMA_signal_8487), .Z1_f (new_AGEMA_signal_8488) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T3), .A0_f (new_AGEMA_signal_6652), .A1_t (new_AGEMA_signal_6653), .A1_f (new_AGEMA_signal_6654), .B0_t (SubBytesIns_Inst_Sbox_10_T16), .B0_f (new_AGEMA_signal_7180), .B1_t (new_AGEMA_signal_7181), .B1_f (new_AGEMA_signal_7182), .Z0_t (SubBytesIns_Inst_Sbox_10_M6), .Z0_f (new_AGEMA_signal_7889), .Z1_t (new_AGEMA_signal_7890), .Z1_f (new_AGEMA_signal_7891) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T22), .A0_f (new_AGEMA_signal_7186), .A1_t (new_AGEMA_signal_7187), .A1_f (new_AGEMA_signal_7188), .B0_t (SubBytesIns_Inst_Sbox_10_T9), .B0_f (new_AGEMA_signal_7171), .B1_t (new_AGEMA_signal_7172), .B1_f (new_AGEMA_signal_7173), .Z0_t (SubBytesIns_Inst_Sbox_10_M7), .Z0_f (new_AGEMA_signal_7892), .Z1_t (new_AGEMA_signal_7893), .Z1_f (new_AGEMA_signal_7894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T26), .A0_f (new_AGEMA_signal_7880), .A1_t (new_AGEMA_signal_7881), .A1_f (new_AGEMA_signal_7882), .B0_t (SubBytesIns_Inst_Sbox_10_M6), .B0_f (new_AGEMA_signal_7889), .B1_t (new_AGEMA_signal_7890), .B1_f (new_AGEMA_signal_7891), .Z0_t (SubBytesIns_Inst_Sbox_10_M8), .Z0_f (new_AGEMA_signal_8489), .Z1_t (new_AGEMA_signal_8490), .Z1_f (new_AGEMA_signal_8491) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T20), .A0_f (new_AGEMA_signal_7874), .A1_t (new_AGEMA_signal_7875), .A1_f (new_AGEMA_signal_7876), .B0_t (SubBytesIns_Inst_Sbox_10_T17), .B0_f (new_AGEMA_signal_7871), .B1_t (new_AGEMA_signal_7872), .B1_f (new_AGEMA_signal_7873), .Z0_t (SubBytesIns_Inst_Sbox_10_M9), .Z0_f (new_AGEMA_signal_8492), .Z1_t (new_AGEMA_signal_8493), .Z1_f (new_AGEMA_signal_8494) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M9), .A0_f (new_AGEMA_signal_8492), .A1_t (new_AGEMA_signal_8493), .A1_f (new_AGEMA_signal_8494), .B0_t (SubBytesIns_Inst_Sbox_10_M6), .B0_f (new_AGEMA_signal_7889), .B1_t (new_AGEMA_signal_7890), .B1_f (new_AGEMA_signal_7891), .Z0_t (SubBytesIns_Inst_Sbox_10_M10), .Z0_f (new_AGEMA_signal_8846), .Z1_t (new_AGEMA_signal_8847), .Z1_f (new_AGEMA_signal_8848) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T1), .A0_f (new_AGEMA_signal_6646), .A1_t (new_AGEMA_signal_6647), .A1_f (new_AGEMA_signal_6648), .B0_t (SubBytesIns_Inst_Sbox_10_T15), .B0_f (new_AGEMA_signal_7177), .B1_t (new_AGEMA_signal_7178), .B1_f (new_AGEMA_signal_7179), .Z0_t (SubBytesIns_Inst_Sbox_10_M11), .Z0_f (new_AGEMA_signal_7895), .Z1_t (new_AGEMA_signal_7896), .Z1_f (new_AGEMA_signal_7897) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T4), .A0_f (new_AGEMA_signal_6655), .A1_t (new_AGEMA_signal_6656), .A1_f (new_AGEMA_signal_6657), .B0_t (SubBytesIns_Inst_Sbox_10_T27), .B0_f (new_AGEMA_signal_7189), .B1_t (new_AGEMA_signal_7190), .B1_f (new_AGEMA_signal_7191), .Z0_t (SubBytesIns_Inst_Sbox_10_M12), .Z0_f (new_AGEMA_signal_7898), .Z1_t (new_AGEMA_signal_7899), .Z1_f (new_AGEMA_signal_7900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M12), .A0_f (new_AGEMA_signal_7898), .A1_t (new_AGEMA_signal_7899), .A1_f (new_AGEMA_signal_7900), .B0_t (SubBytesIns_Inst_Sbox_10_M11), .B0_f (new_AGEMA_signal_7895), .B1_t (new_AGEMA_signal_7896), .B1_f (new_AGEMA_signal_7897), .Z0_t (SubBytesIns_Inst_Sbox_10_M13), .Z0_f (new_AGEMA_signal_8495), .Z1_t (new_AGEMA_signal_8496), .Z1_f (new_AGEMA_signal_8497) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T2), .A0_f (new_AGEMA_signal_6649), .A1_t (new_AGEMA_signal_6650), .A1_f (new_AGEMA_signal_6651), .B0_t (SubBytesIns_Inst_Sbox_10_T10), .B0_f (new_AGEMA_signal_7865), .B1_t (new_AGEMA_signal_7866), .B1_f (new_AGEMA_signal_7867), .Z0_t (SubBytesIns_Inst_Sbox_10_M14), .Z0_f (new_AGEMA_signal_8498), .Z1_t (new_AGEMA_signal_8499), .Z1_f (new_AGEMA_signal_8500) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M14), .A0_f (new_AGEMA_signal_8498), .A1_t (new_AGEMA_signal_8499), .A1_f (new_AGEMA_signal_8500), .B0_t (SubBytesIns_Inst_Sbox_10_M11), .B0_f (new_AGEMA_signal_7895), .B1_t (new_AGEMA_signal_7896), .B1_f (new_AGEMA_signal_7897), .Z0_t (SubBytesIns_Inst_Sbox_10_M15), .Z0_f (new_AGEMA_signal_8849), .Z1_t (new_AGEMA_signal_8850), .Z1_f (new_AGEMA_signal_8851) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M3), .A0_f (new_AGEMA_signal_8483), .A1_t (new_AGEMA_signal_8484), .A1_f (new_AGEMA_signal_8485), .B0_t (SubBytesIns_Inst_Sbox_10_M2), .B0_f (new_AGEMA_signal_8480), .B1_t (new_AGEMA_signal_8481), .B1_f (new_AGEMA_signal_8482), .Z0_t (SubBytesIns_Inst_Sbox_10_M16), .Z0_f (new_AGEMA_signal_8852), .Z1_t (new_AGEMA_signal_8853), .Z1_f (new_AGEMA_signal_8854) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M5), .A0_f (new_AGEMA_signal_8486), .A1_t (new_AGEMA_signal_8487), .A1_f (new_AGEMA_signal_8488), .B0_t (SubBytesIns_Inst_Sbox_10_T24), .B0_f (new_AGEMA_signal_8474), .B1_t (new_AGEMA_signal_8475), .B1_f (new_AGEMA_signal_8476), .Z0_t (SubBytesIns_Inst_Sbox_10_M17), .Z0_f (new_AGEMA_signal_8855), .Z1_t (new_AGEMA_signal_8856), .Z1_f (new_AGEMA_signal_8857) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M8), .A0_f (new_AGEMA_signal_8489), .A1_t (new_AGEMA_signal_8490), .A1_f (new_AGEMA_signal_8491), .B0_t (SubBytesIns_Inst_Sbox_10_M7), .B0_f (new_AGEMA_signal_7892), .B1_t (new_AGEMA_signal_7893), .B1_f (new_AGEMA_signal_7894), .Z0_t (SubBytesIns_Inst_Sbox_10_M18), .Z0_f (new_AGEMA_signal_8858), .Z1_t (new_AGEMA_signal_8859), .Z1_f (new_AGEMA_signal_8860) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M10), .A0_f (new_AGEMA_signal_8846), .A1_t (new_AGEMA_signal_8847), .A1_f (new_AGEMA_signal_8848), .B0_t (SubBytesIns_Inst_Sbox_10_M15), .B0_f (new_AGEMA_signal_8849), .B1_t (new_AGEMA_signal_8850), .B1_f (new_AGEMA_signal_8851), .Z0_t (SubBytesIns_Inst_Sbox_10_M19), .Z0_f (new_AGEMA_signal_9104), .Z1_t (new_AGEMA_signal_9105), .Z1_f (new_AGEMA_signal_9106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M16), .A0_f (new_AGEMA_signal_8852), .A1_t (new_AGEMA_signal_8853), .A1_f (new_AGEMA_signal_8854), .B0_t (SubBytesIns_Inst_Sbox_10_M13), .B0_f (new_AGEMA_signal_8495), .B1_t (new_AGEMA_signal_8496), .B1_f (new_AGEMA_signal_8497), .Z0_t (SubBytesIns_Inst_Sbox_10_M20), .Z0_f (new_AGEMA_signal_9107), .Z1_t (new_AGEMA_signal_9108), .Z1_f (new_AGEMA_signal_9109) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M17), .A0_f (new_AGEMA_signal_8855), .A1_t (new_AGEMA_signal_8856), .A1_f (new_AGEMA_signal_8857), .B0_t (SubBytesIns_Inst_Sbox_10_M15), .B0_f (new_AGEMA_signal_8849), .B1_t (new_AGEMA_signal_8850), .B1_f (new_AGEMA_signal_8851), .Z0_t (SubBytesIns_Inst_Sbox_10_M21), .Z0_f (new_AGEMA_signal_9110), .Z1_t (new_AGEMA_signal_9111), .Z1_f (new_AGEMA_signal_9112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M18), .A0_f (new_AGEMA_signal_8858), .A1_t (new_AGEMA_signal_8859), .A1_f (new_AGEMA_signal_8860), .B0_t (SubBytesIns_Inst_Sbox_10_M13), .B0_f (new_AGEMA_signal_8495), .B1_t (new_AGEMA_signal_8496), .B1_f (new_AGEMA_signal_8497), .Z0_t (SubBytesIns_Inst_Sbox_10_M22), .Z0_f (new_AGEMA_signal_9113), .Z1_t (new_AGEMA_signal_9114), .Z1_f (new_AGEMA_signal_9115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M19), .A0_f (new_AGEMA_signal_9104), .A1_t (new_AGEMA_signal_9105), .A1_f (new_AGEMA_signal_9106), .B0_t (SubBytesIns_Inst_Sbox_10_T25), .B0_f (new_AGEMA_signal_8477), .B1_t (new_AGEMA_signal_8478), .B1_f (new_AGEMA_signal_8479), .Z0_t (SubBytesIns_Inst_Sbox_10_M23), .Z0_f (new_AGEMA_signal_9344), .Z1_t (new_AGEMA_signal_9345), .Z1_f (new_AGEMA_signal_9346) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M22), .A0_f (new_AGEMA_signal_9113), .A1_t (new_AGEMA_signal_9114), .A1_f (new_AGEMA_signal_9115), .B0_t (SubBytesIns_Inst_Sbox_10_M23), .B0_f (new_AGEMA_signal_9344), .B1_t (new_AGEMA_signal_9345), .B1_f (new_AGEMA_signal_9346), .Z0_t (SubBytesIns_Inst_Sbox_10_M24), .Z0_f (new_AGEMA_signal_9626), .Z1_t (new_AGEMA_signal_9627), .Z1_f (new_AGEMA_signal_9628) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M22), .A0_f (new_AGEMA_signal_9113), .A1_t (new_AGEMA_signal_9114), .A1_f (new_AGEMA_signal_9115), .B0_t (SubBytesIns_Inst_Sbox_10_M20), .B0_f (new_AGEMA_signal_9107), .B1_t (new_AGEMA_signal_9108), .B1_f (new_AGEMA_signal_9109), .Z0_t (SubBytesIns_Inst_Sbox_10_M25), .Z0_f (new_AGEMA_signal_9347), .Z1_t (new_AGEMA_signal_9348), .Z1_f (new_AGEMA_signal_9349) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M21), .A0_f (new_AGEMA_signal_9110), .A1_t (new_AGEMA_signal_9111), .A1_f (new_AGEMA_signal_9112), .B0_t (SubBytesIns_Inst_Sbox_10_M25), .B0_f (new_AGEMA_signal_9347), .B1_t (new_AGEMA_signal_9348), .B1_f (new_AGEMA_signal_9349), .Z0_t (SubBytesIns_Inst_Sbox_10_M26), .Z0_f (new_AGEMA_signal_9629), .Z1_t (new_AGEMA_signal_9630), .Z1_f (new_AGEMA_signal_9631) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M20), .A0_f (new_AGEMA_signal_9107), .A1_t (new_AGEMA_signal_9108), .A1_f (new_AGEMA_signal_9109), .B0_t (SubBytesIns_Inst_Sbox_10_M21), .B0_f (new_AGEMA_signal_9110), .B1_t (new_AGEMA_signal_9111), .B1_f (new_AGEMA_signal_9112), .Z0_t (SubBytesIns_Inst_Sbox_10_M27), .Z0_f (new_AGEMA_signal_9350), .Z1_t (new_AGEMA_signal_9351), .Z1_f (new_AGEMA_signal_9352) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M23), .A0_f (new_AGEMA_signal_9344), .A1_t (new_AGEMA_signal_9345), .A1_f (new_AGEMA_signal_9346), .B0_t (SubBytesIns_Inst_Sbox_10_M25), .B0_f (new_AGEMA_signal_9347), .B1_t (new_AGEMA_signal_9348), .B1_f (new_AGEMA_signal_9349), .Z0_t (SubBytesIns_Inst_Sbox_10_M28), .Z0_f (new_AGEMA_signal_9632), .Z1_t (new_AGEMA_signal_9633), .Z1_f (new_AGEMA_signal_9634) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M28), .A0_f (new_AGEMA_signal_9632), .A1_t (new_AGEMA_signal_9633), .A1_f (new_AGEMA_signal_9634), .B0_t (SubBytesIns_Inst_Sbox_10_M27), .B0_f (new_AGEMA_signal_9350), .B1_t (new_AGEMA_signal_9351), .B1_f (new_AGEMA_signal_9352), .Z0_t (SubBytesIns_Inst_Sbox_10_M29), .Z0_f (new_AGEMA_signal_9926), .Z1_t (new_AGEMA_signal_9927), .Z1_f (new_AGEMA_signal_9928) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M26), .A0_f (new_AGEMA_signal_9629), .A1_t (new_AGEMA_signal_9630), .A1_f (new_AGEMA_signal_9631), .B0_t (SubBytesIns_Inst_Sbox_10_M24), .B0_f (new_AGEMA_signal_9626), .B1_t (new_AGEMA_signal_9627), .B1_f (new_AGEMA_signal_9628), .Z0_t (SubBytesIns_Inst_Sbox_10_M30), .Z0_f (new_AGEMA_signal_9929), .Z1_t (new_AGEMA_signal_9930), .Z1_f (new_AGEMA_signal_9931) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M20), .A0_f (new_AGEMA_signal_9107), .A1_t (new_AGEMA_signal_9108), .A1_f (new_AGEMA_signal_9109), .B0_t (SubBytesIns_Inst_Sbox_10_M23), .B0_f (new_AGEMA_signal_9344), .B1_t (new_AGEMA_signal_9345), .B1_f (new_AGEMA_signal_9346), .Z0_t (SubBytesIns_Inst_Sbox_10_M31), .Z0_f (new_AGEMA_signal_9635), .Z1_t (new_AGEMA_signal_9636), .Z1_f (new_AGEMA_signal_9637) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M27), .A0_f (new_AGEMA_signal_9350), .A1_t (new_AGEMA_signal_9351), .A1_f (new_AGEMA_signal_9352), .B0_t (SubBytesIns_Inst_Sbox_10_M31), .B0_f (new_AGEMA_signal_9635), .B1_t (new_AGEMA_signal_9636), .B1_f (new_AGEMA_signal_9637), .Z0_t (SubBytesIns_Inst_Sbox_10_M32), .Z0_f (new_AGEMA_signal_9932), .Z1_t (new_AGEMA_signal_9933), .Z1_f (new_AGEMA_signal_9934) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M27), .A0_f (new_AGEMA_signal_9350), .A1_t (new_AGEMA_signal_9351), .A1_f (new_AGEMA_signal_9352), .B0_t (SubBytesIns_Inst_Sbox_10_M25), .B0_f (new_AGEMA_signal_9347), .B1_t (new_AGEMA_signal_9348), .B1_f (new_AGEMA_signal_9349), .Z0_t (SubBytesIns_Inst_Sbox_10_M33), .Z0_f (new_AGEMA_signal_9638), .Z1_t (new_AGEMA_signal_9639), .Z1_f (new_AGEMA_signal_9640) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M21), .A0_f (new_AGEMA_signal_9110), .A1_t (new_AGEMA_signal_9111), .A1_f (new_AGEMA_signal_9112), .B0_t (SubBytesIns_Inst_Sbox_10_M22), .B0_f (new_AGEMA_signal_9113), .B1_t (new_AGEMA_signal_9114), .B1_f (new_AGEMA_signal_9115), .Z0_t (SubBytesIns_Inst_Sbox_10_M34), .Z0_f (new_AGEMA_signal_9353), .Z1_t (new_AGEMA_signal_9354), .Z1_f (new_AGEMA_signal_9355) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M24), .A0_f (new_AGEMA_signal_9626), .A1_t (new_AGEMA_signal_9627), .A1_f (new_AGEMA_signal_9628), .B0_t (SubBytesIns_Inst_Sbox_10_M34), .B0_f (new_AGEMA_signal_9353), .B1_t (new_AGEMA_signal_9354), .B1_f (new_AGEMA_signal_9355), .Z0_t (SubBytesIns_Inst_Sbox_10_M35), .Z0_f (new_AGEMA_signal_9935), .Z1_t (new_AGEMA_signal_9936), .Z1_f (new_AGEMA_signal_9937) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M24), .A0_f (new_AGEMA_signal_9626), .A1_t (new_AGEMA_signal_9627), .A1_f (new_AGEMA_signal_9628), .B0_t (SubBytesIns_Inst_Sbox_10_M25), .B0_f (new_AGEMA_signal_9347), .B1_t (new_AGEMA_signal_9348), .B1_f (new_AGEMA_signal_9349), .Z0_t (SubBytesIns_Inst_Sbox_10_M36), .Z0_f (new_AGEMA_signal_9938), .Z1_t (new_AGEMA_signal_9939), .Z1_f (new_AGEMA_signal_9940) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M21), .A0_f (new_AGEMA_signal_9110), .A1_t (new_AGEMA_signal_9111), .A1_f (new_AGEMA_signal_9112), .B0_t (SubBytesIns_Inst_Sbox_10_M29), .B0_f (new_AGEMA_signal_9926), .B1_t (new_AGEMA_signal_9927), .B1_f (new_AGEMA_signal_9928), .Z0_t (SubBytesIns_Inst_Sbox_10_M37), .Z0_f (new_AGEMA_signal_10184), .Z1_t (new_AGEMA_signal_10185), .Z1_f (new_AGEMA_signal_10186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M32), .A0_f (new_AGEMA_signal_9932), .A1_t (new_AGEMA_signal_9933), .A1_f (new_AGEMA_signal_9934), .B0_t (SubBytesIns_Inst_Sbox_10_M33), .B0_f (new_AGEMA_signal_9638), .B1_t (new_AGEMA_signal_9639), .B1_f (new_AGEMA_signal_9640), .Z0_t (SubBytesIns_Inst_Sbox_10_M38), .Z0_f (new_AGEMA_signal_10187), .Z1_t (new_AGEMA_signal_10188), .Z1_f (new_AGEMA_signal_10189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M23), .A0_f (new_AGEMA_signal_9344), .A1_t (new_AGEMA_signal_9345), .A1_f (new_AGEMA_signal_9346), .B0_t (SubBytesIns_Inst_Sbox_10_M30), .B0_f (new_AGEMA_signal_9929), .B1_t (new_AGEMA_signal_9930), .B1_f (new_AGEMA_signal_9931), .Z0_t (SubBytesIns_Inst_Sbox_10_M39), .Z0_f (new_AGEMA_signal_10190), .Z1_t (new_AGEMA_signal_10191), .Z1_f (new_AGEMA_signal_10192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M35), .A0_f (new_AGEMA_signal_9935), .A1_t (new_AGEMA_signal_9936), .A1_f (new_AGEMA_signal_9937), .B0_t (SubBytesIns_Inst_Sbox_10_M36), .B0_f (new_AGEMA_signal_9938), .B1_t (new_AGEMA_signal_9939), .B1_f (new_AGEMA_signal_9940), .Z0_t (SubBytesIns_Inst_Sbox_10_M40), .Z0_f (new_AGEMA_signal_10193), .Z1_t (new_AGEMA_signal_10194), .Z1_f (new_AGEMA_signal_10195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M38), .A0_f (new_AGEMA_signal_10187), .A1_t (new_AGEMA_signal_10188), .A1_f (new_AGEMA_signal_10189), .B0_t (SubBytesIns_Inst_Sbox_10_M40), .B0_f (new_AGEMA_signal_10193), .B1_t (new_AGEMA_signal_10194), .B1_f (new_AGEMA_signal_10195), .Z0_t (SubBytesIns_Inst_Sbox_10_M41), .Z0_f (new_AGEMA_signal_10760), .Z1_t (new_AGEMA_signal_10761), .Z1_f (new_AGEMA_signal_10762) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M37), .A0_f (new_AGEMA_signal_10184), .A1_t (new_AGEMA_signal_10185), .A1_f (new_AGEMA_signal_10186), .B0_t (SubBytesIns_Inst_Sbox_10_M39), .B0_f (new_AGEMA_signal_10190), .B1_t (new_AGEMA_signal_10191), .B1_f (new_AGEMA_signal_10192), .Z0_t (SubBytesIns_Inst_Sbox_10_M42), .Z0_f (new_AGEMA_signal_10763), .Z1_t (new_AGEMA_signal_10764), .Z1_f (new_AGEMA_signal_10765) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M37), .A0_f (new_AGEMA_signal_10184), .A1_t (new_AGEMA_signal_10185), .A1_f (new_AGEMA_signal_10186), .B0_t (SubBytesIns_Inst_Sbox_10_M38), .B0_f (new_AGEMA_signal_10187), .B1_t (new_AGEMA_signal_10188), .B1_f (new_AGEMA_signal_10189), .Z0_t (SubBytesIns_Inst_Sbox_10_M43), .Z0_f (new_AGEMA_signal_10766), .Z1_t (new_AGEMA_signal_10767), .Z1_f (new_AGEMA_signal_10768) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M39), .A0_f (new_AGEMA_signal_10190), .A1_t (new_AGEMA_signal_10191), .A1_f (new_AGEMA_signal_10192), .B0_t (SubBytesIns_Inst_Sbox_10_M40), .B0_f (new_AGEMA_signal_10193), .B1_t (new_AGEMA_signal_10194), .B1_f (new_AGEMA_signal_10195), .Z0_t (SubBytesIns_Inst_Sbox_10_M44), .Z0_f (new_AGEMA_signal_10769), .Z1_t (new_AGEMA_signal_10770), .Z1_f (new_AGEMA_signal_10771) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M42), .A0_f (new_AGEMA_signal_10763), .A1_t (new_AGEMA_signal_10764), .A1_f (new_AGEMA_signal_10765), .B0_t (SubBytesIns_Inst_Sbox_10_M41), .B0_f (new_AGEMA_signal_10760), .B1_t (new_AGEMA_signal_10761), .B1_f (new_AGEMA_signal_10762), .Z0_t (SubBytesIns_Inst_Sbox_10_M45), .Z0_f (new_AGEMA_signal_11480), .Z1_t (new_AGEMA_signal_11481), .Z1_f (new_AGEMA_signal_11482) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M44), .A0_f (new_AGEMA_signal_10769), .A1_t (new_AGEMA_signal_10770), .A1_f (new_AGEMA_signal_10771), .B0_t (SubBytesIns_Inst_Sbox_10_T6), .B0_f (new_AGEMA_signal_7168), .B1_t (new_AGEMA_signal_7169), .B1_f (new_AGEMA_signal_7170), .Z0_t (SubBytesIns_Inst_Sbox_10_M46), .Z0_f (new_AGEMA_signal_11483), .Z1_t (new_AGEMA_signal_11484), .Z1_f (new_AGEMA_signal_11485) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M40), .A0_f (new_AGEMA_signal_10193), .A1_t (new_AGEMA_signal_10194), .A1_f (new_AGEMA_signal_10195), .B0_t (SubBytesIns_Inst_Sbox_10_T8), .B0_f (new_AGEMA_signal_7862), .B1_t (new_AGEMA_signal_7863), .B1_f (new_AGEMA_signal_7864), .Z0_t (SubBytesIns_Inst_Sbox_10_M47), .Z0_f (new_AGEMA_signal_10772), .Z1_t (new_AGEMA_signal_10773), .Z1_f (new_AGEMA_signal_10774) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M39), .A0_f (new_AGEMA_signal_10190), .A1_t (new_AGEMA_signal_10191), .A1_f (new_AGEMA_signal_10192), .B0_t (ciphertext_s0_t[80]), .B0_f (ciphertext_s0_f[80]), .B1_t (ciphertext_s1_t[80]), .B1_f (ciphertext_s1_f[80]), .Z0_t (SubBytesIns_Inst_Sbox_10_M48), .Z0_f (new_AGEMA_signal_10775), .Z1_t (new_AGEMA_signal_10776), .Z1_f (new_AGEMA_signal_10777) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M43), .A0_f (new_AGEMA_signal_10766), .A1_t (new_AGEMA_signal_10767), .A1_f (new_AGEMA_signal_10768), .B0_t (SubBytesIns_Inst_Sbox_10_T16), .B0_f (new_AGEMA_signal_7180), .B1_t (new_AGEMA_signal_7181), .B1_f (new_AGEMA_signal_7182), .Z0_t (SubBytesIns_Inst_Sbox_10_M49), .Z0_f (new_AGEMA_signal_11486), .Z1_t (new_AGEMA_signal_11487), .Z1_f (new_AGEMA_signal_11488) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M38), .A0_f (new_AGEMA_signal_10187), .A1_t (new_AGEMA_signal_10188), .A1_f (new_AGEMA_signal_10189), .B0_t (SubBytesIns_Inst_Sbox_10_T9), .B0_f (new_AGEMA_signal_7171), .B1_t (new_AGEMA_signal_7172), .B1_f (new_AGEMA_signal_7173), .Z0_t (SubBytesIns_Inst_Sbox_10_M50), .Z0_f (new_AGEMA_signal_10778), .Z1_t (new_AGEMA_signal_10779), .Z1_f (new_AGEMA_signal_10780) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M37), .A0_f (new_AGEMA_signal_10184), .A1_t (new_AGEMA_signal_10185), .A1_f (new_AGEMA_signal_10186), .B0_t (SubBytesIns_Inst_Sbox_10_T17), .B0_f (new_AGEMA_signal_7871), .B1_t (new_AGEMA_signal_7872), .B1_f (new_AGEMA_signal_7873), .Z0_t (SubBytesIns_Inst_Sbox_10_M51), .Z0_f (new_AGEMA_signal_10781), .Z1_t (new_AGEMA_signal_10782), .Z1_f (new_AGEMA_signal_10783) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M42), .A0_f (new_AGEMA_signal_10763), .A1_t (new_AGEMA_signal_10764), .A1_f (new_AGEMA_signal_10765), .B0_t (SubBytesIns_Inst_Sbox_10_T15), .B0_f (new_AGEMA_signal_7177), .B1_t (new_AGEMA_signal_7178), .B1_f (new_AGEMA_signal_7179), .Z0_t (SubBytesIns_Inst_Sbox_10_M52), .Z0_f (new_AGEMA_signal_11489), .Z1_t (new_AGEMA_signal_11490), .Z1_f (new_AGEMA_signal_11491) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M45), .A0_f (new_AGEMA_signal_11480), .A1_t (new_AGEMA_signal_11481), .A1_f (new_AGEMA_signal_11482), .B0_t (SubBytesIns_Inst_Sbox_10_T27), .B0_f (new_AGEMA_signal_7189), .B1_t (new_AGEMA_signal_7190), .B1_f (new_AGEMA_signal_7191), .Z0_t (SubBytesIns_Inst_Sbox_10_M53), .Z0_f (new_AGEMA_signal_12116), .Z1_t (new_AGEMA_signal_12117), .Z1_f (new_AGEMA_signal_12118) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M41), .A0_f (new_AGEMA_signal_10760), .A1_t (new_AGEMA_signal_10761), .A1_f (new_AGEMA_signal_10762), .B0_t (SubBytesIns_Inst_Sbox_10_T10), .B0_f (new_AGEMA_signal_7865), .B1_t (new_AGEMA_signal_7866), .B1_f (new_AGEMA_signal_7867), .Z0_t (SubBytesIns_Inst_Sbox_10_M54), .Z0_f (new_AGEMA_signal_11492), .Z1_t (new_AGEMA_signal_11493), .Z1_f (new_AGEMA_signal_11494) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M44), .A0_f (new_AGEMA_signal_10769), .A1_t (new_AGEMA_signal_10770), .A1_f (new_AGEMA_signal_10771), .B0_t (SubBytesIns_Inst_Sbox_10_T13), .B0_f (new_AGEMA_signal_7174), .B1_t (new_AGEMA_signal_7175), .B1_f (new_AGEMA_signal_7176), .Z0_t (SubBytesIns_Inst_Sbox_10_M55), .Z0_f (new_AGEMA_signal_11495), .Z1_t (new_AGEMA_signal_11496), .Z1_f (new_AGEMA_signal_11497) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M40), .A0_f (new_AGEMA_signal_10193), .A1_t (new_AGEMA_signal_10194), .A1_f (new_AGEMA_signal_10195), .B0_t (SubBytesIns_Inst_Sbox_10_T23), .B0_f (new_AGEMA_signal_7877), .B1_t (new_AGEMA_signal_7878), .B1_f (new_AGEMA_signal_7879), .Z0_t (SubBytesIns_Inst_Sbox_10_M56), .Z0_f (new_AGEMA_signal_10784), .Z1_t (new_AGEMA_signal_10785), .Z1_f (new_AGEMA_signal_10786) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M39), .A0_f (new_AGEMA_signal_10190), .A1_t (new_AGEMA_signal_10191), .A1_f (new_AGEMA_signal_10192), .B0_t (SubBytesIns_Inst_Sbox_10_T19), .B0_f (new_AGEMA_signal_7183), .B1_t (new_AGEMA_signal_7184), .B1_f (new_AGEMA_signal_7185), .Z0_t (SubBytesIns_Inst_Sbox_10_M57), .Z0_f (new_AGEMA_signal_10787), .Z1_t (new_AGEMA_signal_10788), .Z1_f (new_AGEMA_signal_10789) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M43), .A0_f (new_AGEMA_signal_10766), .A1_t (new_AGEMA_signal_10767), .A1_f (new_AGEMA_signal_10768), .B0_t (SubBytesIns_Inst_Sbox_10_T3), .B0_f (new_AGEMA_signal_6652), .B1_t (new_AGEMA_signal_6653), .B1_f (new_AGEMA_signal_6654), .Z0_t (SubBytesIns_Inst_Sbox_10_M58), .Z0_f (new_AGEMA_signal_11498), .Z1_t (new_AGEMA_signal_11499), .Z1_f (new_AGEMA_signal_11500) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M38), .A0_f (new_AGEMA_signal_10187), .A1_t (new_AGEMA_signal_10188), .A1_f (new_AGEMA_signal_10189), .B0_t (SubBytesIns_Inst_Sbox_10_T22), .B0_f (new_AGEMA_signal_7186), .B1_t (new_AGEMA_signal_7187), .B1_f (new_AGEMA_signal_7188), .Z0_t (SubBytesIns_Inst_Sbox_10_M59), .Z0_f (new_AGEMA_signal_10790), .Z1_t (new_AGEMA_signal_10791), .Z1_f (new_AGEMA_signal_10792) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M37), .A0_f (new_AGEMA_signal_10184), .A1_t (new_AGEMA_signal_10185), .A1_f (new_AGEMA_signal_10186), .B0_t (SubBytesIns_Inst_Sbox_10_T20), .B0_f (new_AGEMA_signal_7874), .B1_t (new_AGEMA_signal_7875), .B1_f (new_AGEMA_signal_7876), .Z0_t (SubBytesIns_Inst_Sbox_10_M60), .Z0_f (new_AGEMA_signal_10793), .Z1_t (new_AGEMA_signal_10794), .Z1_f (new_AGEMA_signal_10795) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M42), .A0_f (new_AGEMA_signal_10763), .A1_t (new_AGEMA_signal_10764), .A1_f (new_AGEMA_signal_10765), .B0_t (SubBytesIns_Inst_Sbox_10_T1), .B0_f (new_AGEMA_signal_6646), .B1_t (new_AGEMA_signal_6647), .B1_f (new_AGEMA_signal_6648), .Z0_t (SubBytesIns_Inst_Sbox_10_M61), .Z0_f (new_AGEMA_signal_11501), .Z1_t (new_AGEMA_signal_11502), .Z1_f (new_AGEMA_signal_11503) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M45), .A0_f (new_AGEMA_signal_11480), .A1_t (new_AGEMA_signal_11481), .A1_f (new_AGEMA_signal_11482), .B0_t (SubBytesIns_Inst_Sbox_10_T4), .B0_f (new_AGEMA_signal_6655), .B1_t (new_AGEMA_signal_6656), .B1_f (new_AGEMA_signal_6657), .Z0_t (SubBytesIns_Inst_Sbox_10_M62), .Z0_f (new_AGEMA_signal_12119), .Z1_t (new_AGEMA_signal_12120), .Z1_f (new_AGEMA_signal_12121) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M41), .A0_f (new_AGEMA_signal_10760), .A1_t (new_AGEMA_signal_10761), .A1_f (new_AGEMA_signal_10762), .B0_t (SubBytesIns_Inst_Sbox_10_T2), .B0_f (new_AGEMA_signal_6649), .B1_t (new_AGEMA_signal_6650), .B1_f (new_AGEMA_signal_6651), .Z0_t (SubBytesIns_Inst_Sbox_10_M63), .Z0_f (new_AGEMA_signal_11504), .Z1_t (new_AGEMA_signal_11505), .Z1_f (new_AGEMA_signal_11506) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M61), .A0_f (new_AGEMA_signal_11501), .A1_t (new_AGEMA_signal_11502), .A1_f (new_AGEMA_signal_11503), .B0_t (SubBytesIns_Inst_Sbox_10_M62), .B0_f (new_AGEMA_signal_12119), .B1_t (new_AGEMA_signal_12120), .B1_f (new_AGEMA_signal_12121), .Z0_t (SubBytesIns_Inst_Sbox_10_L0), .Z0_f (new_AGEMA_signal_12674), .Z1_t (new_AGEMA_signal_12675), .Z1_f (new_AGEMA_signal_12676) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M50), .A0_f (new_AGEMA_signal_10778), .A1_t (new_AGEMA_signal_10779), .A1_f (new_AGEMA_signal_10780), .B0_t (SubBytesIns_Inst_Sbox_10_M56), .B0_f (new_AGEMA_signal_10784), .B1_t (new_AGEMA_signal_10785), .B1_f (new_AGEMA_signal_10786), .Z0_t (SubBytesIns_Inst_Sbox_10_L1), .Z0_f (new_AGEMA_signal_11507), .Z1_t (new_AGEMA_signal_11508), .Z1_f (new_AGEMA_signal_11509) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M46), .A0_f (new_AGEMA_signal_11483), .A1_t (new_AGEMA_signal_11484), .A1_f (new_AGEMA_signal_11485), .B0_t (SubBytesIns_Inst_Sbox_10_M48), .B0_f (new_AGEMA_signal_10775), .B1_t (new_AGEMA_signal_10776), .B1_f (new_AGEMA_signal_10777), .Z0_t (SubBytesIns_Inst_Sbox_10_L2), .Z0_f (new_AGEMA_signal_12122), .Z1_t (new_AGEMA_signal_12123), .Z1_f (new_AGEMA_signal_12124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M47), .A0_f (new_AGEMA_signal_10772), .A1_t (new_AGEMA_signal_10773), .A1_f (new_AGEMA_signal_10774), .B0_t (SubBytesIns_Inst_Sbox_10_M55), .B0_f (new_AGEMA_signal_11495), .B1_t (new_AGEMA_signal_11496), .B1_f (new_AGEMA_signal_11497), .Z0_t (SubBytesIns_Inst_Sbox_10_L3), .Z0_f (new_AGEMA_signal_12125), .Z1_t (new_AGEMA_signal_12126), .Z1_f (new_AGEMA_signal_12127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M54), .A0_f (new_AGEMA_signal_11492), .A1_t (new_AGEMA_signal_11493), .A1_f (new_AGEMA_signal_11494), .B0_t (SubBytesIns_Inst_Sbox_10_M58), .B0_f (new_AGEMA_signal_11498), .B1_t (new_AGEMA_signal_11499), .B1_f (new_AGEMA_signal_11500), .Z0_t (SubBytesIns_Inst_Sbox_10_L4), .Z0_f (new_AGEMA_signal_12128), .Z1_t (new_AGEMA_signal_12129), .Z1_f (new_AGEMA_signal_12130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M49), .A0_f (new_AGEMA_signal_11486), .A1_t (new_AGEMA_signal_11487), .A1_f (new_AGEMA_signal_11488), .B0_t (SubBytesIns_Inst_Sbox_10_M61), .B0_f (new_AGEMA_signal_11501), .B1_t (new_AGEMA_signal_11502), .B1_f (new_AGEMA_signal_11503), .Z0_t (SubBytesIns_Inst_Sbox_10_L5), .Z0_f (new_AGEMA_signal_12131), .Z1_t (new_AGEMA_signal_12132), .Z1_f (new_AGEMA_signal_12133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M62), .A0_f (new_AGEMA_signal_12119), .A1_t (new_AGEMA_signal_12120), .A1_f (new_AGEMA_signal_12121), .B0_t (SubBytesIns_Inst_Sbox_10_L5), .B0_f (new_AGEMA_signal_12131), .B1_t (new_AGEMA_signal_12132), .B1_f (new_AGEMA_signal_12133), .Z0_t (SubBytesIns_Inst_Sbox_10_L6), .Z0_f (new_AGEMA_signal_12677), .Z1_t (new_AGEMA_signal_12678), .Z1_f (new_AGEMA_signal_12679) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M46), .A0_f (new_AGEMA_signal_11483), .A1_t (new_AGEMA_signal_11484), .A1_f (new_AGEMA_signal_11485), .B0_t (SubBytesIns_Inst_Sbox_10_L3), .B0_f (new_AGEMA_signal_12125), .B1_t (new_AGEMA_signal_12126), .B1_f (new_AGEMA_signal_12127), .Z0_t (SubBytesIns_Inst_Sbox_10_L7), .Z0_f (new_AGEMA_signal_12680), .Z1_t (new_AGEMA_signal_12681), .Z1_f (new_AGEMA_signal_12682) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M51), .A0_f (new_AGEMA_signal_10781), .A1_t (new_AGEMA_signal_10782), .A1_f (new_AGEMA_signal_10783), .B0_t (SubBytesIns_Inst_Sbox_10_M59), .B0_f (new_AGEMA_signal_10790), .B1_t (new_AGEMA_signal_10791), .B1_f (new_AGEMA_signal_10792), .Z0_t (SubBytesIns_Inst_Sbox_10_L8), .Z0_f (new_AGEMA_signal_11510), .Z1_t (new_AGEMA_signal_11511), .Z1_f (new_AGEMA_signal_11512) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M52), .A0_f (new_AGEMA_signal_11489), .A1_t (new_AGEMA_signal_11490), .A1_f (new_AGEMA_signal_11491), .B0_t (SubBytesIns_Inst_Sbox_10_M53), .B0_f (new_AGEMA_signal_12116), .B1_t (new_AGEMA_signal_12117), .B1_f (new_AGEMA_signal_12118), .Z0_t (SubBytesIns_Inst_Sbox_10_L9), .Z0_f (new_AGEMA_signal_12683), .Z1_t (new_AGEMA_signal_12684), .Z1_f (new_AGEMA_signal_12685) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M53), .A0_f (new_AGEMA_signal_12116), .A1_t (new_AGEMA_signal_12117), .A1_f (new_AGEMA_signal_12118), .B0_t (SubBytesIns_Inst_Sbox_10_L4), .B0_f (new_AGEMA_signal_12128), .B1_t (new_AGEMA_signal_12129), .B1_f (new_AGEMA_signal_12130), .Z0_t (SubBytesIns_Inst_Sbox_10_L10), .Z0_f (new_AGEMA_signal_12686), .Z1_t (new_AGEMA_signal_12687), .Z1_f (new_AGEMA_signal_12688) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M60), .A0_f (new_AGEMA_signal_10793), .A1_t (new_AGEMA_signal_10794), .A1_f (new_AGEMA_signal_10795), .B0_t (SubBytesIns_Inst_Sbox_10_L2), .B0_f (new_AGEMA_signal_12122), .B1_t (new_AGEMA_signal_12123), .B1_f (new_AGEMA_signal_12124), .Z0_t (SubBytesIns_Inst_Sbox_10_L11), .Z0_f (new_AGEMA_signal_12689), .Z1_t (new_AGEMA_signal_12690), .Z1_f (new_AGEMA_signal_12691) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M48), .A0_f (new_AGEMA_signal_10775), .A1_t (new_AGEMA_signal_10776), .A1_f (new_AGEMA_signal_10777), .B0_t (SubBytesIns_Inst_Sbox_10_M51), .B0_f (new_AGEMA_signal_10781), .B1_t (new_AGEMA_signal_10782), .B1_f (new_AGEMA_signal_10783), .Z0_t (SubBytesIns_Inst_Sbox_10_L12), .Z0_f (new_AGEMA_signal_11513), .Z1_t (new_AGEMA_signal_11514), .Z1_f (new_AGEMA_signal_11515) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M50), .A0_f (new_AGEMA_signal_10778), .A1_t (new_AGEMA_signal_10779), .A1_f (new_AGEMA_signal_10780), .B0_t (SubBytesIns_Inst_Sbox_10_L0), .B0_f (new_AGEMA_signal_12674), .B1_t (new_AGEMA_signal_12675), .B1_f (new_AGEMA_signal_12676), .Z0_t (SubBytesIns_Inst_Sbox_10_L13), .Z0_f (new_AGEMA_signal_13298), .Z1_t (new_AGEMA_signal_13299), .Z1_f (new_AGEMA_signal_13300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M52), .A0_f (new_AGEMA_signal_11489), .A1_t (new_AGEMA_signal_11490), .A1_f (new_AGEMA_signal_11491), .B0_t (SubBytesIns_Inst_Sbox_10_M61), .B0_f (new_AGEMA_signal_11501), .B1_t (new_AGEMA_signal_11502), .B1_f (new_AGEMA_signal_11503), .Z0_t (SubBytesIns_Inst_Sbox_10_L14), .Z0_f (new_AGEMA_signal_12134), .Z1_t (new_AGEMA_signal_12135), .Z1_f (new_AGEMA_signal_12136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M55), .A0_f (new_AGEMA_signal_11495), .A1_t (new_AGEMA_signal_11496), .A1_f (new_AGEMA_signal_11497), .B0_t (SubBytesIns_Inst_Sbox_10_L1), .B0_f (new_AGEMA_signal_11507), .B1_t (new_AGEMA_signal_11508), .B1_f (new_AGEMA_signal_11509), .Z0_t (SubBytesIns_Inst_Sbox_10_L15), .Z0_f (new_AGEMA_signal_12137), .Z1_t (new_AGEMA_signal_12138), .Z1_f (new_AGEMA_signal_12139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M56), .A0_f (new_AGEMA_signal_10784), .A1_t (new_AGEMA_signal_10785), .A1_f (new_AGEMA_signal_10786), .B0_t (SubBytesIns_Inst_Sbox_10_L0), .B0_f (new_AGEMA_signal_12674), .B1_t (new_AGEMA_signal_12675), .B1_f (new_AGEMA_signal_12676), .Z0_t (SubBytesIns_Inst_Sbox_10_L16), .Z0_f (new_AGEMA_signal_13301), .Z1_t (new_AGEMA_signal_13302), .Z1_f (new_AGEMA_signal_13303) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M57), .A0_f (new_AGEMA_signal_10787), .A1_t (new_AGEMA_signal_10788), .A1_f (new_AGEMA_signal_10789), .B0_t (SubBytesIns_Inst_Sbox_10_L1), .B0_f (new_AGEMA_signal_11507), .B1_t (new_AGEMA_signal_11508), .B1_f (new_AGEMA_signal_11509), .Z0_t (SubBytesIns_Inst_Sbox_10_L17), .Z0_f (new_AGEMA_signal_12140), .Z1_t (new_AGEMA_signal_12141), .Z1_f (new_AGEMA_signal_12142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M58), .A0_f (new_AGEMA_signal_11498), .A1_t (new_AGEMA_signal_11499), .A1_f (new_AGEMA_signal_11500), .B0_t (SubBytesIns_Inst_Sbox_10_L8), .B0_f (new_AGEMA_signal_11510), .B1_t (new_AGEMA_signal_11511), .B1_f (new_AGEMA_signal_11512), .Z0_t (SubBytesIns_Inst_Sbox_10_L18), .Z0_f (new_AGEMA_signal_12143), .Z1_t (new_AGEMA_signal_12144), .Z1_f (new_AGEMA_signal_12145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M63), .A0_f (new_AGEMA_signal_11504), .A1_t (new_AGEMA_signal_11505), .A1_f (new_AGEMA_signal_11506), .B0_t (SubBytesIns_Inst_Sbox_10_L4), .B0_f (new_AGEMA_signal_12128), .B1_t (new_AGEMA_signal_12129), .B1_f (new_AGEMA_signal_12130), .Z0_t (SubBytesIns_Inst_Sbox_10_L19), .Z0_f (new_AGEMA_signal_12692), .Z1_t (new_AGEMA_signal_12693), .Z1_f (new_AGEMA_signal_12694) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L0), .A0_f (new_AGEMA_signal_12674), .A1_t (new_AGEMA_signal_12675), .A1_f (new_AGEMA_signal_12676), .B0_t (SubBytesIns_Inst_Sbox_10_L1), .B0_f (new_AGEMA_signal_11507), .B1_t (new_AGEMA_signal_11508), .B1_f (new_AGEMA_signal_11509), .Z0_t (SubBytesIns_Inst_Sbox_10_L20), .Z0_f (new_AGEMA_signal_13304), .Z1_t (new_AGEMA_signal_13305), .Z1_f (new_AGEMA_signal_13306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L1), .A0_f (new_AGEMA_signal_11507), .A1_t (new_AGEMA_signal_11508), .A1_f (new_AGEMA_signal_11509), .B0_t (SubBytesIns_Inst_Sbox_10_L7), .B0_f (new_AGEMA_signal_12680), .B1_t (new_AGEMA_signal_12681), .B1_f (new_AGEMA_signal_12682), .Z0_t (SubBytesIns_Inst_Sbox_10_L21), .Z0_f (new_AGEMA_signal_13307), .Z1_t (new_AGEMA_signal_13308), .Z1_f (new_AGEMA_signal_13309) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L3), .A0_f (new_AGEMA_signal_12125), .A1_t (new_AGEMA_signal_12126), .A1_f (new_AGEMA_signal_12127), .B0_t (SubBytesIns_Inst_Sbox_10_L12), .B0_f (new_AGEMA_signal_11513), .B1_t (new_AGEMA_signal_11514), .B1_f (new_AGEMA_signal_11515), .Z0_t (SubBytesIns_Inst_Sbox_10_L22), .Z0_f (new_AGEMA_signal_12695), .Z1_t (new_AGEMA_signal_12696), .Z1_f (new_AGEMA_signal_12697) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L18), .A0_f (new_AGEMA_signal_12143), .A1_t (new_AGEMA_signal_12144), .A1_f (new_AGEMA_signal_12145), .B0_t (SubBytesIns_Inst_Sbox_10_L2), .B0_f (new_AGEMA_signal_12122), .B1_t (new_AGEMA_signal_12123), .B1_f (new_AGEMA_signal_12124), .Z0_t (SubBytesIns_Inst_Sbox_10_L23), .Z0_f (new_AGEMA_signal_12698), .Z1_t (new_AGEMA_signal_12699), .Z1_f (new_AGEMA_signal_12700) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L15), .A0_f (new_AGEMA_signal_12137), .A1_t (new_AGEMA_signal_12138), .A1_f (new_AGEMA_signal_12139), .B0_t (SubBytesIns_Inst_Sbox_10_L9), .B0_f (new_AGEMA_signal_12683), .B1_t (new_AGEMA_signal_12684), .B1_f (new_AGEMA_signal_12685), .Z0_t (SubBytesIns_Inst_Sbox_10_L24), .Z0_f (new_AGEMA_signal_13310), .Z1_t (new_AGEMA_signal_13311), .Z1_f (new_AGEMA_signal_13312) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L6), .A0_f (new_AGEMA_signal_12677), .A1_t (new_AGEMA_signal_12678), .A1_f (new_AGEMA_signal_12679), .B0_t (SubBytesIns_Inst_Sbox_10_L10), .B0_f (new_AGEMA_signal_12686), .B1_t (new_AGEMA_signal_12687), .B1_f (new_AGEMA_signal_12688), .Z0_t (SubBytesIns_Inst_Sbox_10_L25), .Z0_f (new_AGEMA_signal_13313), .Z1_t (new_AGEMA_signal_13314), .Z1_f (new_AGEMA_signal_13315) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L7), .A0_f (new_AGEMA_signal_12680), .A1_t (new_AGEMA_signal_12681), .A1_f (new_AGEMA_signal_12682), .B0_t (SubBytesIns_Inst_Sbox_10_L9), .B0_f (new_AGEMA_signal_12683), .B1_t (new_AGEMA_signal_12684), .B1_f (new_AGEMA_signal_12685), .Z0_t (SubBytesIns_Inst_Sbox_10_L26), .Z0_f (new_AGEMA_signal_13316), .Z1_t (new_AGEMA_signal_13317), .Z1_f (new_AGEMA_signal_13318) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L8), .A0_f (new_AGEMA_signal_11510), .A1_t (new_AGEMA_signal_11511), .A1_f (new_AGEMA_signal_11512), .B0_t (SubBytesIns_Inst_Sbox_10_L10), .B0_f (new_AGEMA_signal_12686), .B1_t (new_AGEMA_signal_12687), .B1_f (new_AGEMA_signal_12688), .Z0_t (SubBytesIns_Inst_Sbox_10_L27), .Z0_f (new_AGEMA_signal_13319), .Z1_t (new_AGEMA_signal_13320), .Z1_f (new_AGEMA_signal_13321) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L11), .A0_f (new_AGEMA_signal_12689), .A1_t (new_AGEMA_signal_12690), .A1_f (new_AGEMA_signal_12691), .B0_t (SubBytesIns_Inst_Sbox_10_L14), .B0_f (new_AGEMA_signal_12134), .B1_t (new_AGEMA_signal_12135), .B1_f (new_AGEMA_signal_12136), .Z0_t (SubBytesIns_Inst_Sbox_10_L28), .Z0_f (new_AGEMA_signal_13322), .Z1_t (new_AGEMA_signal_13323), .Z1_f (new_AGEMA_signal_13324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L11), .A0_f (new_AGEMA_signal_12689), .A1_t (new_AGEMA_signal_12690), .A1_f (new_AGEMA_signal_12691), .B0_t (SubBytesIns_Inst_Sbox_10_L17), .B0_f (new_AGEMA_signal_12140), .B1_t (new_AGEMA_signal_12141), .B1_f (new_AGEMA_signal_12142), .Z0_t (SubBytesIns_Inst_Sbox_10_L29), .Z0_f (new_AGEMA_signal_13325), .Z1_t (new_AGEMA_signal_13326), .Z1_f (new_AGEMA_signal_13327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L6), .A0_f (new_AGEMA_signal_12677), .A1_t (new_AGEMA_signal_12678), .A1_f (new_AGEMA_signal_12679), .B0_t (SubBytesIns_Inst_Sbox_10_L24), .B0_f (new_AGEMA_signal_13310), .B1_t (new_AGEMA_signal_13311), .B1_f (new_AGEMA_signal_13312), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .Z0_f (new_AGEMA_signal_13850), .Z1_t (new_AGEMA_signal_13851), .Z1_f (new_AGEMA_signal_13852) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L16), .A0_f (new_AGEMA_signal_13301), .A1_t (new_AGEMA_signal_13302), .A1_f (new_AGEMA_signal_13303), .B0_t (SubBytesIns_Inst_Sbox_10_L26), .B0_f (new_AGEMA_signal_13316), .B1_t (new_AGEMA_signal_13317), .B1_f (new_AGEMA_signal_13318), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .Z0_f (new_AGEMA_signal_13853), .Z1_t (new_AGEMA_signal_13854), .Z1_f (new_AGEMA_signal_13855) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L19), .A0_f (new_AGEMA_signal_12692), .A1_t (new_AGEMA_signal_12693), .A1_f (new_AGEMA_signal_12694), .B0_t (SubBytesIns_Inst_Sbox_10_L28), .B0_f (new_AGEMA_signal_13322), .B1_t (new_AGEMA_signal_13323), .B1_f (new_AGEMA_signal_13324), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .Z0_f (new_AGEMA_signal_13856), .Z1_t (new_AGEMA_signal_13857), .Z1_f (new_AGEMA_signal_13858) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L6), .A0_f (new_AGEMA_signal_12677), .A1_t (new_AGEMA_signal_12678), .A1_f (new_AGEMA_signal_12679), .B0_t (SubBytesIns_Inst_Sbox_10_L21), .B0_f (new_AGEMA_signal_13307), .B1_t (new_AGEMA_signal_13308), .B1_f (new_AGEMA_signal_13309), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .Z0_f (new_AGEMA_signal_13859), .Z1_t (new_AGEMA_signal_13860), .Z1_f (new_AGEMA_signal_13861) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L20), .A0_f (new_AGEMA_signal_13304), .A1_t (new_AGEMA_signal_13305), .A1_f (new_AGEMA_signal_13306), .B0_t (SubBytesIns_Inst_Sbox_10_L22), .B0_f (new_AGEMA_signal_12695), .B1_t (new_AGEMA_signal_12696), .B1_f (new_AGEMA_signal_12697), .Z0_t (MixColumnsInput[115]), .Z0_f (new_AGEMA_signal_13862), .Z1_t (new_AGEMA_signal_13863), .Z1_f (new_AGEMA_signal_13864) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L25), .A0_f (new_AGEMA_signal_13313), .A1_t (new_AGEMA_signal_13314), .A1_f (new_AGEMA_signal_13315), .B0_t (SubBytesIns_Inst_Sbox_10_L29), .B0_f (new_AGEMA_signal_13325), .B1_t (new_AGEMA_signal_13326), .B1_f (new_AGEMA_signal_13327), .Z0_t (MixColumnsInput[114]), .Z0_f (new_AGEMA_signal_13865), .Z1_t (new_AGEMA_signal_13866), .Z1_f (new_AGEMA_signal_13867) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L13), .A0_f (new_AGEMA_signal_13298), .A1_t (new_AGEMA_signal_13299), .A1_f (new_AGEMA_signal_13300), .B0_t (SubBytesIns_Inst_Sbox_10_L27), .B0_f (new_AGEMA_signal_13319), .B1_t (new_AGEMA_signal_13320), .B1_f (new_AGEMA_signal_13321), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .Z0_f (new_AGEMA_signal_13868), .Z1_t (new_AGEMA_signal_13869), .Z1_f (new_AGEMA_signal_13870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L6), .A0_f (new_AGEMA_signal_12677), .A1_t (new_AGEMA_signal_12678), .A1_f (new_AGEMA_signal_12679), .B0_t (SubBytesIns_Inst_Sbox_10_L23), .B0_f (new_AGEMA_signal_12698), .B1_t (new_AGEMA_signal_12699), .B1_f (new_AGEMA_signal_12700), .Z0_t (MixColumnsInput[112]), .Z0_f (new_AGEMA_signal_13328), .Z1_t (new_AGEMA_signal_13329), .Z1_f (new_AGEMA_signal_13330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[95]), .A0_f (ciphertext_s0_f[95]), .A1_t (ciphertext_s1_t[95]), .A1_f (ciphertext_s1_f[95]), .B0_t (ciphertext_s0_t[92]), .B0_f (ciphertext_s0_f[92]), .B1_t (ciphertext_s1_t[92]), .B1_f (ciphertext_s1_f[92]), .Z0_t (SubBytesIns_Inst_Sbox_11_T1), .Z0_f (new_AGEMA_signal_6676), .Z1_t (new_AGEMA_signal_6677), .Z1_f (new_AGEMA_signal_6678) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[95]), .A0_f (ciphertext_s0_f[95]), .A1_t (ciphertext_s1_t[95]), .A1_f (ciphertext_s1_f[95]), .B0_t (ciphertext_s0_t[90]), .B0_f (ciphertext_s0_f[90]), .B1_t (ciphertext_s1_t[90]), .B1_f (ciphertext_s1_f[90]), .Z0_t (SubBytesIns_Inst_Sbox_11_T2), .Z0_f (new_AGEMA_signal_6679), .Z1_t (new_AGEMA_signal_6680), .Z1_f (new_AGEMA_signal_6681) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[95]), .A0_f (ciphertext_s0_f[95]), .A1_t (ciphertext_s1_t[95]), .A1_f (ciphertext_s1_f[95]), .B0_t (ciphertext_s0_t[89]), .B0_f (ciphertext_s0_f[89]), .B1_t (ciphertext_s1_t[89]), .B1_f (ciphertext_s1_f[89]), .Z0_t (SubBytesIns_Inst_Sbox_11_T3), .Z0_f (new_AGEMA_signal_6682), .Z1_t (new_AGEMA_signal_6683), .Z1_f (new_AGEMA_signal_6684) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[92]), .A0_f (ciphertext_s0_f[92]), .A1_t (ciphertext_s1_t[92]), .A1_f (ciphertext_s1_f[92]), .B0_t (ciphertext_s0_t[90]), .B0_f (ciphertext_s0_f[90]), .B1_t (ciphertext_s1_t[90]), .B1_f (ciphertext_s1_f[90]), .Z0_t (SubBytesIns_Inst_Sbox_11_T4), .Z0_f (new_AGEMA_signal_6685), .Z1_t (new_AGEMA_signal_6686), .Z1_f (new_AGEMA_signal_6687) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[91]), .A0_f (ciphertext_s0_f[91]), .A1_t (ciphertext_s1_t[91]), .A1_f (ciphertext_s1_f[91]), .B0_t (ciphertext_s0_t[89]), .B0_f (ciphertext_s0_f[89]), .B1_t (ciphertext_s1_t[89]), .B1_f (ciphertext_s1_f[89]), .Z0_t (SubBytesIns_Inst_Sbox_11_T5), .Z0_f (new_AGEMA_signal_6688), .Z1_t (new_AGEMA_signal_6689), .Z1_f (new_AGEMA_signal_6690) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T1), .A0_f (new_AGEMA_signal_6676), .A1_t (new_AGEMA_signal_6677), .A1_f (new_AGEMA_signal_6678), .B0_t (SubBytesIns_Inst_Sbox_11_T5), .B0_f (new_AGEMA_signal_6688), .B1_t (new_AGEMA_signal_6689), .B1_f (new_AGEMA_signal_6690), .Z0_t (SubBytesIns_Inst_Sbox_11_T6), .Z0_f (new_AGEMA_signal_7192), .Z1_t (new_AGEMA_signal_7193), .Z1_f (new_AGEMA_signal_7194) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[94]), .A0_f (ciphertext_s0_f[94]), .A1_t (ciphertext_s1_t[94]), .A1_f (ciphertext_s1_f[94]), .B0_t (ciphertext_s0_t[93]), .B0_f (ciphertext_s0_f[93]), .B1_t (ciphertext_s1_t[93]), .B1_f (ciphertext_s1_f[93]), .Z0_t (SubBytesIns_Inst_Sbox_11_T7), .Z0_f (new_AGEMA_signal_6691), .Z1_t (new_AGEMA_signal_6692), .Z1_f (new_AGEMA_signal_6693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[88]), .A0_f (ciphertext_s0_f[88]), .A1_t (ciphertext_s1_t[88]), .A1_f (ciphertext_s1_f[88]), .B0_t (SubBytesIns_Inst_Sbox_11_T6), .B0_f (new_AGEMA_signal_7192), .B1_t (new_AGEMA_signal_7193), .B1_f (new_AGEMA_signal_7194), .Z0_t (SubBytesIns_Inst_Sbox_11_T8), .Z0_f (new_AGEMA_signal_7901), .Z1_t (new_AGEMA_signal_7902), .Z1_f (new_AGEMA_signal_7903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[88]), .A0_f (ciphertext_s0_f[88]), .A1_t (ciphertext_s1_t[88]), .A1_f (ciphertext_s1_f[88]), .B0_t (SubBytesIns_Inst_Sbox_11_T7), .B0_f (new_AGEMA_signal_6691), .B1_t (new_AGEMA_signal_6692), .B1_f (new_AGEMA_signal_6693), .Z0_t (SubBytesIns_Inst_Sbox_11_T9), .Z0_f (new_AGEMA_signal_7195), .Z1_t (new_AGEMA_signal_7196), .Z1_f (new_AGEMA_signal_7197) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T6), .A0_f (new_AGEMA_signal_7192), .A1_t (new_AGEMA_signal_7193), .A1_f (new_AGEMA_signal_7194), .B0_t (SubBytesIns_Inst_Sbox_11_T7), .B0_f (new_AGEMA_signal_6691), .B1_t (new_AGEMA_signal_6692), .B1_f (new_AGEMA_signal_6693), .Z0_t (SubBytesIns_Inst_Sbox_11_T10), .Z0_f (new_AGEMA_signal_7904), .Z1_t (new_AGEMA_signal_7905), .Z1_f (new_AGEMA_signal_7906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[94]), .A0_f (ciphertext_s0_f[94]), .A1_t (ciphertext_s1_t[94]), .A1_f (ciphertext_s1_f[94]), .B0_t (ciphertext_s0_t[90]), .B0_f (ciphertext_s0_f[90]), .B1_t (ciphertext_s1_t[90]), .B1_f (ciphertext_s1_f[90]), .Z0_t (SubBytesIns_Inst_Sbox_11_T11), .Z0_f (new_AGEMA_signal_6694), .Z1_t (new_AGEMA_signal_6695), .Z1_f (new_AGEMA_signal_6696) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[93]), .A0_f (ciphertext_s0_f[93]), .A1_t (ciphertext_s1_t[93]), .A1_f (ciphertext_s1_f[93]), .B0_t (ciphertext_s0_t[90]), .B0_f (ciphertext_s0_f[90]), .B1_t (ciphertext_s1_t[90]), .B1_f (ciphertext_s1_f[90]), .Z0_t (SubBytesIns_Inst_Sbox_11_T12), .Z0_f (new_AGEMA_signal_6697), .Z1_t (new_AGEMA_signal_6698), .Z1_f (new_AGEMA_signal_6699) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T3), .A0_f (new_AGEMA_signal_6682), .A1_t (new_AGEMA_signal_6683), .A1_f (new_AGEMA_signal_6684), .B0_t (SubBytesIns_Inst_Sbox_11_T4), .B0_f (new_AGEMA_signal_6685), .B1_t (new_AGEMA_signal_6686), .B1_f (new_AGEMA_signal_6687), .Z0_t (SubBytesIns_Inst_Sbox_11_T13), .Z0_f (new_AGEMA_signal_7198), .Z1_t (new_AGEMA_signal_7199), .Z1_f (new_AGEMA_signal_7200) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T6), .A0_f (new_AGEMA_signal_7192), .A1_t (new_AGEMA_signal_7193), .A1_f (new_AGEMA_signal_7194), .B0_t (SubBytesIns_Inst_Sbox_11_T11), .B0_f (new_AGEMA_signal_6694), .B1_t (new_AGEMA_signal_6695), .B1_f (new_AGEMA_signal_6696), .Z0_t (SubBytesIns_Inst_Sbox_11_T14), .Z0_f (new_AGEMA_signal_7907), .Z1_t (new_AGEMA_signal_7908), .Z1_f (new_AGEMA_signal_7909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T5), .A0_f (new_AGEMA_signal_6688), .A1_t (new_AGEMA_signal_6689), .A1_f (new_AGEMA_signal_6690), .B0_t (SubBytesIns_Inst_Sbox_11_T11), .B0_f (new_AGEMA_signal_6694), .B1_t (new_AGEMA_signal_6695), .B1_f (new_AGEMA_signal_6696), .Z0_t (SubBytesIns_Inst_Sbox_11_T15), .Z0_f (new_AGEMA_signal_7201), .Z1_t (new_AGEMA_signal_7202), .Z1_f (new_AGEMA_signal_7203) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T5), .A0_f (new_AGEMA_signal_6688), .A1_t (new_AGEMA_signal_6689), .A1_f (new_AGEMA_signal_6690), .B0_t (SubBytesIns_Inst_Sbox_11_T12), .B0_f (new_AGEMA_signal_6697), .B1_t (new_AGEMA_signal_6698), .B1_f (new_AGEMA_signal_6699), .Z0_t (SubBytesIns_Inst_Sbox_11_T16), .Z0_f (new_AGEMA_signal_7204), .Z1_t (new_AGEMA_signal_7205), .Z1_f (new_AGEMA_signal_7206) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T9), .A0_f (new_AGEMA_signal_7195), .A1_t (new_AGEMA_signal_7196), .A1_f (new_AGEMA_signal_7197), .B0_t (SubBytesIns_Inst_Sbox_11_T16), .B0_f (new_AGEMA_signal_7204), .B1_t (new_AGEMA_signal_7205), .B1_f (new_AGEMA_signal_7206), .Z0_t (SubBytesIns_Inst_Sbox_11_T17), .Z0_f (new_AGEMA_signal_7910), .Z1_t (new_AGEMA_signal_7911), .Z1_f (new_AGEMA_signal_7912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[92]), .A0_f (ciphertext_s0_f[92]), .A1_t (ciphertext_s1_t[92]), .A1_f (ciphertext_s1_f[92]), .B0_t (ciphertext_s0_t[88]), .B0_f (ciphertext_s0_f[88]), .B1_t (ciphertext_s1_t[88]), .B1_f (ciphertext_s1_f[88]), .Z0_t (SubBytesIns_Inst_Sbox_11_T18), .Z0_f (new_AGEMA_signal_6700), .Z1_t (new_AGEMA_signal_6701), .Z1_f (new_AGEMA_signal_6702) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T7), .A0_f (new_AGEMA_signal_6691), .A1_t (new_AGEMA_signal_6692), .A1_f (new_AGEMA_signal_6693), .B0_t (SubBytesIns_Inst_Sbox_11_T18), .B0_f (new_AGEMA_signal_6700), .B1_t (new_AGEMA_signal_6701), .B1_f (new_AGEMA_signal_6702), .Z0_t (SubBytesIns_Inst_Sbox_11_T19), .Z0_f (new_AGEMA_signal_7207), .Z1_t (new_AGEMA_signal_7208), .Z1_f (new_AGEMA_signal_7209) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T1), .A0_f (new_AGEMA_signal_6676), .A1_t (new_AGEMA_signal_6677), .A1_f (new_AGEMA_signal_6678), .B0_t (SubBytesIns_Inst_Sbox_11_T19), .B0_f (new_AGEMA_signal_7207), .B1_t (new_AGEMA_signal_7208), .B1_f (new_AGEMA_signal_7209), .Z0_t (SubBytesIns_Inst_Sbox_11_T20), .Z0_f (new_AGEMA_signal_7913), .Z1_t (new_AGEMA_signal_7914), .Z1_f (new_AGEMA_signal_7915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[89]), .A0_f (ciphertext_s0_f[89]), .A1_t (ciphertext_s1_t[89]), .A1_f (ciphertext_s1_f[89]), .B0_t (ciphertext_s0_t[88]), .B0_f (ciphertext_s0_f[88]), .B1_t (ciphertext_s1_t[88]), .B1_f (ciphertext_s1_f[88]), .Z0_t (SubBytesIns_Inst_Sbox_11_T21), .Z0_f (new_AGEMA_signal_6703), .Z1_t (new_AGEMA_signal_6704), .Z1_f (new_AGEMA_signal_6705) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T7), .A0_f (new_AGEMA_signal_6691), .A1_t (new_AGEMA_signal_6692), .A1_f (new_AGEMA_signal_6693), .B0_t (SubBytesIns_Inst_Sbox_11_T21), .B0_f (new_AGEMA_signal_6703), .B1_t (new_AGEMA_signal_6704), .B1_f (new_AGEMA_signal_6705), .Z0_t (SubBytesIns_Inst_Sbox_11_T22), .Z0_f (new_AGEMA_signal_7210), .Z1_t (new_AGEMA_signal_7211), .Z1_f (new_AGEMA_signal_7212) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T2), .A0_f (new_AGEMA_signal_6679), .A1_t (new_AGEMA_signal_6680), .A1_f (new_AGEMA_signal_6681), .B0_t (SubBytesIns_Inst_Sbox_11_T22), .B0_f (new_AGEMA_signal_7210), .B1_t (new_AGEMA_signal_7211), .B1_f (new_AGEMA_signal_7212), .Z0_t (SubBytesIns_Inst_Sbox_11_T23), .Z0_f (new_AGEMA_signal_7916), .Z1_t (new_AGEMA_signal_7917), .Z1_f (new_AGEMA_signal_7918) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T2), .A0_f (new_AGEMA_signal_6679), .A1_t (new_AGEMA_signal_6680), .A1_f (new_AGEMA_signal_6681), .B0_t (SubBytesIns_Inst_Sbox_11_T10), .B0_f (new_AGEMA_signal_7904), .B1_t (new_AGEMA_signal_7905), .B1_f (new_AGEMA_signal_7906), .Z0_t (SubBytesIns_Inst_Sbox_11_T24), .Z0_f (new_AGEMA_signal_8501), .Z1_t (new_AGEMA_signal_8502), .Z1_f (new_AGEMA_signal_8503) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T20), .A0_f (new_AGEMA_signal_7913), .A1_t (new_AGEMA_signal_7914), .A1_f (new_AGEMA_signal_7915), .B0_t (SubBytesIns_Inst_Sbox_11_T17), .B0_f (new_AGEMA_signal_7910), .B1_t (new_AGEMA_signal_7911), .B1_f (new_AGEMA_signal_7912), .Z0_t (SubBytesIns_Inst_Sbox_11_T25), .Z0_f (new_AGEMA_signal_8504), .Z1_t (new_AGEMA_signal_8505), .Z1_f (new_AGEMA_signal_8506) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T3), .A0_f (new_AGEMA_signal_6682), .A1_t (new_AGEMA_signal_6683), .A1_f (new_AGEMA_signal_6684), .B0_t (SubBytesIns_Inst_Sbox_11_T16), .B0_f (new_AGEMA_signal_7204), .B1_t (new_AGEMA_signal_7205), .B1_f (new_AGEMA_signal_7206), .Z0_t (SubBytesIns_Inst_Sbox_11_T26), .Z0_f (new_AGEMA_signal_7919), .Z1_t (new_AGEMA_signal_7920), .Z1_f (new_AGEMA_signal_7921) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T1), .A0_f (new_AGEMA_signal_6676), .A1_t (new_AGEMA_signal_6677), .A1_f (new_AGEMA_signal_6678), .B0_t (SubBytesIns_Inst_Sbox_11_T12), .B0_f (new_AGEMA_signal_6697), .B1_t (new_AGEMA_signal_6698), .B1_f (new_AGEMA_signal_6699), .Z0_t (SubBytesIns_Inst_Sbox_11_T27), .Z0_f (new_AGEMA_signal_7213), .Z1_t (new_AGEMA_signal_7214), .Z1_f (new_AGEMA_signal_7215) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T13), .A0_f (new_AGEMA_signal_7198), .A1_t (new_AGEMA_signal_7199), .A1_f (new_AGEMA_signal_7200), .B0_t (SubBytesIns_Inst_Sbox_11_T6), .B0_f (new_AGEMA_signal_7192), .B1_t (new_AGEMA_signal_7193), .B1_f (new_AGEMA_signal_7194), .Z0_t (SubBytesIns_Inst_Sbox_11_M1), .Z0_f (new_AGEMA_signal_7922), .Z1_t (new_AGEMA_signal_7923), .Z1_f (new_AGEMA_signal_7924) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T23), .A0_f (new_AGEMA_signal_7916), .A1_t (new_AGEMA_signal_7917), .A1_f (new_AGEMA_signal_7918), .B0_t (SubBytesIns_Inst_Sbox_11_T8), .B0_f (new_AGEMA_signal_7901), .B1_t (new_AGEMA_signal_7902), .B1_f (new_AGEMA_signal_7903), .Z0_t (SubBytesIns_Inst_Sbox_11_M2), .Z0_f (new_AGEMA_signal_8507), .Z1_t (new_AGEMA_signal_8508), .Z1_f (new_AGEMA_signal_8509) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T14), .A0_f (new_AGEMA_signal_7907), .A1_t (new_AGEMA_signal_7908), .A1_f (new_AGEMA_signal_7909), .B0_t (SubBytesIns_Inst_Sbox_11_M1), .B0_f (new_AGEMA_signal_7922), .B1_t (new_AGEMA_signal_7923), .B1_f (new_AGEMA_signal_7924), .Z0_t (SubBytesIns_Inst_Sbox_11_M3), .Z0_f (new_AGEMA_signal_8510), .Z1_t (new_AGEMA_signal_8511), .Z1_f (new_AGEMA_signal_8512) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T19), .A0_f (new_AGEMA_signal_7207), .A1_t (new_AGEMA_signal_7208), .A1_f (new_AGEMA_signal_7209), .B0_t (ciphertext_s0_t[88]), .B0_f (ciphertext_s0_f[88]), .B1_t (ciphertext_s1_t[88]), .B1_f (ciphertext_s1_f[88]), .Z0_t (SubBytesIns_Inst_Sbox_11_M4), .Z0_f (new_AGEMA_signal_7925), .Z1_t (new_AGEMA_signal_7926), .Z1_f (new_AGEMA_signal_7927) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M4), .A0_f (new_AGEMA_signal_7925), .A1_t (new_AGEMA_signal_7926), .A1_f (new_AGEMA_signal_7927), .B0_t (SubBytesIns_Inst_Sbox_11_M1), .B0_f (new_AGEMA_signal_7922), .B1_t (new_AGEMA_signal_7923), .B1_f (new_AGEMA_signal_7924), .Z0_t (SubBytesIns_Inst_Sbox_11_M5), .Z0_f (new_AGEMA_signal_8513), .Z1_t (new_AGEMA_signal_8514), .Z1_f (new_AGEMA_signal_8515) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T3), .A0_f (new_AGEMA_signal_6682), .A1_t (new_AGEMA_signal_6683), .A1_f (new_AGEMA_signal_6684), .B0_t (SubBytesIns_Inst_Sbox_11_T16), .B0_f (new_AGEMA_signal_7204), .B1_t (new_AGEMA_signal_7205), .B1_f (new_AGEMA_signal_7206), .Z0_t (SubBytesIns_Inst_Sbox_11_M6), .Z0_f (new_AGEMA_signal_7928), .Z1_t (new_AGEMA_signal_7929), .Z1_f (new_AGEMA_signal_7930) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T22), .A0_f (new_AGEMA_signal_7210), .A1_t (new_AGEMA_signal_7211), .A1_f (new_AGEMA_signal_7212), .B0_t (SubBytesIns_Inst_Sbox_11_T9), .B0_f (new_AGEMA_signal_7195), .B1_t (new_AGEMA_signal_7196), .B1_f (new_AGEMA_signal_7197), .Z0_t (SubBytesIns_Inst_Sbox_11_M7), .Z0_f (new_AGEMA_signal_7931), .Z1_t (new_AGEMA_signal_7932), .Z1_f (new_AGEMA_signal_7933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T26), .A0_f (new_AGEMA_signal_7919), .A1_t (new_AGEMA_signal_7920), .A1_f (new_AGEMA_signal_7921), .B0_t (SubBytesIns_Inst_Sbox_11_M6), .B0_f (new_AGEMA_signal_7928), .B1_t (new_AGEMA_signal_7929), .B1_f (new_AGEMA_signal_7930), .Z0_t (SubBytesIns_Inst_Sbox_11_M8), .Z0_f (new_AGEMA_signal_8516), .Z1_t (new_AGEMA_signal_8517), .Z1_f (new_AGEMA_signal_8518) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T20), .A0_f (new_AGEMA_signal_7913), .A1_t (new_AGEMA_signal_7914), .A1_f (new_AGEMA_signal_7915), .B0_t (SubBytesIns_Inst_Sbox_11_T17), .B0_f (new_AGEMA_signal_7910), .B1_t (new_AGEMA_signal_7911), .B1_f (new_AGEMA_signal_7912), .Z0_t (SubBytesIns_Inst_Sbox_11_M9), .Z0_f (new_AGEMA_signal_8519), .Z1_t (new_AGEMA_signal_8520), .Z1_f (new_AGEMA_signal_8521) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M9), .A0_f (new_AGEMA_signal_8519), .A1_t (new_AGEMA_signal_8520), .A1_f (new_AGEMA_signal_8521), .B0_t (SubBytesIns_Inst_Sbox_11_M6), .B0_f (new_AGEMA_signal_7928), .B1_t (new_AGEMA_signal_7929), .B1_f (new_AGEMA_signal_7930), .Z0_t (SubBytesIns_Inst_Sbox_11_M10), .Z0_f (new_AGEMA_signal_8861), .Z1_t (new_AGEMA_signal_8862), .Z1_f (new_AGEMA_signal_8863) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T1), .A0_f (new_AGEMA_signal_6676), .A1_t (new_AGEMA_signal_6677), .A1_f (new_AGEMA_signal_6678), .B0_t (SubBytesIns_Inst_Sbox_11_T15), .B0_f (new_AGEMA_signal_7201), .B1_t (new_AGEMA_signal_7202), .B1_f (new_AGEMA_signal_7203), .Z0_t (SubBytesIns_Inst_Sbox_11_M11), .Z0_f (new_AGEMA_signal_7934), .Z1_t (new_AGEMA_signal_7935), .Z1_f (new_AGEMA_signal_7936) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T4), .A0_f (new_AGEMA_signal_6685), .A1_t (new_AGEMA_signal_6686), .A1_f (new_AGEMA_signal_6687), .B0_t (SubBytesIns_Inst_Sbox_11_T27), .B0_f (new_AGEMA_signal_7213), .B1_t (new_AGEMA_signal_7214), .B1_f (new_AGEMA_signal_7215), .Z0_t (SubBytesIns_Inst_Sbox_11_M12), .Z0_f (new_AGEMA_signal_7937), .Z1_t (new_AGEMA_signal_7938), .Z1_f (new_AGEMA_signal_7939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M12), .A0_f (new_AGEMA_signal_7937), .A1_t (new_AGEMA_signal_7938), .A1_f (new_AGEMA_signal_7939), .B0_t (SubBytesIns_Inst_Sbox_11_M11), .B0_f (new_AGEMA_signal_7934), .B1_t (new_AGEMA_signal_7935), .B1_f (new_AGEMA_signal_7936), .Z0_t (SubBytesIns_Inst_Sbox_11_M13), .Z0_f (new_AGEMA_signal_8522), .Z1_t (new_AGEMA_signal_8523), .Z1_f (new_AGEMA_signal_8524) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T2), .A0_f (new_AGEMA_signal_6679), .A1_t (new_AGEMA_signal_6680), .A1_f (new_AGEMA_signal_6681), .B0_t (SubBytesIns_Inst_Sbox_11_T10), .B0_f (new_AGEMA_signal_7904), .B1_t (new_AGEMA_signal_7905), .B1_f (new_AGEMA_signal_7906), .Z0_t (SubBytesIns_Inst_Sbox_11_M14), .Z0_f (new_AGEMA_signal_8525), .Z1_t (new_AGEMA_signal_8526), .Z1_f (new_AGEMA_signal_8527) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M14), .A0_f (new_AGEMA_signal_8525), .A1_t (new_AGEMA_signal_8526), .A1_f (new_AGEMA_signal_8527), .B0_t (SubBytesIns_Inst_Sbox_11_M11), .B0_f (new_AGEMA_signal_7934), .B1_t (new_AGEMA_signal_7935), .B1_f (new_AGEMA_signal_7936), .Z0_t (SubBytesIns_Inst_Sbox_11_M15), .Z0_f (new_AGEMA_signal_8864), .Z1_t (new_AGEMA_signal_8865), .Z1_f (new_AGEMA_signal_8866) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M3), .A0_f (new_AGEMA_signal_8510), .A1_t (new_AGEMA_signal_8511), .A1_f (new_AGEMA_signal_8512), .B0_t (SubBytesIns_Inst_Sbox_11_M2), .B0_f (new_AGEMA_signal_8507), .B1_t (new_AGEMA_signal_8508), .B1_f (new_AGEMA_signal_8509), .Z0_t (SubBytesIns_Inst_Sbox_11_M16), .Z0_f (new_AGEMA_signal_8867), .Z1_t (new_AGEMA_signal_8868), .Z1_f (new_AGEMA_signal_8869) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M5), .A0_f (new_AGEMA_signal_8513), .A1_t (new_AGEMA_signal_8514), .A1_f (new_AGEMA_signal_8515), .B0_t (SubBytesIns_Inst_Sbox_11_T24), .B0_f (new_AGEMA_signal_8501), .B1_t (new_AGEMA_signal_8502), .B1_f (new_AGEMA_signal_8503), .Z0_t (SubBytesIns_Inst_Sbox_11_M17), .Z0_f (new_AGEMA_signal_8870), .Z1_t (new_AGEMA_signal_8871), .Z1_f (new_AGEMA_signal_8872) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M8), .A0_f (new_AGEMA_signal_8516), .A1_t (new_AGEMA_signal_8517), .A1_f (new_AGEMA_signal_8518), .B0_t (SubBytesIns_Inst_Sbox_11_M7), .B0_f (new_AGEMA_signal_7931), .B1_t (new_AGEMA_signal_7932), .B1_f (new_AGEMA_signal_7933), .Z0_t (SubBytesIns_Inst_Sbox_11_M18), .Z0_f (new_AGEMA_signal_8873), .Z1_t (new_AGEMA_signal_8874), .Z1_f (new_AGEMA_signal_8875) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M10), .A0_f (new_AGEMA_signal_8861), .A1_t (new_AGEMA_signal_8862), .A1_f (new_AGEMA_signal_8863), .B0_t (SubBytesIns_Inst_Sbox_11_M15), .B0_f (new_AGEMA_signal_8864), .B1_t (new_AGEMA_signal_8865), .B1_f (new_AGEMA_signal_8866), .Z0_t (SubBytesIns_Inst_Sbox_11_M19), .Z0_f (new_AGEMA_signal_9116), .Z1_t (new_AGEMA_signal_9117), .Z1_f (new_AGEMA_signal_9118) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M16), .A0_f (new_AGEMA_signal_8867), .A1_t (new_AGEMA_signal_8868), .A1_f (new_AGEMA_signal_8869), .B0_t (SubBytesIns_Inst_Sbox_11_M13), .B0_f (new_AGEMA_signal_8522), .B1_t (new_AGEMA_signal_8523), .B1_f (new_AGEMA_signal_8524), .Z0_t (SubBytesIns_Inst_Sbox_11_M20), .Z0_f (new_AGEMA_signal_9119), .Z1_t (new_AGEMA_signal_9120), .Z1_f (new_AGEMA_signal_9121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M17), .A0_f (new_AGEMA_signal_8870), .A1_t (new_AGEMA_signal_8871), .A1_f (new_AGEMA_signal_8872), .B0_t (SubBytesIns_Inst_Sbox_11_M15), .B0_f (new_AGEMA_signal_8864), .B1_t (new_AGEMA_signal_8865), .B1_f (new_AGEMA_signal_8866), .Z0_t (SubBytesIns_Inst_Sbox_11_M21), .Z0_f (new_AGEMA_signal_9122), .Z1_t (new_AGEMA_signal_9123), .Z1_f (new_AGEMA_signal_9124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M18), .A0_f (new_AGEMA_signal_8873), .A1_t (new_AGEMA_signal_8874), .A1_f (new_AGEMA_signal_8875), .B0_t (SubBytesIns_Inst_Sbox_11_M13), .B0_f (new_AGEMA_signal_8522), .B1_t (new_AGEMA_signal_8523), .B1_f (new_AGEMA_signal_8524), .Z0_t (SubBytesIns_Inst_Sbox_11_M22), .Z0_f (new_AGEMA_signal_9125), .Z1_t (new_AGEMA_signal_9126), .Z1_f (new_AGEMA_signal_9127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M19), .A0_f (new_AGEMA_signal_9116), .A1_t (new_AGEMA_signal_9117), .A1_f (new_AGEMA_signal_9118), .B0_t (SubBytesIns_Inst_Sbox_11_T25), .B0_f (new_AGEMA_signal_8504), .B1_t (new_AGEMA_signal_8505), .B1_f (new_AGEMA_signal_8506), .Z0_t (SubBytesIns_Inst_Sbox_11_M23), .Z0_f (new_AGEMA_signal_9356), .Z1_t (new_AGEMA_signal_9357), .Z1_f (new_AGEMA_signal_9358) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M22), .A0_f (new_AGEMA_signal_9125), .A1_t (new_AGEMA_signal_9126), .A1_f (new_AGEMA_signal_9127), .B0_t (SubBytesIns_Inst_Sbox_11_M23), .B0_f (new_AGEMA_signal_9356), .B1_t (new_AGEMA_signal_9357), .B1_f (new_AGEMA_signal_9358), .Z0_t (SubBytesIns_Inst_Sbox_11_M24), .Z0_f (new_AGEMA_signal_9641), .Z1_t (new_AGEMA_signal_9642), .Z1_f (new_AGEMA_signal_9643) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M22), .A0_f (new_AGEMA_signal_9125), .A1_t (new_AGEMA_signal_9126), .A1_f (new_AGEMA_signal_9127), .B0_t (SubBytesIns_Inst_Sbox_11_M20), .B0_f (new_AGEMA_signal_9119), .B1_t (new_AGEMA_signal_9120), .B1_f (new_AGEMA_signal_9121), .Z0_t (SubBytesIns_Inst_Sbox_11_M25), .Z0_f (new_AGEMA_signal_9359), .Z1_t (new_AGEMA_signal_9360), .Z1_f (new_AGEMA_signal_9361) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M21), .A0_f (new_AGEMA_signal_9122), .A1_t (new_AGEMA_signal_9123), .A1_f (new_AGEMA_signal_9124), .B0_t (SubBytesIns_Inst_Sbox_11_M25), .B0_f (new_AGEMA_signal_9359), .B1_t (new_AGEMA_signal_9360), .B1_f (new_AGEMA_signal_9361), .Z0_t (SubBytesIns_Inst_Sbox_11_M26), .Z0_f (new_AGEMA_signal_9644), .Z1_t (new_AGEMA_signal_9645), .Z1_f (new_AGEMA_signal_9646) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M20), .A0_f (new_AGEMA_signal_9119), .A1_t (new_AGEMA_signal_9120), .A1_f (new_AGEMA_signal_9121), .B0_t (SubBytesIns_Inst_Sbox_11_M21), .B0_f (new_AGEMA_signal_9122), .B1_t (new_AGEMA_signal_9123), .B1_f (new_AGEMA_signal_9124), .Z0_t (SubBytesIns_Inst_Sbox_11_M27), .Z0_f (new_AGEMA_signal_9362), .Z1_t (new_AGEMA_signal_9363), .Z1_f (new_AGEMA_signal_9364) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M23), .A0_f (new_AGEMA_signal_9356), .A1_t (new_AGEMA_signal_9357), .A1_f (new_AGEMA_signal_9358), .B0_t (SubBytesIns_Inst_Sbox_11_M25), .B0_f (new_AGEMA_signal_9359), .B1_t (new_AGEMA_signal_9360), .B1_f (new_AGEMA_signal_9361), .Z0_t (SubBytesIns_Inst_Sbox_11_M28), .Z0_f (new_AGEMA_signal_9647), .Z1_t (new_AGEMA_signal_9648), .Z1_f (new_AGEMA_signal_9649) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M28), .A0_f (new_AGEMA_signal_9647), .A1_t (new_AGEMA_signal_9648), .A1_f (new_AGEMA_signal_9649), .B0_t (SubBytesIns_Inst_Sbox_11_M27), .B0_f (new_AGEMA_signal_9362), .B1_t (new_AGEMA_signal_9363), .B1_f (new_AGEMA_signal_9364), .Z0_t (SubBytesIns_Inst_Sbox_11_M29), .Z0_f (new_AGEMA_signal_9941), .Z1_t (new_AGEMA_signal_9942), .Z1_f (new_AGEMA_signal_9943) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M26), .A0_f (new_AGEMA_signal_9644), .A1_t (new_AGEMA_signal_9645), .A1_f (new_AGEMA_signal_9646), .B0_t (SubBytesIns_Inst_Sbox_11_M24), .B0_f (new_AGEMA_signal_9641), .B1_t (new_AGEMA_signal_9642), .B1_f (new_AGEMA_signal_9643), .Z0_t (SubBytesIns_Inst_Sbox_11_M30), .Z0_f (new_AGEMA_signal_9944), .Z1_t (new_AGEMA_signal_9945), .Z1_f (new_AGEMA_signal_9946) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M20), .A0_f (new_AGEMA_signal_9119), .A1_t (new_AGEMA_signal_9120), .A1_f (new_AGEMA_signal_9121), .B0_t (SubBytesIns_Inst_Sbox_11_M23), .B0_f (new_AGEMA_signal_9356), .B1_t (new_AGEMA_signal_9357), .B1_f (new_AGEMA_signal_9358), .Z0_t (SubBytesIns_Inst_Sbox_11_M31), .Z0_f (new_AGEMA_signal_9650), .Z1_t (new_AGEMA_signal_9651), .Z1_f (new_AGEMA_signal_9652) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M27), .A0_f (new_AGEMA_signal_9362), .A1_t (new_AGEMA_signal_9363), .A1_f (new_AGEMA_signal_9364), .B0_t (SubBytesIns_Inst_Sbox_11_M31), .B0_f (new_AGEMA_signal_9650), .B1_t (new_AGEMA_signal_9651), .B1_f (new_AGEMA_signal_9652), .Z0_t (SubBytesIns_Inst_Sbox_11_M32), .Z0_f (new_AGEMA_signal_9947), .Z1_t (new_AGEMA_signal_9948), .Z1_f (new_AGEMA_signal_9949) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M27), .A0_f (new_AGEMA_signal_9362), .A1_t (new_AGEMA_signal_9363), .A1_f (new_AGEMA_signal_9364), .B0_t (SubBytesIns_Inst_Sbox_11_M25), .B0_f (new_AGEMA_signal_9359), .B1_t (new_AGEMA_signal_9360), .B1_f (new_AGEMA_signal_9361), .Z0_t (SubBytesIns_Inst_Sbox_11_M33), .Z0_f (new_AGEMA_signal_9653), .Z1_t (new_AGEMA_signal_9654), .Z1_f (new_AGEMA_signal_9655) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M21), .A0_f (new_AGEMA_signal_9122), .A1_t (new_AGEMA_signal_9123), .A1_f (new_AGEMA_signal_9124), .B0_t (SubBytesIns_Inst_Sbox_11_M22), .B0_f (new_AGEMA_signal_9125), .B1_t (new_AGEMA_signal_9126), .B1_f (new_AGEMA_signal_9127), .Z0_t (SubBytesIns_Inst_Sbox_11_M34), .Z0_f (new_AGEMA_signal_9365), .Z1_t (new_AGEMA_signal_9366), .Z1_f (new_AGEMA_signal_9367) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M24), .A0_f (new_AGEMA_signal_9641), .A1_t (new_AGEMA_signal_9642), .A1_f (new_AGEMA_signal_9643), .B0_t (SubBytesIns_Inst_Sbox_11_M34), .B0_f (new_AGEMA_signal_9365), .B1_t (new_AGEMA_signal_9366), .B1_f (new_AGEMA_signal_9367), .Z0_t (SubBytesIns_Inst_Sbox_11_M35), .Z0_f (new_AGEMA_signal_9950), .Z1_t (new_AGEMA_signal_9951), .Z1_f (new_AGEMA_signal_9952) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M24), .A0_f (new_AGEMA_signal_9641), .A1_t (new_AGEMA_signal_9642), .A1_f (new_AGEMA_signal_9643), .B0_t (SubBytesIns_Inst_Sbox_11_M25), .B0_f (new_AGEMA_signal_9359), .B1_t (new_AGEMA_signal_9360), .B1_f (new_AGEMA_signal_9361), .Z0_t (SubBytesIns_Inst_Sbox_11_M36), .Z0_f (new_AGEMA_signal_9953), .Z1_t (new_AGEMA_signal_9954), .Z1_f (new_AGEMA_signal_9955) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M21), .A0_f (new_AGEMA_signal_9122), .A1_t (new_AGEMA_signal_9123), .A1_f (new_AGEMA_signal_9124), .B0_t (SubBytesIns_Inst_Sbox_11_M29), .B0_f (new_AGEMA_signal_9941), .B1_t (new_AGEMA_signal_9942), .B1_f (new_AGEMA_signal_9943), .Z0_t (SubBytesIns_Inst_Sbox_11_M37), .Z0_f (new_AGEMA_signal_10196), .Z1_t (new_AGEMA_signal_10197), .Z1_f (new_AGEMA_signal_10198) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M32), .A0_f (new_AGEMA_signal_9947), .A1_t (new_AGEMA_signal_9948), .A1_f (new_AGEMA_signal_9949), .B0_t (SubBytesIns_Inst_Sbox_11_M33), .B0_f (new_AGEMA_signal_9653), .B1_t (new_AGEMA_signal_9654), .B1_f (new_AGEMA_signal_9655), .Z0_t (SubBytesIns_Inst_Sbox_11_M38), .Z0_f (new_AGEMA_signal_10199), .Z1_t (new_AGEMA_signal_10200), .Z1_f (new_AGEMA_signal_10201) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M23), .A0_f (new_AGEMA_signal_9356), .A1_t (new_AGEMA_signal_9357), .A1_f (new_AGEMA_signal_9358), .B0_t (SubBytesIns_Inst_Sbox_11_M30), .B0_f (new_AGEMA_signal_9944), .B1_t (new_AGEMA_signal_9945), .B1_f (new_AGEMA_signal_9946), .Z0_t (SubBytesIns_Inst_Sbox_11_M39), .Z0_f (new_AGEMA_signal_10202), .Z1_t (new_AGEMA_signal_10203), .Z1_f (new_AGEMA_signal_10204) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M35), .A0_f (new_AGEMA_signal_9950), .A1_t (new_AGEMA_signal_9951), .A1_f (new_AGEMA_signal_9952), .B0_t (SubBytesIns_Inst_Sbox_11_M36), .B0_f (new_AGEMA_signal_9953), .B1_t (new_AGEMA_signal_9954), .B1_f (new_AGEMA_signal_9955), .Z0_t (SubBytesIns_Inst_Sbox_11_M40), .Z0_f (new_AGEMA_signal_10205), .Z1_t (new_AGEMA_signal_10206), .Z1_f (new_AGEMA_signal_10207) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M38), .A0_f (new_AGEMA_signal_10199), .A1_t (new_AGEMA_signal_10200), .A1_f (new_AGEMA_signal_10201), .B0_t (SubBytesIns_Inst_Sbox_11_M40), .B0_f (new_AGEMA_signal_10205), .B1_t (new_AGEMA_signal_10206), .B1_f (new_AGEMA_signal_10207), .Z0_t (SubBytesIns_Inst_Sbox_11_M41), .Z0_f (new_AGEMA_signal_10796), .Z1_t (new_AGEMA_signal_10797), .Z1_f (new_AGEMA_signal_10798) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M37), .A0_f (new_AGEMA_signal_10196), .A1_t (new_AGEMA_signal_10197), .A1_f (new_AGEMA_signal_10198), .B0_t (SubBytesIns_Inst_Sbox_11_M39), .B0_f (new_AGEMA_signal_10202), .B1_t (new_AGEMA_signal_10203), .B1_f (new_AGEMA_signal_10204), .Z0_t (SubBytesIns_Inst_Sbox_11_M42), .Z0_f (new_AGEMA_signal_10799), .Z1_t (new_AGEMA_signal_10800), .Z1_f (new_AGEMA_signal_10801) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M37), .A0_f (new_AGEMA_signal_10196), .A1_t (new_AGEMA_signal_10197), .A1_f (new_AGEMA_signal_10198), .B0_t (SubBytesIns_Inst_Sbox_11_M38), .B0_f (new_AGEMA_signal_10199), .B1_t (new_AGEMA_signal_10200), .B1_f (new_AGEMA_signal_10201), .Z0_t (SubBytesIns_Inst_Sbox_11_M43), .Z0_f (new_AGEMA_signal_10802), .Z1_t (new_AGEMA_signal_10803), .Z1_f (new_AGEMA_signal_10804) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M39), .A0_f (new_AGEMA_signal_10202), .A1_t (new_AGEMA_signal_10203), .A1_f (new_AGEMA_signal_10204), .B0_t (SubBytesIns_Inst_Sbox_11_M40), .B0_f (new_AGEMA_signal_10205), .B1_t (new_AGEMA_signal_10206), .B1_f (new_AGEMA_signal_10207), .Z0_t (SubBytesIns_Inst_Sbox_11_M44), .Z0_f (new_AGEMA_signal_10805), .Z1_t (new_AGEMA_signal_10806), .Z1_f (new_AGEMA_signal_10807) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M42), .A0_f (new_AGEMA_signal_10799), .A1_t (new_AGEMA_signal_10800), .A1_f (new_AGEMA_signal_10801), .B0_t (SubBytesIns_Inst_Sbox_11_M41), .B0_f (new_AGEMA_signal_10796), .B1_t (new_AGEMA_signal_10797), .B1_f (new_AGEMA_signal_10798), .Z0_t (SubBytesIns_Inst_Sbox_11_M45), .Z0_f (new_AGEMA_signal_11516), .Z1_t (new_AGEMA_signal_11517), .Z1_f (new_AGEMA_signal_11518) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M44), .A0_f (new_AGEMA_signal_10805), .A1_t (new_AGEMA_signal_10806), .A1_f (new_AGEMA_signal_10807), .B0_t (SubBytesIns_Inst_Sbox_11_T6), .B0_f (new_AGEMA_signal_7192), .B1_t (new_AGEMA_signal_7193), .B1_f (new_AGEMA_signal_7194), .Z0_t (SubBytesIns_Inst_Sbox_11_M46), .Z0_f (new_AGEMA_signal_11519), .Z1_t (new_AGEMA_signal_11520), .Z1_f (new_AGEMA_signal_11521) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M40), .A0_f (new_AGEMA_signal_10205), .A1_t (new_AGEMA_signal_10206), .A1_f (new_AGEMA_signal_10207), .B0_t (SubBytesIns_Inst_Sbox_11_T8), .B0_f (new_AGEMA_signal_7901), .B1_t (new_AGEMA_signal_7902), .B1_f (new_AGEMA_signal_7903), .Z0_t (SubBytesIns_Inst_Sbox_11_M47), .Z0_f (new_AGEMA_signal_10808), .Z1_t (new_AGEMA_signal_10809), .Z1_f (new_AGEMA_signal_10810) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M39), .A0_f (new_AGEMA_signal_10202), .A1_t (new_AGEMA_signal_10203), .A1_f (new_AGEMA_signal_10204), .B0_t (ciphertext_s0_t[88]), .B0_f (ciphertext_s0_f[88]), .B1_t (ciphertext_s1_t[88]), .B1_f (ciphertext_s1_f[88]), .Z0_t (SubBytesIns_Inst_Sbox_11_M48), .Z0_f (new_AGEMA_signal_10811), .Z1_t (new_AGEMA_signal_10812), .Z1_f (new_AGEMA_signal_10813) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M43), .A0_f (new_AGEMA_signal_10802), .A1_t (new_AGEMA_signal_10803), .A1_f (new_AGEMA_signal_10804), .B0_t (SubBytesIns_Inst_Sbox_11_T16), .B0_f (new_AGEMA_signal_7204), .B1_t (new_AGEMA_signal_7205), .B1_f (new_AGEMA_signal_7206), .Z0_t (SubBytesIns_Inst_Sbox_11_M49), .Z0_f (new_AGEMA_signal_11522), .Z1_t (new_AGEMA_signal_11523), .Z1_f (new_AGEMA_signal_11524) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M38), .A0_f (new_AGEMA_signal_10199), .A1_t (new_AGEMA_signal_10200), .A1_f (new_AGEMA_signal_10201), .B0_t (SubBytesIns_Inst_Sbox_11_T9), .B0_f (new_AGEMA_signal_7195), .B1_t (new_AGEMA_signal_7196), .B1_f (new_AGEMA_signal_7197), .Z0_t (SubBytesIns_Inst_Sbox_11_M50), .Z0_f (new_AGEMA_signal_10814), .Z1_t (new_AGEMA_signal_10815), .Z1_f (new_AGEMA_signal_10816) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M37), .A0_f (new_AGEMA_signal_10196), .A1_t (new_AGEMA_signal_10197), .A1_f (new_AGEMA_signal_10198), .B0_t (SubBytesIns_Inst_Sbox_11_T17), .B0_f (new_AGEMA_signal_7910), .B1_t (new_AGEMA_signal_7911), .B1_f (new_AGEMA_signal_7912), .Z0_t (SubBytesIns_Inst_Sbox_11_M51), .Z0_f (new_AGEMA_signal_10817), .Z1_t (new_AGEMA_signal_10818), .Z1_f (new_AGEMA_signal_10819) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M42), .A0_f (new_AGEMA_signal_10799), .A1_t (new_AGEMA_signal_10800), .A1_f (new_AGEMA_signal_10801), .B0_t (SubBytesIns_Inst_Sbox_11_T15), .B0_f (new_AGEMA_signal_7201), .B1_t (new_AGEMA_signal_7202), .B1_f (new_AGEMA_signal_7203), .Z0_t (SubBytesIns_Inst_Sbox_11_M52), .Z0_f (new_AGEMA_signal_11525), .Z1_t (new_AGEMA_signal_11526), .Z1_f (new_AGEMA_signal_11527) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M45), .A0_f (new_AGEMA_signal_11516), .A1_t (new_AGEMA_signal_11517), .A1_f (new_AGEMA_signal_11518), .B0_t (SubBytesIns_Inst_Sbox_11_T27), .B0_f (new_AGEMA_signal_7213), .B1_t (new_AGEMA_signal_7214), .B1_f (new_AGEMA_signal_7215), .Z0_t (SubBytesIns_Inst_Sbox_11_M53), .Z0_f (new_AGEMA_signal_12146), .Z1_t (new_AGEMA_signal_12147), .Z1_f (new_AGEMA_signal_12148) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M41), .A0_f (new_AGEMA_signal_10796), .A1_t (new_AGEMA_signal_10797), .A1_f (new_AGEMA_signal_10798), .B0_t (SubBytesIns_Inst_Sbox_11_T10), .B0_f (new_AGEMA_signal_7904), .B1_t (new_AGEMA_signal_7905), .B1_f (new_AGEMA_signal_7906), .Z0_t (SubBytesIns_Inst_Sbox_11_M54), .Z0_f (new_AGEMA_signal_11528), .Z1_t (new_AGEMA_signal_11529), .Z1_f (new_AGEMA_signal_11530) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M44), .A0_f (new_AGEMA_signal_10805), .A1_t (new_AGEMA_signal_10806), .A1_f (new_AGEMA_signal_10807), .B0_t (SubBytesIns_Inst_Sbox_11_T13), .B0_f (new_AGEMA_signal_7198), .B1_t (new_AGEMA_signal_7199), .B1_f (new_AGEMA_signal_7200), .Z0_t (SubBytesIns_Inst_Sbox_11_M55), .Z0_f (new_AGEMA_signal_11531), .Z1_t (new_AGEMA_signal_11532), .Z1_f (new_AGEMA_signal_11533) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M40), .A0_f (new_AGEMA_signal_10205), .A1_t (new_AGEMA_signal_10206), .A1_f (new_AGEMA_signal_10207), .B0_t (SubBytesIns_Inst_Sbox_11_T23), .B0_f (new_AGEMA_signal_7916), .B1_t (new_AGEMA_signal_7917), .B1_f (new_AGEMA_signal_7918), .Z0_t (SubBytesIns_Inst_Sbox_11_M56), .Z0_f (new_AGEMA_signal_10820), .Z1_t (new_AGEMA_signal_10821), .Z1_f (new_AGEMA_signal_10822) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M39), .A0_f (new_AGEMA_signal_10202), .A1_t (new_AGEMA_signal_10203), .A1_f (new_AGEMA_signal_10204), .B0_t (SubBytesIns_Inst_Sbox_11_T19), .B0_f (new_AGEMA_signal_7207), .B1_t (new_AGEMA_signal_7208), .B1_f (new_AGEMA_signal_7209), .Z0_t (SubBytesIns_Inst_Sbox_11_M57), .Z0_f (new_AGEMA_signal_10823), .Z1_t (new_AGEMA_signal_10824), .Z1_f (new_AGEMA_signal_10825) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M43), .A0_f (new_AGEMA_signal_10802), .A1_t (new_AGEMA_signal_10803), .A1_f (new_AGEMA_signal_10804), .B0_t (SubBytesIns_Inst_Sbox_11_T3), .B0_f (new_AGEMA_signal_6682), .B1_t (new_AGEMA_signal_6683), .B1_f (new_AGEMA_signal_6684), .Z0_t (SubBytesIns_Inst_Sbox_11_M58), .Z0_f (new_AGEMA_signal_11534), .Z1_t (new_AGEMA_signal_11535), .Z1_f (new_AGEMA_signal_11536) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M38), .A0_f (new_AGEMA_signal_10199), .A1_t (new_AGEMA_signal_10200), .A1_f (new_AGEMA_signal_10201), .B0_t (SubBytesIns_Inst_Sbox_11_T22), .B0_f (new_AGEMA_signal_7210), .B1_t (new_AGEMA_signal_7211), .B1_f (new_AGEMA_signal_7212), .Z0_t (SubBytesIns_Inst_Sbox_11_M59), .Z0_f (new_AGEMA_signal_10826), .Z1_t (new_AGEMA_signal_10827), .Z1_f (new_AGEMA_signal_10828) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M37), .A0_f (new_AGEMA_signal_10196), .A1_t (new_AGEMA_signal_10197), .A1_f (new_AGEMA_signal_10198), .B0_t (SubBytesIns_Inst_Sbox_11_T20), .B0_f (new_AGEMA_signal_7913), .B1_t (new_AGEMA_signal_7914), .B1_f (new_AGEMA_signal_7915), .Z0_t (SubBytesIns_Inst_Sbox_11_M60), .Z0_f (new_AGEMA_signal_10829), .Z1_t (new_AGEMA_signal_10830), .Z1_f (new_AGEMA_signal_10831) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M42), .A0_f (new_AGEMA_signal_10799), .A1_t (new_AGEMA_signal_10800), .A1_f (new_AGEMA_signal_10801), .B0_t (SubBytesIns_Inst_Sbox_11_T1), .B0_f (new_AGEMA_signal_6676), .B1_t (new_AGEMA_signal_6677), .B1_f (new_AGEMA_signal_6678), .Z0_t (SubBytesIns_Inst_Sbox_11_M61), .Z0_f (new_AGEMA_signal_11537), .Z1_t (new_AGEMA_signal_11538), .Z1_f (new_AGEMA_signal_11539) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M45), .A0_f (new_AGEMA_signal_11516), .A1_t (new_AGEMA_signal_11517), .A1_f (new_AGEMA_signal_11518), .B0_t (SubBytesIns_Inst_Sbox_11_T4), .B0_f (new_AGEMA_signal_6685), .B1_t (new_AGEMA_signal_6686), .B1_f (new_AGEMA_signal_6687), .Z0_t (SubBytesIns_Inst_Sbox_11_M62), .Z0_f (new_AGEMA_signal_12149), .Z1_t (new_AGEMA_signal_12150), .Z1_f (new_AGEMA_signal_12151) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M41), .A0_f (new_AGEMA_signal_10796), .A1_t (new_AGEMA_signal_10797), .A1_f (new_AGEMA_signal_10798), .B0_t (SubBytesIns_Inst_Sbox_11_T2), .B0_f (new_AGEMA_signal_6679), .B1_t (new_AGEMA_signal_6680), .B1_f (new_AGEMA_signal_6681), .Z0_t (SubBytesIns_Inst_Sbox_11_M63), .Z0_f (new_AGEMA_signal_11540), .Z1_t (new_AGEMA_signal_11541), .Z1_f (new_AGEMA_signal_11542) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M61), .A0_f (new_AGEMA_signal_11537), .A1_t (new_AGEMA_signal_11538), .A1_f (new_AGEMA_signal_11539), .B0_t (SubBytesIns_Inst_Sbox_11_M62), .B0_f (new_AGEMA_signal_12149), .B1_t (new_AGEMA_signal_12150), .B1_f (new_AGEMA_signal_12151), .Z0_t (SubBytesIns_Inst_Sbox_11_L0), .Z0_f (new_AGEMA_signal_12701), .Z1_t (new_AGEMA_signal_12702), .Z1_f (new_AGEMA_signal_12703) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M50), .A0_f (new_AGEMA_signal_10814), .A1_t (new_AGEMA_signal_10815), .A1_f (new_AGEMA_signal_10816), .B0_t (SubBytesIns_Inst_Sbox_11_M56), .B0_f (new_AGEMA_signal_10820), .B1_t (new_AGEMA_signal_10821), .B1_f (new_AGEMA_signal_10822), .Z0_t (SubBytesIns_Inst_Sbox_11_L1), .Z0_f (new_AGEMA_signal_11543), .Z1_t (new_AGEMA_signal_11544), .Z1_f (new_AGEMA_signal_11545) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M46), .A0_f (new_AGEMA_signal_11519), .A1_t (new_AGEMA_signal_11520), .A1_f (new_AGEMA_signal_11521), .B0_t (SubBytesIns_Inst_Sbox_11_M48), .B0_f (new_AGEMA_signal_10811), .B1_t (new_AGEMA_signal_10812), .B1_f (new_AGEMA_signal_10813), .Z0_t (SubBytesIns_Inst_Sbox_11_L2), .Z0_f (new_AGEMA_signal_12152), .Z1_t (new_AGEMA_signal_12153), .Z1_f (new_AGEMA_signal_12154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M47), .A0_f (new_AGEMA_signal_10808), .A1_t (new_AGEMA_signal_10809), .A1_f (new_AGEMA_signal_10810), .B0_t (SubBytesIns_Inst_Sbox_11_M55), .B0_f (new_AGEMA_signal_11531), .B1_t (new_AGEMA_signal_11532), .B1_f (new_AGEMA_signal_11533), .Z0_t (SubBytesIns_Inst_Sbox_11_L3), .Z0_f (new_AGEMA_signal_12155), .Z1_t (new_AGEMA_signal_12156), .Z1_f (new_AGEMA_signal_12157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M54), .A0_f (new_AGEMA_signal_11528), .A1_t (new_AGEMA_signal_11529), .A1_f (new_AGEMA_signal_11530), .B0_t (SubBytesIns_Inst_Sbox_11_M58), .B0_f (new_AGEMA_signal_11534), .B1_t (new_AGEMA_signal_11535), .B1_f (new_AGEMA_signal_11536), .Z0_t (SubBytesIns_Inst_Sbox_11_L4), .Z0_f (new_AGEMA_signal_12158), .Z1_t (new_AGEMA_signal_12159), .Z1_f (new_AGEMA_signal_12160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M49), .A0_f (new_AGEMA_signal_11522), .A1_t (new_AGEMA_signal_11523), .A1_f (new_AGEMA_signal_11524), .B0_t (SubBytesIns_Inst_Sbox_11_M61), .B0_f (new_AGEMA_signal_11537), .B1_t (new_AGEMA_signal_11538), .B1_f (new_AGEMA_signal_11539), .Z0_t (SubBytesIns_Inst_Sbox_11_L5), .Z0_f (new_AGEMA_signal_12161), .Z1_t (new_AGEMA_signal_12162), .Z1_f (new_AGEMA_signal_12163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M62), .A0_f (new_AGEMA_signal_12149), .A1_t (new_AGEMA_signal_12150), .A1_f (new_AGEMA_signal_12151), .B0_t (SubBytesIns_Inst_Sbox_11_L5), .B0_f (new_AGEMA_signal_12161), .B1_t (new_AGEMA_signal_12162), .B1_f (new_AGEMA_signal_12163), .Z0_t (SubBytesIns_Inst_Sbox_11_L6), .Z0_f (new_AGEMA_signal_12704), .Z1_t (new_AGEMA_signal_12705), .Z1_f (new_AGEMA_signal_12706) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M46), .A0_f (new_AGEMA_signal_11519), .A1_t (new_AGEMA_signal_11520), .A1_f (new_AGEMA_signal_11521), .B0_t (SubBytesIns_Inst_Sbox_11_L3), .B0_f (new_AGEMA_signal_12155), .B1_t (new_AGEMA_signal_12156), .B1_f (new_AGEMA_signal_12157), .Z0_t (SubBytesIns_Inst_Sbox_11_L7), .Z0_f (new_AGEMA_signal_12707), .Z1_t (new_AGEMA_signal_12708), .Z1_f (new_AGEMA_signal_12709) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M51), .A0_f (new_AGEMA_signal_10817), .A1_t (new_AGEMA_signal_10818), .A1_f (new_AGEMA_signal_10819), .B0_t (SubBytesIns_Inst_Sbox_11_M59), .B0_f (new_AGEMA_signal_10826), .B1_t (new_AGEMA_signal_10827), .B1_f (new_AGEMA_signal_10828), .Z0_t (SubBytesIns_Inst_Sbox_11_L8), .Z0_f (new_AGEMA_signal_11546), .Z1_t (new_AGEMA_signal_11547), .Z1_f (new_AGEMA_signal_11548) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M52), .A0_f (new_AGEMA_signal_11525), .A1_t (new_AGEMA_signal_11526), .A1_f (new_AGEMA_signal_11527), .B0_t (SubBytesIns_Inst_Sbox_11_M53), .B0_f (new_AGEMA_signal_12146), .B1_t (new_AGEMA_signal_12147), .B1_f (new_AGEMA_signal_12148), .Z0_t (SubBytesIns_Inst_Sbox_11_L9), .Z0_f (new_AGEMA_signal_12710), .Z1_t (new_AGEMA_signal_12711), .Z1_f (new_AGEMA_signal_12712) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M53), .A0_f (new_AGEMA_signal_12146), .A1_t (new_AGEMA_signal_12147), .A1_f (new_AGEMA_signal_12148), .B0_t (SubBytesIns_Inst_Sbox_11_L4), .B0_f (new_AGEMA_signal_12158), .B1_t (new_AGEMA_signal_12159), .B1_f (new_AGEMA_signal_12160), .Z0_t (SubBytesIns_Inst_Sbox_11_L10), .Z0_f (new_AGEMA_signal_12713), .Z1_t (new_AGEMA_signal_12714), .Z1_f (new_AGEMA_signal_12715) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M60), .A0_f (new_AGEMA_signal_10829), .A1_t (new_AGEMA_signal_10830), .A1_f (new_AGEMA_signal_10831), .B0_t (SubBytesIns_Inst_Sbox_11_L2), .B0_f (new_AGEMA_signal_12152), .B1_t (new_AGEMA_signal_12153), .B1_f (new_AGEMA_signal_12154), .Z0_t (SubBytesIns_Inst_Sbox_11_L11), .Z0_f (new_AGEMA_signal_12716), .Z1_t (new_AGEMA_signal_12717), .Z1_f (new_AGEMA_signal_12718) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M48), .A0_f (new_AGEMA_signal_10811), .A1_t (new_AGEMA_signal_10812), .A1_f (new_AGEMA_signal_10813), .B0_t (SubBytesIns_Inst_Sbox_11_M51), .B0_f (new_AGEMA_signal_10817), .B1_t (new_AGEMA_signal_10818), .B1_f (new_AGEMA_signal_10819), .Z0_t (SubBytesIns_Inst_Sbox_11_L12), .Z0_f (new_AGEMA_signal_11549), .Z1_t (new_AGEMA_signal_11550), .Z1_f (new_AGEMA_signal_11551) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M50), .A0_f (new_AGEMA_signal_10814), .A1_t (new_AGEMA_signal_10815), .A1_f (new_AGEMA_signal_10816), .B0_t (SubBytesIns_Inst_Sbox_11_L0), .B0_f (new_AGEMA_signal_12701), .B1_t (new_AGEMA_signal_12702), .B1_f (new_AGEMA_signal_12703), .Z0_t (SubBytesIns_Inst_Sbox_11_L13), .Z0_f (new_AGEMA_signal_13331), .Z1_t (new_AGEMA_signal_13332), .Z1_f (new_AGEMA_signal_13333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M52), .A0_f (new_AGEMA_signal_11525), .A1_t (new_AGEMA_signal_11526), .A1_f (new_AGEMA_signal_11527), .B0_t (SubBytesIns_Inst_Sbox_11_M61), .B0_f (new_AGEMA_signal_11537), .B1_t (new_AGEMA_signal_11538), .B1_f (new_AGEMA_signal_11539), .Z0_t (SubBytesIns_Inst_Sbox_11_L14), .Z0_f (new_AGEMA_signal_12164), .Z1_t (new_AGEMA_signal_12165), .Z1_f (new_AGEMA_signal_12166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M55), .A0_f (new_AGEMA_signal_11531), .A1_t (new_AGEMA_signal_11532), .A1_f (new_AGEMA_signal_11533), .B0_t (SubBytesIns_Inst_Sbox_11_L1), .B0_f (new_AGEMA_signal_11543), .B1_t (new_AGEMA_signal_11544), .B1_f (new_AGEMA_signal_11545), .Z0_t (SubBytesIns_Inst_Sbox_11_L15), .Z0_f (new_AGEMA_signal_12167), .Z1_t (new_AGEMA_signal_12168), .Z1_f (new_AGEMA_signal_12169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M56), .A0_f (new_AGEMA_signal_10820), .A1_t (new_AGEMA_signal_10821), .A1_f (new_AGEMA_signal_10822), .B0_t (SubBytesIns_Inst_Sbox_11_L0), .B0_f (new_AGEMA_signal_12701), .B1_t (new_AGEMA_signal_12702), .B1_f (new_AGEMA_signal_12703), .Z0_t (SubBytesIns_Inst_Sbox_11_L16), .Z0_f (new_AGEMA_signal_13334), .Z1_t (new_AGEMA_signal_13335), .Z1_f (new_AGEMA_signal_13336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M57), .A0_f (new_AGEMA_signal_10823), .A1_t (new_AGEMA_signal_10824), .A1_f (new_AGEMA_signal_10825), .B0_t (SubBytesIns_Inst_Sbox_11_L1), .B0_f (new_AGEMA_signal_11543), .B1_t (new_AGEMA_signal_11544), .B1_f (new_AGEMA_signal_11545), .Z0_t (SubBytesIns_Inst_Sbox_11_L17), .Z0_f (new_AGEMA_signal_12170), .Z1_t (new_AGEMA_signal_12171), .Z1_f (new_AGEMA_signal_12172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M58), .A0_f (new_AGEMA_signal_11534), .A1_t (new_AGEMA_signal_11535), .A1_f (new_AGEMA_signal_11536), .B0_t (SubBytesIns_Inst_Sbox_11_L8), .B0_f (new_AGEMA_signal_11546), .B1_t (new_AGEMA_signal_11547), .B1_f (new_AGEMA_signal_11548), .Z0_t (SubBytesIns_Inst_Sbox_11_L18), .Z0_f (new_AGEMA_signal_12173), .Z1_t (new_AGEMA_signal_12174), .Z1_f (new_AGEMA_signal_12175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M63), .A0_f (new_AGEMA_signal_11540), .A1_t (new_AGEMA_signal_11541), .A1_f (new_AGEMA_signal_11542), .B0_t (SubBytesIns_Inst_Sbox_11_L4), .B0_f (new_AGEMA_signal_12158), .B1_t (new_AGEMA_signal_12159), .B1_f (new_AGEMA_signal_12160), .Z0_t (SubBytesIns_Inst_Sbox_11_L19), .Z0_f (new_AGEMA_signal_12719), .Z1_t (new_AGEMA_signal_12720), .Z1_f (new_AGEMA_signal_12721) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L0), .A0_f (new_AGEMA_signal_12701), .A1_t (new_AGEMA_signal_12702), .A1_f (new_AGEMA_signal_12703), .B0_t (SubBytesIns_Inst_Sbox_11_L1), .B0_f (new_AGEMA_signal_11543), .B1_t (new_AGEMA_signal_11544), .B1_f (new_AGEMA_signal_11545), .Z0_t (SubBytesIns_Inst_Sbox_11_L20), .Z0_f (new_AGEMA_signal_13337), .Z1_t (new_AGEMA_signal_13338), .Z1_f (new_AGEMA_signal_13339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L1), .A0_f (new_AGEMA_signal_11543), .A1_t (new_AGEMA_signal_11544), .A1_f (new_AGEMA_signal_11545), .B0_t (SubBytesIns_Inst_Sbox_11_L7), .B0_f (new_AGEMA_signal_12707), .B1_t (new_AGEMA_signal_12708), .B1_f (new_AGEMA_signal_12709), .Z0_t (SubBytesIns_Inst_Sbox_11_L21), .Z0_f (new_AGEMA_signal_13340), .Z1_t (new_AGEMA_signal_13341), .Z1_f (new_AGEMA_signal_13342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L3), .A0_f (new_AGEMA_signal_12155), .A1_t (new_AGEMA_signal_12156), .A1_f (new_AGEMA_signal_12157), .B0_t (SubBytesIns_Inst_Sbox_11_L12), .B0_f (new_AGEMA_signal_11549), .B1_t (new_AGEMA_signal_11550), .B1_f (new_AGEMA_signal_11551), .Z0_t (SubBytesIns_Inst_Sbox_11_L22), .Z0_f (new_AGEMA_signal_12722), .Z1_t (new_AGEMA_signal_12723), .Z1_f (new_AGEMA_signal_12724) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L18), .A0_f (new_AGEMA_signal_12173), .A1_t (new_AGEMA_signal_12174), .A1_f (new_AGEMA_signal_12175), .B0_t (SubBytesIns_Inst_Sbox_11_L2), .B0_f (new_AGEMA_signal_12152), .B1_t (new_AGEMA_signal_12153), .B1_f (new_AGEMA_signal_12154), .Z0_t (SubBytesIns_Inst_Sbox_11_L23), .Z0_f (new_AGEMA_signal_12725), .Z1_t (new_AGEMA_signal_12726), .Z1_f (new_AGEMA_signal_12727) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L15), .A0_f (new_AGEMA_signal_12167), .A1_t (new_AGEMA_signal_12168), .A1_f (new_AGEMA_signal_12169), .B0_t (SubBytesIns_Inst_Sbox_11_L9), .B0_f (new_AGEMA_signal_12710), .B1_t (new_AGEMA_signal_12711), .B1_f (new_AGEMA_signal_12712), .Z0_t (SubBytesIns_Inst_Sbox_11_L24), .Z0_f (new_AGEMA_signal_13343), .Z1_t (new_AGEMA_signal_13344), .Z1_f (new_AGEMA_signal_13345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L6), .A0_f (new_AGEMA_signal_12704), .A1_t (new_AGEMA_signal_12705), .A1_f (new_AGEMA_signal_12706), .B0_t (SubBytesIns_Inst_Sbox_11_L10), .B0_f (new_AGEMA_signal_12713), .B1_t (new_AGEMA_signal_12714), .B1_f (new_AGEMA_signal_12715), .Z0_t (SubBytesIns_Inst_Sbox_11_L25), .Z0_f (new_AGEMA_signal_13346), .Z1_t (new_AGEMA_signal_13347), .Z1_f (new_AGEMA_signal_13348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L7), .A0_f (new_AGEMA_signal_12707), .A1_t (new_AGEMA_signal_12708), .A1_f (new_AGEMA_signal_12709), .B0_t (SubBytesIns_Inst_Sbox_11_L9), .B0_f (new_AGEMA_signal_12710), .B1_t (new_AGEMA_signal_12711), .B1_f (new_AGEMA_signal_12712), .Z0_t (SubBytesIns_Inst_Sbox_11_L26), .Z0_f (new_AGEMA_signal_13349), .Z1_t (new_AGEMA_signal_13350), .Z1_f (new_AGEMA_signal_13351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L8), .A0_f (new_AGEMA_signal_11546), .A1_t (new_AGEMA_signal_11547), .A1_f (new_AGEMA_signal_11548), .B0_t (SubBytesIns_Inst_Sbox_11_L10), .B0_f (new_AGEMA_signal_12713), .B1_t (new_AGEMA_signal_12714), .B1_f (new_AGEMA_signal_12715), .Z0_t (SubBytesIns_Inst_Sbox_11_L27), .Z0_f (new_AGEMA_signal_13352), .Z1_t (new_AGEMA_signal_13353), .Z1_f (new_AGEMA_signal_13354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L11), .A0_f (new_AGEMA_signal_12716), .A1_t (new_AGEMA_signal_12717), .A1_f (new_AGEMA_signal_12718), .B0_t (SubBytesIns_Inst_Sbox_11_L14), .B0_f (new_AGEMA_signal_12164), .B1_t (new_AGEMA_signal_12165), .B1_f (new_AGEMA_signal_12166), .Z0_t (SubBytesIns_Inst_Sbox_11_L28), .Z0_f (new_AGEMA_signal_13355), .Z1_t (new_AGEMA_signal_13356), .Z1_f (new_AGEMA_signal_13357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L11), .A0_f (new_AGEMA_signal_12716), .A1_t (new_AGEMA_signal_12717), .A1_f (new_AGEMA_signal_12718), .B0_t (SubBytesIns_Inst_Sbox_11_L17), .B0_f (new_AGEMA_signal_12170), .B1_t (new_AGEMA_signal_12171), .B1_f (new_AGEMA_signal_12172), .Z0_t (SubBytesIns_Inst_Sbox_11_L29), .Z0_f (new_AGEMA_signal_13358), .Z1_t (new_AGEMA_signal_13359), .Z1_f (new_AGEMA_signal_13360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L6), .A0_f (new_AGEMA_signal_12704), .A1_t (new_AGEMA_signal_12705), .A1_f (new_AGEMA_signal_12706), .B0_t (SubBytesIns_Inst_Sbox_11_L24), .B0_f (new_AGEMA_signal_13343), .B1_t (new_AGEMA_signal_13344), .B1_f (new_AGEMA_signal_13345), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .Z0_f (new_AGEMA_signal_13871), .Z1_t (new_AGEMA_signal_13872), .Z1_f (new_AGEMA_signal_13873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L16), .A0_f (new_AGEMA_signal_13334), .A1_t (new_AGEMA_signal_13335), .A1_f (new_AGEMA_signal_13336), .B0_t (SubBytesIns_Inst_Sbox_11_L26), .B0_f (new_AGEMA_signal_13349), .B1_t (new_AGEMA_signal_13350), .B1_f (new_AGEMA_signal_13351), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .Z0_f (new_AGEMA_signal_13874), .Z1_t (new_AGEMA_signal_13875), .Z1_f (new_AGEMA_signal_13876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L19), .A0_f (new_AGEMA_signal_12719), .A1_t (new_AGEMA_signal_12720), .A1_f (new_AGEMA_signal_12721), .B0_t (SubBytesIns_Inst_Sbox_11_L28), .B0_f (new_AGEMA_signal_13355), .B1_t (new_AGEMA_signal_13356), .B1_f (new_AGEMA_signal_13357), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .Z0_f (new_AGEMA_signal_13877), .Z1_t (new_AGEMA_signal_13878), .Z1_f (new_AGEMA_signal_13879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L6), .A0_f (new_AGEMA_signal_12704), .A1_t (new_AGEMA_signal_12705), .A1_f (new_AGEMA_signal_12706), .B0_t (SubBytesIns_Inst_Sbox_11_L21), .B0_f (new_AGEMA_signal_13340), .B1_t (new_AGEMA_signal_13341), .B1_f (new_AGEMA_signal_13342), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .Z0_f (new_AGEMA_signal_13880), .Z1_t (new_AGEMA_signal_13881), .Z1_f (new_AGEMA_signal_13882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L20), .A0_f (new_AGEMA_signal_13337), .A1_t (new_AGEMA_signal_13338), .A1_f (new_AGEMA_signal_13339), .B0_t (SubBytesIns_Inst_Sbox_11_L22), .B0_f (new_AGEMA_signal_12722), .B1_t (new_AGEMA_signal_12723), .B1_f (new_AGEMA_signal_12724), .Z0_t (MixColumnsInput[91]), .Z0_f (new_AGEMA_signal_13883), .Z1_t (new_AGEMA_signal_13884), .Z1_f (new_AGEMA_signal_13885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L25), .A0_f (new_AGEMA_signal_13346), .A1_t (new_AGEMA_signal_13347), .A1_f (new_AGEMA_signal_13348), .B0_t (SubBytesIns_Inst_Sbox_11_L29), .B0_f (new_AGEMA_signal_13358), .B1_t (new_AGEMA_signal_13359), .B1_f (new_AGEMA_signal_13360), .Z0_t (MixColumnsInput[90]), .Z0_f (new_AGEMA_signal_13886), .Z1_t (new_AGEMA_signal_13887), .Z1_f (new_AGEMA_signal_13888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L13), .A0_f (new_AGEMA_signal_13331), .A1_t (new_AGEMA_signal_13332), .A1_f (new_AGEMA_signal_13333), .B0_t (SubBytesIns_Inst_Sbox_11_L27), .B0_f (new_AGEMA_signal_13352), .B1_t (new_AGEMA_signal_13353), .B1_f (new_AGEMA_signal_13354), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .Z0_f (new_AGEMA_signal_13889), .Z1_t (new_AGEMA_signal_13890), .Z1_f (new_AGEMA_signal_13891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L6), .A0_f (new_AGEMA_signal_12704), .A1_t (new_AGEMA_signal_12705), .A1_f (new_AGEMA_signal_12706), .B0_t (SubBytesIns_Inst_Sbox_11_L23), .B0_f (new_AGEMA_signal_12725), .B1_t (new_AGEMA_signal_12726), .B1_f (new_AGEMA_signal_12727), .Z0_t (MixColumnsInput[88]), .Z0_f (new_AGEMA_signal_13361), .Z1_t (new_AGEMA_signal_13362), .Z1_f (new_AGEMA_signal_13363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (ciphertext_s0_t[100]), .B0_f (ciphertext_s0_f[100]), .B1_t (ciphertext_s1_t[100]), .B1_f (ciphertext_s1_f[100]), .Z0_t (SubBytesIns_Inst_Sbox_12_T1), .Z0_f (new_AGEMA_signal_6706), .Z1_t (new_AGEMA_signal_6707), .Z1_f (new_AGEMA_signal_6708) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (ciphertext_s0_t[98]), .B0_f (ciphertext_s0_f[98]), .B1_t (ciphertext_s1_t[98]), .B1_f (ciphertext_s1_f[98]), .Z0_t (SubBytesIns_Inst_Sbox_12_T2), .Z0_f (new_AGEMA_signal_6709), .Z1_t (new_AGEMA_signal_6710), .Z1_f (new_AGEMA_signal_6711) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (ciphertext_s0_t[97]), .B0_f (ciphertext_s0_f[97]), .B1_t (ciphertext_s1_t[97]), .B1_f (ciphertext_s1_f[97]), .Z0_t (SubBytesIns_Inst_Sbox_12_T3), .Z0_f (new_AGEMA_signal_6712), .Z1_t (new_AGEMA_signal_6713), .Z1_f (new_AGEMA_signal_6714) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[100]), .A0_f (ciphertext_s0_f[100]), .A1_t (ciphertext_s1_t[100]), .A1_f (ciphertext_s1_f[100]), .B0_t (ciphertext_s0_t[98]), .B0_f (ciphertext_s0_f[98]), .B1_t (ciphertext_s1_t[98]), .B1_f (ciphertext_s1_f[98]), .Z0_t (SubBytesIns_Inst_Sbox_12_T4), .Z0_f (new_AGEMA_signal_6715), .Z1_t (new_AGEMA_signal_6716), .Z1_f (new_AGEMA_signal_6717) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[99]), .A0_f (ciphertext_s0_f[99]), .A1_t (ciphertext_s1_t[99]), .A1_f (ciphertext_s1_f[99]), .B0_t (ciphertext_s0_t[97]), .B0_f (ciphertext_s0_f[97]), .B1_t (ciphertext_s1_t[97]), .B1_f (ciphertext_s1_f[97]), .Z0_t (SubBytesIns_Inst_Sbox_12_T5), .Z0_f (new_AGEMA_signal_6718), .Z1_t (new_AGEMA_signal_6719), .Z1_f (new_AGEMA_signal_6720) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T1), .A0_f (new_AGEMA_signal_6706), .A1_t (new_AGEMA_signal_6707), .A1_f (new_AGEMA_signal_6708), .B0_t (SubBytesIns_Inst_Sbox_12_T5), .B0_f (new_AGEMA_signal_6718), .B1_t (new_AGEMA_signal_6719), .B1_f (new_AGEMA_signal_6720), .Z0_t (SubBytesIns_Inst_Sbox_12_T6), .Z0_f (new_AGEMA_signal_7216), .Z1_t (new_AGEMA_signal_7217), .Z1_f (new_AGEMA_signal_7218) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[102]), .A0_f (ciphertext_s0_f[102]), .A1_t (ciphertext_s1_t[102]), .A1_f (ciphertext_s1_f[102]), .B0_t (ciphertext_s0_t[101]), .B0_f (ciphertext_s0_f[101]), .B1_t (ciphertext_s1_t[101]), .B1_f (ciphertext_s1_f[101]), .Z0_t (SubBytesIns_Inst_Sbox_12_T7), .Z0_f (new_AGEMA_signal_6721), .Z1_t (new_AGEMA_signal_6722), .Z1_f (new_AGEMA_signal_6723) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[96]), .A0_f (ciphertext_s0_f[96]), .A1_t (ciphertext_s1_t[96]), .A1_f (ciphertext_s1_f[96]), .B0_t (SubBytesIns_Inst_Sbox_12_T6), .B0_f (new_AGEMA_signal_7216), .B1_t (new_AGEMA_signal_7217), .B1_f (new_AGEMA_signal_7218), .Z0_t (SubBytesIns_Inst_Sbox_12_T8), .Z0_f (new_AGEMA_signal_7940), .Z1_t (new_AGEMA_signal_7941), .Z1_f (new_AGEMA_signal_7942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[96]), .A0_f (ciphertext_s0_f[96]), .A1_t (ciphertext_s1_t[96]), .A1_f (ciphertext_s1_f[96]), .B0_t (SubBytesIns_Inst_Sbox_12_T7), .B0_f (new_AGEMA_signal_6721), .B1_t (new_AGEMA_signal_6722), .B1_f (new_AGEMA_signal_6723), .Z0_t (SubBytesIns_Inst_Sbox_12_T9), .Z0_f (new_AGEMA_signal_7219), .Z1_t (new_AGEMA_signal_7220), .Z1_f (new_AGEMA_signal_7221) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T6), .A0_f (new_AGEMA_signal_7216), .A1_t (new_AGEMA_signal_7217), .A1_f (new_AGEMA_signal_7218), .B0_t (SubBytesIns_Inst_Sbox_12_T7), .B0_f (new_AGEMA_signal_6721), .B1_t (new_AGEMA_signal_6722), .B1_f (new_AGEMA_signal_6723), .Z0_t (SubBytesIns_Inst_Sbox_12_T10), .Z0_f (new_AGEMA_signal_7943), .Z1_t (new_AGEMA_signal_7944), .Z1_f (new_AGEMA_signal_7945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[102]), .A0_f (ciphertext_s0_f[102]), .A1_t (ciphertext_s1_t[102]), .A1_f (ciphertext_s1_f[102]), .B0_t (ciphertext_s0_t[98]), .B0_f (ciphertext_s0_f[98]), .B1_t (ciphertext_s1_t[98]), .B1_f (ciphertext_s1_f[98]), .Z0_t (SubBytesIns_Inst_Sbox_12_T11), .Z0_f (new_AGEMA_signal_6724), .Z1_t (new_AGEMA_signal_6725), .Z1_f (new_AGEMA_signal_6726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[101]), .A0_f (ciphertext_s0_f[101]), .A1_t (ciphertext_s1_t[101]), .A1_f (ciphertext_s1_f[101]), .B0_t (ciphertext_s0_t[98]), .B0_f (ciphertext_s0_f[98]), .B1_t (ciphertext_s1_t[98]), .B1_f (ciphertext_s1_f[98]), .Z0_t (SubBytesIns_Inst_Sbox_12_T12), .Z0_f (new_AGEMA_signal_6727), .Z1_t (new_AGEMA_signal_6728), .Z1_f (new_AGEMA_signal_6729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T3), .A0_f (new_AGEMA_signal_6712), .A1_t (new_AGEMA_signal_6713), .A1_f (new_AGEMA_signal_6714), .B0_t (SubBytesIns_Inst_Sbox_12_T4), .B0_f (new_AGEMA_signal_6715), .B1_t (new_AGEMA_signal_6716), .B1_f (new_AGEMA_signal_6717), .Z0_t (SubBytesIns_Inst_Sbox_12_T13), .Z0_f (new_AGEMA_signal_7222), .Z1_t (new_AGEMA_signal_7223), .Z1_f (new_AGEMA_signal_7224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T6), .A0_f (new_AGEMA_signal_7216), .A1_t (new_AGEMA_signal_7217), .A1_f (new_AGEMA_signal_7218), .B0_t (SubBytesIns_Inst_Sbox_12_T11), .B0_f (new_AGEMA_signal_6724), .B1_t (new_AGEMA_signal_6725), .B1_f (new_AGEMA_signal_6726), .Z0_t (SubBytesIns_Inst_Sbox_12_T14), .Z0_f (new_AGEMA_signal_7946), .Z1_t (new_AGEMA_signal_7947), .Z1_f (new_AGEMA_signal_7948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T5), .A0_f (new_AGEMA_signal_6718), .A1_t (new_AGEMA_signal_6719), .A1_f (new_AGEMA_signal_6720), .B0_t (SubBytesIns_Inst_Sbox_12_T11), .B0_f (new_AGEMA_signal_6724), .B1_t (new_AGEMA_signal_6725), .B1_f (new_AGEMA_signal_6726), .Z0_t (SubBytesIns_Inst_Sbox_12_T15), .Z0_f (new_AGEMA_signal_7225), .Z1_t (new_AGEMA_signal_7226), .Z1_f (new_AGEMA_signal_7227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T5), .A0_f (new_AGEMA_signal_6718), .A1_t (new_AGEMA_signal_6719), .A1_f (new_AGEMA_signal_6720), .B0_t (SubBytesIns_Inst_Sbox_12_T12), .B0_f (new_AGEMA_signal_6727), .B1_t (new_AGEMA_signal_6728), .B1_f (new_AGEMA_signal_6729), .Z0_t (SubBytesIns_Inst_Sbox_12_T16), .Z0_f (new_AGEMA_signal_7228), .Z1_t (new_AGEMA_signal_7229), .Z1_f (new_AGEMA_signal_7230) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T9), .A0_f (new_AGEMA_signal_7219), .A1_t (new_AGEMA_signal_7220), .A1_f (new_AGEMA_signal_7221), .B0_t (SubBytesIns_Inst_Sbox_12_T16), .B0_f (new_AGEMA_signal_7228), .B1_t (new_AGEMA_signal_7229), .B1_f (new_AGEMA_signal_7230), .Z0_t (SubBytesIns_Inst_Sbox_12_T17), .Z0_f (new_AGEMA_signal_7949), .Z1_t (new_AGEMA_signal_7950), .Z1_f (new_AGEMA_signal_7951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[100]), .A0_f (ciphertext_s0_f[100]), .A1_t (ciphertext_s1_t[100]), .A1_f (ciphertext_s1_f[100]), .B0_t (ciphertext_s0_t[96]), .B0_f (ciphertext_s0_f[96]), .B1_t (ciphertext_s1_t[96]), .B1_f (ciphertext_s1_f[96]), .Z0_t (SubBytesIns_Inst_Sbox_12_T18), .Z0_f (new_AGEMA_signal_6730), .Z1_t (new_AGEMA_signal_6731), .Z1_f (new_AGEMA_signal_6732) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T7), .A0_f (new_AGEMA_signal_6721), .A1_t (new_AGEMA_signal_6722), .A1_f (new_AGEMA_signal_6723), .B0_t (SubBytesIns_Inst_Sbox_12_T18), .B0_f (new_AGEMA_signal_6730), .B1_t (new_AGEMA_signal_6731), .B1_f (new_AGEMA_signal_6732), .Z0_t (SubBytesIns_Inst_Sbox_12_T19), .Z0_f (new_AGEMA_signal_7231), .Z1_t (new_AGEMA_signal_7232), .Z1_f (new_AGEMA_signal_7233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T1), .A0_f (new_AGEMA_signal_6706), .A1_t (new_AGEMA_signal_6707), .A1_f (new_AGEMA_signal_6708), .B0_t (SubBytesIns_Inst_Sbox_12_T19), .B0_f (new_AGEMA_signal_7231), .B1_t (new_AGEMA_signal_7232), .B1_f (new_AGEMA_signal_7233), .Z0_t (SubBytesIns_Inst_Sbox_12_T20), .Z0_f (new_AGEMA_signal_7952), .Z1_t (new_AGEMA_signal_7953), .Z1_f (new_AGEMA_signal_7954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[97]), .A0_f (ciphertext_s0_f[97]), .A1_t (ciphertext_s1_t[97]), .A1_f (ciphertext_s1_f[97]), .B0_t (ciphertext_s0_t[96]), .B0_f (ciphertext_s0_f[96]), .B1_t (ciphertext_s1_t[96]), .B1_f (ciphertext_s1_f[96]), .Z0_t (SubBytesIns_Inst_Sbox_12_T21), .Z0_f (new_AGEMA_signal_6733), .Z1_t (new_AGEMA_signal_6734), .Z1_f (new_AGEMA_signal_6735) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T7), .A0_f (new_AGEMA_signal_6721), .A1_t (new_AGEMA_signal_6722), .A1_f (new_AGEMA_signal_6723), .B0_t (SubBytesIns_Inst_Sbox_12_T21), .B0_f (new_AGEMA_signal_6733), .B1_t (new_AGEMA_signal_6734), .B1_f (new_AGEMA_signal_6735), .Z0_t (SubBytesIns_Inst_Sbox_12_T22), .Z0_f (new_AGEMA_signal_7234), .Z1_t (new_AGEMA_signal_7235), .Z1_f (new_AGEMA_signal_7236) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T2), .A0_f (new_AGEMA_signal_6709), .A1_t (new_AGEMA_signal_6710), .A1_f (new_AGEMA_signal_6711), .B0_t (SubBytesIns_Inst_Sbox_12_T22), .B0_f (new_AGEMA_signal_7234), .B1_t (new_AGEMA_signal_7235), .B1_f (new_AGEMA_signal_7236), .Z0_t (SubBytesIns_Inst_Sbox_12_T23), .Z0_f (new_AGEMA_signal_7955), .Z1_t (new_AGEMA_signal_7956), .Z1_f (new_AGEMA_signal_7957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T2), .A0_f (new_AGEMA_signal_6709), .A1_t (new_AGEMA_signal_6710), .A1_f (new_AGEMA_signal_6711), .B0_t (SubBytesIns_Inst_Sbox_12_T10), .B0_f (new_AGEMA_signal_7943), .B1_t (new_AGEMA_signal_7944), .B1_f (new_AGEMA_signal_7945), .Z0_t (SubBytesIns_Inst_Sbox_12_T24), .Z0_f (new_AGEMA_signal_8528), .Z1_t (new_AGEMA_signal_8529), .Z1_f (new_AGEMA_signal_8530) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T20), .A0_f (new_AGEMA_signal_7952), .A1_t (new_AGEMA_signal_7953), .A1_f (new_AGEMA_signal_7954), .B0_t (SubBytesIns_Inst_Sbox_12_T17), .B0_f (new_AGEMA_signal_7949), .B1_t (new_AGEMA_signal_7950), .B1_f (new_AGEMA_signal_7951), .Z0_t (SubBytesIns_Inst_Sbox_12_T25), .Z0_f (new_AGEMA_signal_8531), .Z1_t (new_AGEMA_signal_8532), .Z1_f (new_AGEMA_signal_8533) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T3), .A0_f (new_AGEMA_signal_6712), .A1_t (new_AGEMA_signal_6713), .A1_f (new_AGEMA_signal_6714), .B0_t (SubBytesIns_Inst_Sbox_12_T16), .B0_f (new_AGEMA_signal_7228), .B1_t (new_AGEMA_signal_7229), .B1_f (new_AGEMA_signal_7230), .Z0_t (SubBytesIns_Inst_Sbox_12_T26), .Z0_f (new_AGEMA_signal_7958), .Z1_t (new_AGEMA_signal_7959), .Z1_f (new_AGEMA_signal_7960) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T1), .A0_f (new_AGEMA_signal_6706), .A1_t (new_AGEMA_signal_6707), .A1_f (new_AGEMA_signal_6708), .B0_t (SubBytesIns_Inst_Sbox_12_T12), .B0_f (new_AGEMA_signal_6727), .B1_t (new_AGEMA_signal_6728), .B1_f (new_AGEMA_signal_6729), .Z0_t (SubBytesIns_Inst_Sbox_12_T27), .Z0_f (new_AGEMA_signal_7237), .Z1_t (new_AGEMA_signal_7238), .Z1_f (new_AGEMA_signal_7239) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T13), .A0_f (new_AGEMA_signal_7222), .A1_t (new_AGEMA_signal_7223), .A1_f (new_AGEMA_signal_7224), .B0_t (SubBytesIns_Inst_Sbox_12_T6), .B0_f (new_AGEMA_signal_7216), .B1_t (new_AGEMA_signal_7217), .B1_f (new_AGEMA_signal_7218), .Z0_t (SubBytesIns_Inst_Sbox_12_M1), .Z0_f (new_AGEMA_signal_7961), .Z1_t (new_AGEMA_signal_7962), .Z1_f (new_AGEMA_signal_7963) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T23), .A0_f (new_AGEMA_signal_7955), .A1_t (new_AGEMA_signal_7956), .A1_f (new_AGEMA_signal_7957), .B0_t (SubBytesIns_Inst_Sbox_12_T8), .B0_f (new_AGEMA_signal_7940), .B1_t (new_AGEMA_signal_7941), .B1_f (new_AGEMA_signal_7942), .Z0_t (SubBytesIns_Inst_Sbox_12_M2), .Z0_f (new_AGEMA_signal_8534), .Z1_t (new_AGEMA_signal_8535), .Z1_f (new_AGEMA_signal_8536) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T14), .A0_f (new_AGEMA_signal_7946), .A1_t (new_AGEMA_signal_7947), .A1_f (new_AGEMA_signal_7948), .B0_t (SubBytesIns_Inst_Sbox_12_M1), .B0_f (new_AGEMA_signal_7961), .B1_t (new_AGEMA_signal_7962), .B1_f (new_AGEMA_signal_7963), .Z0_t (SubBytesIns_Inst_Sbox_12_M3), .Z0_f (new_AGEMA_signal_8537), .Z1_t (new_AGEMA_signal_8538), .Z1_f (new_AGEMA_signal_8539) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T19), .A0_f (new_AGEMA_signal_7231), .A1_t (new_AGEMA_signal_7232), .A1_f (new_AGEMA_signal_7233), .B0_t (ciphertext_s0_t[96]), .B0_f (ciphertext_s0_f[96]), .B1_t (ciphertext_s1_t[96]), .B1_f (ciphertext_s1_f[96]), .Z0_t (SubBytesIns_Inst_Sbox_12_M4), .Z0_f (new_AGEMA_signal_7964), .Z1_t (new_AGEMA_signal_7965), .Z1_f (new_AGEMA_signal_7966) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M4), .A0_f (new_AGEMA_signal_7964), .A1_t (new_AGEMA_signal_7965), .A1_f (new_AGEMA_signal_7966), .B0_t (SubBytesIns_Inst_Sbox_12_M1), .B0_f (new_AGEMA_signal_7961), .B1_t (new_AGEMA_signal_7962), .B1_f (new_AGEMA_signal_7963), .Z0_t (SubBytesIns_Inst_Sbox_12_M5), .Z0_f (new_AGEMA_signal_8540), .Z1_t (new_AGEMA_signal_8541), .Z1_f (new_AGEMA_signal_8542) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T3), .A0_f (new_AGEMA_signal_6712), .A1_t (new_AGEMA_signal_6713), .A1_f (new_AGEMA_signal_6714), .B0_t (SubBytesIns_Inst_Sbox_12_T16), .B0_f (new_AGEMA_signal_7228), .B1_t (new_AGEMA_signal_7229), .B1_f (new_AGEMA_signal_7230), .Z0_t (SubBytesIns_Inst_Sbox_12_M6), .Z0_f (new_AGEMA_signal_7967), .Z1_t (new_AGEMA_signal_7968), .Z1_f (new_AGEMA_signal_7969) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T22), .A0_f (new_AGEMA_signal_7234), .A1_t (new_AGEMA_signal_7235), .A1_f (new_AGEMA_signal_7236), .B0_t (SubBytesIns_Inst_Sbox_12_T9), .B0_f (new_AGEMA_signal_7219), .B1_t (new_AGEMA_signal_7220), .B1_f (new_AGEMA_signal_7221), .Z0_t (SubBytesIns_Inst_Sbox_12_M7), .Z0_f (new_AGEMA_signal_7970), .Z1_t (new_AGEMA_signal_7971), .Z1_f (new_AGEMA_signal_7972) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T26), .A0_f (new_AGEMA_signal_7958), .A1_t (new_AGEMA_signal_7959), .A1_f (new_AGEMA_signal_7960), .B0_t (SubBytesIns_Inst_Sbox_12_M6), .B0_f (new_AGEMA_signal_7967), .B1_t (new_AGEMA_signal_7968), .B1_f (new_AGEMA_signal_7969), .Z0_t (SubBytesIns_Inst_Sbox_12_M8), .Z0_f (new_AGEMA_signal_8543), .Z1_t (new_AGEMA_signal_8544), .Z1_f (new_AGEMA_signal_8545) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T20), .A0_f (new_AGEMA_signal_7952), .A1_t (new_AGEMA_signal_7953), .A1_f (new_AGEMA_signal_7954), .B0_t (SubBytesIns_Inst_Sbox_12_T17), .B0_f (new_AGEMA_signal_7949), .B1_t (new_AGEMA_signal_7950), .B1_f (new_AGEMA_signal_7951), .Z0_t (SubBytesIns_Inst_Sbox_12_M9), .Z0_f (new_AGEMA_signal_8546), .Z1_t (new_AGEMA_signal_8547), .Z1_f (new_AGEMA_signal_8548) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M9), .A0_f (new_AGEMA_signal_8546), .A1_t (new_AGEMA_signal_8547), .A1_f (new_AGEMA_signal_8548), .B0_t (SubBytesIns_Inst_Sbox_12_M6), .B0_f (new_AGEMA_signal_7967), .B1_t (new_AGEMA_signal_7968), .B1_f (new_AGEMA_signal_7969), .Z0_t (SubBytesIns_Inst_Sbox_12_M10), .Z0_f (new_AGEMA_signal_8876), .Z1_t (new_AGEMA_signal_8877), .Z1_f (new_AGEMA_signal_8878) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T1), .A0_f (new_AGEMA_signal_6706), .A1_t (new_AGEMA_signal_6707), .A1_f (new_AGEMA_signal_6708), .B0_t (SubBytesIns_Inst_Sbox_12_T15), .B0_f (new_AGEMA_signal_7225), .B1_t (new_AGEMA_signal_7226), .B1_f (new_AGEMA_signal_7227), .Z0_t (SubBytesIns_Inst_Sbox_12_M11), .Z0_f (new_AGEMA_signal_7973), .Z1_t (new_AGEMA_signal_7974), .Z1_f (new_AGEMA_signal_7975) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T4), .A0_f (new_AGEMA_signal_6715), .A1_t (new_AGEMA_signal_6716), .A1_f (new_AGEMA_signal_6717), .B0_t (SubBytesIns_Inst_Sbox_12_T27), .B0_f (new_AGEMA_signal_7237), .B1_t (new_AGEMA_signal_7238), .B1_f (new_AGEMA_signal_7239), .Z0_t (SubBytesIns_Inst_Sbox_12_M12), .Z0_f (new_AGEMA_signal_7976), .Z1_t (new_AGEMA_signal_7977), .Z1_f (new_AGEMA_signal_7978) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M12), .A0_f (new_AGEMA_signal_7976), .A1_t (new_AGEMA_signal_7977), .A1_f (new_AGEMA_signal_7978), .B0_t (SubBytesIns_Inst_Sbox_12_M11), .B0_f (new_AGEMA_signal_7973), .B1_t (new_AGEMA_signal_7974), .B1_f (new_AGEMA_signal_7975), .Z0_t (SubBytesIns_Inst_Sbox_12_M13), .Z0_f (new_AGEMA_signal_8549), .Z1_t (new_AGEMA_signal_8550), .Z1_f (new_AGEMA_signal_8551) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T2), .A0_f (new_AGEMA_signal_6709), .A1_t (new_AGEMA_signal_6710), .A1_f (new_AGEMA_signal_6711), .B0_t (SubBytesIns_Inst_Sbox_12_T10), .B0_f (new_AGEMA_signal_7943), .B1_t (new_AGEMA_signal_7944), .B1_f (new_AGEMA_signal_7945), .Z0_t (SubBytesIns_Inst_Sbox_12_M14), .Z0_f (new_AGEMA_signal_8552), .Z1_t (new_AGEMA_signal_8553), .Z1_f (new_AGEMA_signal_8554) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M14), .A0_f (new_AGEMA_signal_8552), .A1_t (new_AGEMA_signal_8553), .A1_f (new_AGEMA_signal_8554), .B0_t (SubBytesIns_Inst_Sbox_12_M11), .B0_f (new_AGEMA_signal_7973), .B1_t (new_AGEMA_signal_7974), .B1_f (new_AGEMA_signal_7975), .Z0_t (SubBytesIns_Inst_Sbox_12_M15), .Z0_f (new_AGEMA_signal_8879), .Z1_t (new_AGEMA_signal_8880), .Z1_f (new_AGEMA_signal_8881) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M3), .A0_f (new_AGEMA_signal_8537), .A1_t (new_AGEMA_signal_8538), .A1_f (new_AGEMA_signal_8539), .B0_t (SubBytesIns_Inst_Sbox_12_M2), .B0_f (new_AGEMA_signal_8534), .B1_t (new_AGEMA_signal_8535), .B1_f (new_AGEMA_signal_8536), .Z0_t (SubBytesIns_Inst_Sbox_12_M16), .Z0_f (new_AGEMA_signal_8882), .Z1_t (new_AGEMA_signal_8883), .Z1_f (new_AGEMA_signal_8884) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M5), .A0_f (new_AGEMA_signal_8540), .A1_t (new_AGEMA_signal_8541), .A1_f (new_AGEMA_signal_8542), .B0_t (SubBytesIns_Inst_Sbox_12_T24), .B0_f (new_AGEMA_signal_8528), .B1_t (new_AGEMA_signal_8529), .B1_f (new_AGEMA_signal_8530), .Z0_t (SubBytesIns_Inst_Sbox_12_M17), .Z0_f (new_AGEMA_signal_8885), .Z1_t (new_AGEMA_signal_8886), .Z1_f (new_AGEMA_signal_8887) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M8), .A0_f (new_AGEMA_signal_8543), .A1_t (new_AGEMA_signal_8544), .A1_f (new_AGEMA_signal_8545), .B0_t (SubBytesIns_Inst_Sbox_12_M7), .B0_f (new_AGEMA_signal_7970), .B1_t (new_AGEMA_signal_7971), .B1_f (new_AGEMA_signal_7972), .Z0_t (SubBytesIns_Inst_Sbox_12_M18), .Z0_f (new_AGEMA_signal_8888), .Z1_t (new_AGEMA_signal_8889), .Z1_f (new_AGEMA_signal_8890) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M10), .A0_f (new_AGEMA_signal_8876), .A1_t (new_AGEMA_signal_8877), .A1_f (new_AGEMA_signal_8878), .B0_t (SubBytesIns_Inst_Sbox_12_M15), .B0_f (new_AGEMA_signal_8879), .B1_t (new_AGEMA_signal_8880), .B1_f (new_AGEMA_signal_8881), .Z0_t (SubBytesIns_Inst_Sbox_12_M19), .Z0_f (new_AGEMA_signal_9128), .Z1_t (new_AGEMA_signal_9129), .Z1_f (new_AGEMA_signal_9130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M16), .A0_f (new_AGEMA_signal_8882), .A1_t (new_AGEMA_signal_8883), .A1_f (new_AGEMA_signal_8884), .B0_t (SubBytesIns_Inst_Sbox_12_M13), .B0_f (new_AGEMA_signal_8549), .B1_t (new_AGEMA_signal_8550), .B1_f (new_AGEMA_signal_8551), .Z0_t (SubBytesIns_Inst_Sbox_12_M20), .Z0_f (new_AGEMA_signal_9131), .Z1_t (new_AGEMA_signal_9132), .Z1_f (new_AGEMA_signal_9133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M17), .A0_f (new_AGEMA_signal_8885), .A1_t (new_AGEMA_signal_8886), .A1_f (new_AGEMA_signal_8887), .B0_t (SubBytesIns_Inst_Sbox_12_M15), .B0_f (new_AGEMA_signal_8879), .B1_t (new_AGEMA_signal_8880), .B1_f (new_AGEMA_signal_8881), .Z0_t (SubBytesIns_Inst_Sbox_12_M21), .Z0_f (new_AGEMA_signal_9134), .Z1_t (new_AGEMA_signal_9135), .Z1_f (new_AGEMA_signal_9136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M18), .A0_f (new_AGEMA_signal_8888), .A1_t (new_AGEMA_signal_8889), .A1_f (new_AGEMA_signal_8890), .B0_t (SubBytesIns_Inst_Sbox_12_M13), .B0_f (new_AGEMA_signal_8549), .B1_t (new_AGEMA_signal_8550), .B1_f (new_AGEMA_signal_8551), .Z0_t (SubBytesIns_Inst_Sbox_12_M22), .Z0_f (new_AGEMA_signal_9137), .Z1_t (new_AGEMA_signal_9138), .Z1_f (new_AGEMA_signal_9139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M19), .A0_f (new_AGEMA_signal_9128), .A1_t (new_AGEMA_signal_9129), .A1_f (new_AGEMA_signal_9130), .B0_t (SubBytesIns_Inst_Sbox_12_T25), .B0_f (new_AGEMA_signal_8531), .B1_t (new_AGEMA_signal_8532), .B1_f (new_AGEMA_signal_8533), .Z0_t (SubBytesIns_Inst_Sbox_12_M23), .Z0_f (new_AGEMA_signal_9368), .Z1_t (new_AGEMA_signal_9369), .Z1_f (new_AGEMA_signal_9370) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M22), .A0_f (new_AGEMA_signal_9137), .A1_t (new_AGEMA_signal_9138), .A1_f (new_AGEMA_signal_9139), .B0_t (SubBytesIns_Inst_Sbox_12_M23), .B0_f (new_AGEMA_signal_9368), .B1_t (new_AGEMA_signal_9369), .B1_f (new_AGEMA_signal_9370), .Z0_t (SubBytesIns_Inst_Sbox_12_M24), .Z0_f (new_AGEMA_signal_9656), .Z1_t (new_AGEMA_signal_9657), .Z1_f (new_AGEMA_signal_9658) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M22), .A0_f (new_AGEMA_signal_9137), .A1_t (new_AGEMA_signal_9138), .A1_f (new_AGEMA_signal_9139), .B0_t (SubBytesIns_Inst_Sbox_12_M20), .B0_f (new_AGEMA_signal_9131), .B1_t (new_AGEMA_signal_9132), .B1_f (new_AGEMA_signal_9133), .Z0_t (SubBytesIns_Inst_Sbox_12_M25), .Z0_f (new_AGEMA_signal_9371), .Z1_t (new_AGEMA_signal_9372), .Z1_f (new_AGEMA_signal_9373) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M21), .A0_f (new_AGEMA_signal_9134), .A1_t (new_AGEMA_signal_9135), .A1_f (new_AGEMA_signal_9136), .B0_t (SubBytesIns_Inst_Sbox_12_M25), .B0_f (new_AGEMA_signal_9371), .B1_t (new_AGEMA_signal_9372), .B1_f (new_AGEMA_signal_9373), .Z0_t (SubBytesIns_Inst_Sbox_12_M26), .Z0_f (new_AGEMA_signal_9659), .Z1_t (new_AGEMA_signal_9660), .Z1_f (new_AGEMA_signal_9661) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M20), .A0_f (new_AGEMA_signal_9131), .A1_t (new_AGEMA_signal_9132), .A1_f (new_AGEMA_signal_9133), .B0_t (SubBytesIns_Inst_Sbox_12_M21), .B0_f (new_AGEMA_signal_9134), .B1_t (new_AGEMA_signal_9135), .B1_f (new_AGEMA_signal_9136), .Z0_t (SubBytesIns_Inst_Sbox_12_M27), .Z0_f (new_AGEMA_signal_9374), .Z1_t (new_AGEMA_signal_9375), .Z1_f (new_AGEMA_signal_9376) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M23), .A0_f (new_AGEMA_signal_9368), .A1_t (new_AGEMA_signal_9369), .A1_f (new_AGEMA_signal_9370), .B0_t (SubBytesIns_Inst_Sbox_12_M25), .B0_f (new_AGEMA_signal_9371), .B1_t (new_AGEMA_signal_9372), .B1_f (new_AGEMA_signal_9373), .Z0_t (SubBytesIns_Inst_Sbox_12_M28), .Z0_f (new_AGEMA_signal_9662), .Z1_t (new_AGEMA_signal_9663), .Z1_f (new_AGEMA_signal_9664) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M28), .A0_f (new_AGEMA_signal_9662), .A1_t (new_AGEMA_signal_9663), .A1_f (new_AGEMA_signal_9664), .B0_t (SubBytesIns_Inst_Sbox_12_M27), .B0_f (new_AGEMA_signal_9374), .B1_t (new_AGEMA_signal_9375), .B1_f (new_AGEMA_signal_9376), .Z0_t (SubBytesIns_Inst_Sbox_12_M29), .Z0_f (new_AGEMA_signal_9956), .Z1_t (new_AGEMA_signal_9957), .Z1_f (new_AGEMA_signal_9958) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M26), .A0_f (new_AGEMA_signal_9659), .A1_t (new_AGEMA_signal_9660), .A1_f (new_AGEMA_signal_9661), .B0_t (SubBytesIns_Inst_Sbox_12_M24), .B0_f (new_AGEMA_signal_9656), .B1_t (new_AGEMA_signal_9657), .B1_f (new_AGEMA_signal_9658), .Z0_t (SubBytesIns_Inst_Sbox_12_M30), .Z0_f (new_AGEMA_signal_9959), .Z1_t (new_AGEMA_signal_9960), .Z1_f (new_AGEMA_signal_9961) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M20), .A0_f (new_AGEMA_signal_9131), .A1_t (new_AGEMA_signal_9132), .A1_f (new_AGEMA_signal_9133), .B0_t (SubBytesIns_Inst_Sbox_12_M23), .B0_f (new_AGEMA_signal_9368), .B1_t (new_AGEMA_signal_9369), .B1_f (new_AGEMA_signal_9370), .Z0_t (SubBytesIns_Inst_Sbox_12_M31), .Z0_f (new_AGEMA_signal_9665), .Z1_t (new_AGEMA_signal_9666), .Z1_f (new_AGEMA_signal_9667) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M27), .A0_f (new_AGEMA_signal_9374), .A1_t (new_AGEMA_signal_9375), .A1_f (new_AGEMA_signal_9376), .B0_t (SubBytesIns_Inst_Sbox_12_M31), .B0_f (new_AGEMA_signal_9665), .B1_t (new_AGEMA_signal_9666), .B1_f (new_AGEMA_signal_9667), .Z0_t (SubBytesIns_Inst_Sbox_12_M32), .Z0_f (new_AGEMA_signal_9962), .Z1_t (new_AGEMA_signal_9963), .Z1_f (new_AGEMA_signal_9964) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M27), .A0_f (new_AGEMA_signal_9374), .A1_t (new_AGEMA_signal_9375), .A1_f (new_AGEMA_signal_9376), .B0_t (SubBytesIns_Inst_Sbox_12_M25), .B0_f (new_AGEMA_signal_9371), .B1_t (new_AGEMA_signal_9372), .B1_f (new_AGEMA_signal_9373), .Z0_t (SubBytesIns_Inst_Sbox_12_M33), .Z0_f (new_AGEMA_signal_9668), .Z1_t (new_AGEMA_signal_9669), .Z1_f (new_AGEMA_signal_9670) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M21), .A0_f (new_AGEMA_signal_9134), .A1_t (new_AGEMA_signal_9135), .A1_f (new_AGEMA_signal_9136), .B0_t (SubBytesIns_Inst_Sbox_12_M22), .B0_f (new_AGEMA_signal_9137), .B1_t (new_AGEMA_signal_9138), .B1_f (new_AGEMA_signal_9139), .Z0_t (SubBytesIns_Inst_Sbox_12_M34), .Z0_f (new_AGEMA_signal_9377), .Z1_t (new_AGEMA_signal_9378), .Z1_f (new_AGEMA_signal_9379) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M24), .A0_f (new_AGEMA_signal_9656), .A1_t (new_AGEMA_signal_9657), .A1_f (new_AGEMA_signal_9658), .B0_t (SubBytesIns_Inst_Sbox_12_M34), .B0_f (new_AGEMA_signal_9377), .B1_t (new_AGEMA_signal_9378), .B1_f (new_AGEMA_signal_9379), .Z0_t (SubBytesIns_Inst_Sbox_12_M35), .Z0_f (new_AGEMA_signal_9965), .Z1_t (new_AGEMA_signal_9966), .Z1_f (new_AGEMA_signal_9967) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M24), .A0_f (new_AGEMA_signal_9656), .A1_t (new_AGEMA_signal_9657), .A1_f (new_AGEMA_signal_9658), .B0_t (SubBytesIns_Inst_Sbox_12_M25), .B0_f (new_AGEMA_signal_9371), .B1_t (new_AGEMA_signal_9372), .B1_f (new_AGEMA_signal_9373), .Z0_t (SubBytesIns_Inst_Sbox_12_M36), .Z0_f (new_AGEMA_signal_9968), .Z1_t (new_AGEMA_signal_9969), .Z1_f (new_AGEMA_signal_9970) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M21), .A0_f (new_AGEMA_signal_9134), .A1_t (new_AGEMA_signal_9135), .A1_f (new_AGEMA_signal_9136), .B0_t (SubBytesIns_Inst_Sbox_12_M29), .B0_f (new_AGEMA_signal_9956), .B1_t (new_AGEMA_signal_9957), .B1_f (new_AGEMA_signal_9958), .Z0_t (SubBytesIns_Inst_Sbox_12_M37), .Z0_f (new_AGEMA_signal_10208), .Z1_t (new_AGEMA_signal_10209), .Z1_f (new_AGEMA_signal_10210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M32), .A0_f (new_AGEMA_signal_9962), .A1_t (new_AGEMA_signal_9963), .A1_f (new_AGEMA_signal_9964), .B0_t (SubBytesIns_Inst_Sbox_12_M33), .B0_f (new_AGEMA_signal_9668), .B1_t (new_AGEMA_signal_9669), .B1_f (new_AGEMA_signal_9670), .Z0_t (SubBytesIns_Inst_Sbox_12_M38), .Z0_f (new_AGEMA_signal_10211), .Z1_t (new_AGEMA_signal_10212), .Z1_f (new_AGEMA_signal_10213) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M23), .A0_f (new_AGEMA_signal_9368), .A1_t (new_AGEMA_signal_9369), .A1_f (new_AGEMA_signal_9370), .B0_t (SubBytesIns_Inst_Sbox_12_M30), .B0_f (new_AGEMA_signal_9959), .B1_t (new_AGEMA_signal_9960), .B1_f (new_AGEMA_signal_9961), .Z0_t (SubBytesIns_Inst_Sbox_12_M39), .Z0_f (new_AGEMA_signal_10214), .Z1_t (new_AGEMA_signal_10215), .Z1_f (new_AGEMA_signal_10216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M35), .A0_f (new_AGEMA_signal_9965), .A1_t (new_AGEMA_signal_9966), .A1_f (new_AGEMA_signal_9967), .B0_t (SubBytesIns_Inst_Sbox_12_M36), .B0_f (new_AGEMA_signal_9968), .B1_t (new_AGEMA_signal_9969), .B1_f (new_AGEMA_signal_9970), .Z0_t (SubBytesIns_Inst_Sbox_12_M40), .Z0_f (new_AGEMA_signal_10217), .Z1_t (new_AGEMA_signal_10218), .Z1_f (new_AGEMA_signal_10219) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M38), .A0_f (new_AGEMA_signal_10211), .A1_t (new_AGEMA_signal_10212), .A1_f (new_AGEMA_signal_10213), .B0_t (SubBytesIns_Inst_Sbox_12_M40), .B0_f (new_AGEMA_signal_10217), .B1_t (new_AGEMA_signal_10218), .B1_f (new_AGEMA_signal_10219), .Z0_t (SubBytesIns_Inst_Sbox_12_M41), .Z0_f (new_AGEMA_signal_10832), .Z1_t (new_AGEMA_signal_10833), .Z1_f (new_AGEMA_signal_10834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M37), .A0_f (new_AGEMA_signal_10208), .A1_t (new_AGEMA_signal_10209), .A1_f (new_AGEMA_signal_10210), .B0_t (SubBytesIns_Inst_Sbox_12_M39), .B0_f (new_AGEMA_signal_10214), .B1_t (new_AGEMA_signal_10215), .B1_f (new_AGEMA_signal_10216), .Z0_t (SubBytesIns_Inst_Sbox_12_M42), .Z0_f (new_AGEMA_signal_10835), .Z1_t (new_AGEMA_signal_10836), .Z1_f (new_AGEMA_signal_10837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M37), .A0_f (new_AGEMA_signal_10208), .A1_t (new_AGEMA_signal_10209), .A1_f (new_AGEMA_signal_10210), .B0_t (SubBytesIns_Inst_Sbox_12_M38), .B0_f (new_AGEMA_signal_10211), .B1_t (new_AGEMA_signal_10212), .B1_f (new_AGEMA_signal_10213), .Z0_t (SubBytesIns_Inst_Sbox_12_M43), .Z0_f (new_AGEMA_signal_10838), .Z1_t (new_AGEMA_signal_10839), .Z1_f (new_AGEMA_signal_10840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M39), .A0_f (new_AGEMA_signal_10214), .A1_t (new_AGEMA_signal_10215), .A1_f (new_AGEMA_signal_10216), .B0_t (SubBytesIns_Inst_Sbox_12_M40), .B0_f (new_AGEMA_signal_10217), .B1_t (new_AGEMA_signal_10218), .B1_f (new_AGEMA_signal_10219), .Z0_t (SubBytesIns_Inst_Sbox_12_M44), .Z0_f (new_AGEMA_signal_10841), .Z1_t (new_AGEMA_signal_10842), .Z1_f (new_AGEMA_signal_10843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M42), .A0_f (new_AGEMA_signal_10835), .A1_t (new_AGEMA_signal_10836), .A1_f (new_AGEMA_signal_10837), .B0_t (SubBytesIns_Inst_Sbox_12_M41), .B0_f (new_AGEMA_signal_10832), .B1_t (new_AGEMA_signal_10833), .B1_f (new_AGEMA_signal_10834), .Z0_t (SubBytesIns_Inst_Sbox_12_M45), .Z0_f (new_AGEMA_signal_11552), .Z1_t (new_AGEMA_signal_11553), .Z1_f (new_AGEMA_signal_11554) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M44), .A0_f (new_AGEMA_signal_10841), .A1_t (new_AGEMA_signal_10842), .A1_f (new_AGEMA_signal_10843), .B0_t (SubBytesIns_Inst_Sbox_12_T6), .B0_f (new_AGEMA_signal_7216), .B1_t (new_AGEMA_signal_7217), .B1_f (new_AGEMA_signal_7218), .Z0_t (SubBytesIns_Inst_Sbox_12_M46), .Z0_f (new_AGEMA_signal_11555), .Z1_t (new_AGEMA_signal_11556), .Z1_f (new_AGEMA_signal_11557) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M40), .A0_f (new_AGEMA_signal_10217), .A1_t (new_AGEMA_signal_10218), .A1_f (new_AGEMA_signal_10219), .B0_t (SubBytesIns_Inst_Sbox_12_T8), .B0_f (new_AGEMA_signal_7940), .B1_t (new_AGEMA_signal_7941), .B1_f (new_AGEMA_signal_7942), .Z0_t (SubBytesIns_Inst_Sbox_12_M47), .Z0_f (new_AGEMA_signal_10844), .Z1_t (new_AGEMA_signal_10845), .Z1_f (new_AGEMA_signal_10846) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M39), .A0_f (new_AGEMA_signal_10214), .A1_t (new_AGEMA_signal_10215), .A1_f (new_AGEMA_signal_10216), .B0_t (ciphertext_s0_t[96]), .B0_f (ciphertext_s0_f[96]), .B1_t (ciphertext_s1_t[96]), .B1_f (ciphertext_s1_f[96]), .Z0_t (SubBytesIns_Inst_Sbox_12_M48), .Z0_f (new_AGEMA_signal_10847), .Z1_t (new_AGEMA_signal_10848), .Z1_f (new_AGEMA_signal_10849) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M43), .A0_f (new_AGEMA_signal_10838), .A1_t (new_AGEMA_signal_10839), .A1_f (new_AGEMA_signal_10840), .B0_t (SubBytesIns_Inst_Sbox_12_T16), .B0_f (new_AGEMA_signal_7228), .B1_t (new_AGEMA_signal_7229), .B1_f (new_AGEMA_signal_7230), .Z0_t (SubBytesIns_Inst_Sbox_12_M49), .Z0_f (new_AGEMA_signal_11558), .Z1_t (new_AGEMA_signal_11559), .Z1_f (new_AGEMA_signal_11560) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M38), .A0_f (new_AGEMA_signal_10211), .A1_t (new_AGEMA_signal_10212), .A1_f (new_AGEMA_signal_10213), .B0_t (SubBytesIns_Inst_Sbox_12_T9), .B0_f (new_AGEMA_signal_7219), .B1_t (new_AGEMA_signal_7220), .B1_f (new_AGEMA_signal_7221), .Z0_t (SubBytesIns_Inst_Sbox_12_M50), .Z0_f (new_AGEMA_signal_10850), .Z1_t (new_AGEMA_signal_10851), .Z1_f (new_AGEMA_signal_10852) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M37), .A0_f (new_AGEMA_signal_10208), .A1_t (new_AGEMA_signal_10209), .A1_f (new_AGEMA_signal_10210), .B0_t (SubBytesIns_Inst_Sbox_12_T17), .B0_f (new_AGEMA_signal_7949), .B1_t (new_AGEMA_signal_7950), .B1_f (new_AGEMA_signal_7951), .Z0_t (SubBytesIns_Inst_Sbox_12_M51), .Z0_f (new_AGEMA_signal_10853), .Z1_t (new_AGEMA_signal_10854), .Z1_f (new_AGEMA_signal_10855) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M42), .A0_f (new_AGEMA_signal_10835), .A1_t (new_AGEMA_signal_10836), .A1_f (new_AGEMA_signal_10837), .B0_t (SubBytesIns_Inst_Sbox_12_T15), .B0_f (new_AGEMA_signal_7225), .B1_t (new_AGEMA_signal_7226), .B1_f (new_AGEMA_signal_7227), .Z0_t (SubBytesIns_Inst_Sbox_12_M52), .Z0_f (new_AGEMA_signal_11561), .Z1_t (new_AGEMA_signal_11562), .Z1_f (new_AGEMA_signal_11563) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M45), .A0_f (new_AGEMA_signal_11552), .A1_t (new_AGEMA_signal_11553), .A1_f (new_AGEMA_signal_11554), .B0_t (SubBytesIns_Inst_Sbox_12_T27), .B0_f (new_AGEMA_signal_7237), .B1_t (new_AGEMA_signal_7238), .B1_f (new_AGEMA_signal_7239), .Z0_t (SubBytesIns_Inst_Sbox_12_M53), .Z0_f (new_AGEMA_signal_12176), .Z1_t (new_AGEMA_signal_12177), .Z1_f (new_AGEMA_signal_12178) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M41), .A0_f (new_AGEMA_signal_10832), .A1_t (new_AGEMA_signal_10833), .A1_f (new_AGEMA_signal_10834), .B0_t (SubBytesIns_Inst_Sbox_12_T10), .B0_f (new_AGEMA_signal_7943), .B1_t (new_AGEMA_signal_7944), .B1_f (new_AGEMA_signal_7945), .Z0_t (SubBytesIns_Inst_Sbox_12_M54), .Z0_f (new_AGEMA_signal_11564), .Z1_t (new_AGEMA_signal_11565), .Z1_f (new_AGEMA_signal_11566) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M44), .A0_f (new_AGEMA_signal_10841), .A1_t (new_AGEMA_signal_10842), .A1_f (new_AGEMA_signal_10843), .B0_t (SubBytesIns_Inst_Sbox_12_T13), .B0_f (new_AGEMA_signal_7222), .B1_t (new_AGEMA_signal_7223), .B1_f (new_AGEMA_signal_7224), .Z0_t (SubBytesIns_Inst_Sbox_12_M55), .Z0_f (new_AGEMA_signal_11567), .Z1_t (new_AGEMA_signal_11568), .Z1_f (new_AGEMA_signal_11569) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M40), .A0_f (new_AGEMA_signal_10217), .A1_t (new_AGEMA_signal_10218), .A1_f (new_AGEMA_signal_10219), .B0_t (SubBytesIns_Inst_Sbox_12_T23), .B0_f (new_AGEMA_signal_7955), .B1_t (new_AGEMA_signal_7956), .B1_f (new_AGEMA_signal_7957), .Z0_t (SubBytesIns_Inst_Sbox_12_M56), .Z0_f (new_AGEMA_signal_10856), .Z1_t (new_AGEMA_signal_10857), .Z1_f (new_AGEMA_signal_10858) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M39), .A0_f (new_AGEMA_signal_10214), .A1_t (new_AGEMA_signal_10215), .A1_f (new_AGEMA_signal_10216), .B0_t (SubBytesIns_Inst_Sbox_12_T19), .B0_f (new_AGEMA_signal_7231), .B1_t (new_AGEMA_signal_7232), .B1_f (new_AGEMA_signal_7233), .Z0_t (SubBytesIns_Inst_Sbox_12_M57), .Z0_f (new_AGEMA_signal_10859), .Z1_t (new_AGEMA_signal_10860), .Z1_f (new_AGEMA_signal_10861) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M43), .A0_f (new_AGEMA_signal_10838), .A1_t (new_AGEMA_signal_10839), .A1_f (new_AGEMA_signal_10840), .B0_t (SubBytesIns_Inst_Sbox_12_T3), .B0_f (new_AGEMA_signal_6712), .B1_t (new_AGEMA_signal_6713), .B1_f (new_AGEMA_signal_6714), .Z0_t (SubBytesIns_Inst_Sbox_12_M58), .Z0_f (new_AGEMA_signal_11570), .Z1_t (new_AGEMA_signal_11571), .Z1_f (new_AGEMA_signal_11572) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M38), .A0_f (new_AGEMA_signal_10211), .A1_t (new_AGEMA_signal_10212), .A1_f (new_AGEMA_signal_10213), .B0_t (SubBytesIns_Inst_Sbox_12_T22), .B0_f (new_AGEMA_signal_7234), .B1_t (new_AGEMA_signal_7235), .B1_f (new_AGEMA_signal_7236), .Z0_t (SubBytesIns_Inst_Sbox_12_M59), .Z0_f (new_AGEMA_signal_10862), .Z1_t (new_AGEMA_signal_10863), .Z1_f (new_AGEMA_signal_10864) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M37), .A0_f (new_AGEMA_signal_10208), .A1_t (new_AGEMA_signal_10209), .A1_f (new_AGEMA_signal_10210), .B0_t (SubBytesIns_Inst_Sbox_12_T20), .B0_f (new_AGEMA_signal_7952), .B1_t (new_AGEMA_signal_7953), .B1_f (new_AGEMA_signal_7954), .Z0_t (SubBytesIns_Inst_Sbox_12_M60), .Z0_f (new_AGEMA_signal_10865), .Z1_t (new_AGEMA_signal_10866), .Z1_f (new_AGEMA_signal_10867) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M42), .A0_f (new_AGEMA_signal_10835), .A1_t (new_AGEMA_signal_10836), .A1_f (new_AGEMA_signal_10837), .B0_t (SubBytesIns_Inst_Sbox_12_T1), .B0_f (new_AGEMA_signal_6706), .B1_t (new_AGEMA_signal_6707), .B1_f (new_AGEMA_signal_6708), .Z0_t (SubBytesIns_Inst_Sbox_12_M61), .Z0_f (new_AGEMA_signal_11573), .Z1_t (new_AGEMA_signal_11574), .Z1_f (new_AGEMA_signal_11575) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M45), .A0_f (new_AGEMA_signal_11552), .A1_t (new_AGEMA_signal_11553), .A1_f (new_AGEMA_signal_11554), .B0_t (SubBytesIns_Inst_Sbox_12_T4), .B0_f (new_AGEMA_signal_6715), .B1_t (new_AGEMA_signal_6716), .B1_f (new_AGEMA_signal_6717), .Z0_t (SubBytesIns_Inst_Sbox_12_M62), .Z0_f (new_AGEMA_signal_12179), .Z1_t (new_AGEMA_signal_12180), .Z1_f (new_AGEMA_signal_12181) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M41), .A0_f (new_AGEMA_signal_10832), .A1_t (new_AGEMA_signal_10833), .A1_f (new_AGEMA_signal_10834), .B0_t (SubBytesIns_Inst_Sbox_12_T2), .B0_f (new_AGEMA_signal_6709), .B1_t (new_AGEMA_signal_6710), .B1_f (new_AGEMA_signal_6711), .Z0_t (SubBytesIns_Inst_Sbox_12_M63), .Z0_f (new_AGEMA_signal_11576), .Z1_t (new_AGEMA_signal_11577), .Z1_f (new_AGEMA_signal_11578) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M61), .A0_f (new_AGEMA_signal_11573), .A1_t (new_AGEMA_signal_11574), .A1_f (new_AGEMA_signal_11575), .B0_t (SubBytesIns_Inst_Sbox_12_M62), .B0_f (new_AGEMA_signal_12179), .B1_t (new_AGEMA_signal_12180), .B1_f (new_AGEMA_signal_12181), .Z0_t (SubBytesIns_Inst_Sbox_12_L0), .Z0_f (new_AGEMA_signal_12728), .Z1_t (new_AGEMA_signal_12729), .Z1_f (new_AGEMA_signal_12730) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M50), .A0_f (new_AGEMA_signal_10850), .A1_t (new_AGEMA_signal_10851), .A1_f (new_AGEMA_signal_10852), .B0_t (SubBytesIns_Inst_Sbox_12_M56), .B0_f (new_AGEMA_signal_10856), .B1_t (new_AGEMA_signal_10857), .B1_f (new_AGEMA_signal_10858), .Z0_t (SubBytesIns_Inst_Sbox_12_L1), .Z0_f (new_AGEMA_signal_11579), .Z1_t (new_AGEMA_signal_11580), .Z1_f (new_AGEMA_signal_11581) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M46), .A0_f (new_AGEMA_signal_11555), .A1_t (new_AGEMA_signal_11556), .A1_f (new_AGEMA_signal_11557), .B0_t (SubBytesIns_Inst_Sbox_12_M48), .B0_f (new_AGEMA_signal_10847), .B1_t (new_AGEMA_signal_10848), .B1_f (new_AGEMA_signal_10849), .Z0_t (SubBytesIns_Inst_Sbox_12_L2), .Z0_f (new_AGEMA_signal_12182), .Z1_t (new_AGEMA_signal_12183), .Z1_f (new_AGEMA_signal_12184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M47), .A0_f (new_AGEMA_signal_10844), .A1_t (new_AGEMA_signal_10845), .A1_f (new_AGEMA_signal_10846), .B0_t (SubBytesIns_Inst_Sbox_12_M55), .B0_f (new_AGEMA_signal_11567), .B1_t (new_AGEMA_signal_11568), .B1_f (new_AGEMA_signal_11569), .Z0_t (SubBytesIns_Inst_Sbox_12_L3), .Z0_f (new_AGEMA_signal_12185), .Z1_t (new_AGEMA_signal_12186), .Z1_f (new_AGEMA_signal_12187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M54), .A0_f (new_AGEMA_signal_11564), .A1_t (new_AGEMA_signal_11565), .A1_f (new_AGEMA_signal_11566), .B0_t (SubBytesIns_Inst_Sbox_12_M58), .B0_f (new_AGEMA_signal_11570), .B1_t (new_AGEMA_signal_11571), .B1_f (new_AGEMA_signal_11572), .Z0_t (SubBytesIns_Inst_Sbox_12_L4), .Z0_f (new_AGEMA_signal_12188), .Z1_t (new_AGEMA_signal_12189), .Z1_f (new_AGEMA_signal_12190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M49), .A0_f (new_AGEMA_signal_11558), .A1_t (new_AGEMA_signal_11559), .A1_f (new_AGEMA_signal_11560), .B0_t (SubBytesIns_Inst_Sbox_12_M61), .B0_f (new_AGEMA_signal_11573), .B1_t (new_AGEMA_signal_11574), .B1_f (new_AGEMA_signal_11575), .Z0_t (SubBytesIns_Inst_Sbox_12_L5), .Z0_f (new_AGEMA_signal_12191), .Z1_t (new_AGEMA_signal_12192), .Z1_f (new_AGEMA_signal_12193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M62), .A0_f (new_AGEMA_signal_12179), .A1_t (new_AGEMA_signal_12180), .A1_f (new_AGEMA_signal_12181), .B0_t (SubBytesIns_Inst_Sbox_12_L5), .B0_f (new_AGEMA_signal_12191), .B1_t (new_AGEMA_signal_12192), .B1_f (new_AGEMA_signal_12193), .Z0_t (SubBytesIns_Inst_Sbox_12_L6), .Z0_f (new_AGEMA_signal_12731), .Z1_t (new_AGEMA_signal_12732), .Z1_f (new_AGEMA_signal_12733) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M46), .A0_f (new_AGEMA_signal_11555), .A1_t (new_AGEMA_signal_11556), .A1_f (new_AGEMA_signal_11557), .B0_t (SubBytesIns_Inst_Sbox_12_L3), .B0_f (new_AGEMA_signal_12185), .B1_t (new_AGEMA_signal_12186), .B1_f (new_AGEMA_signal_12187), .Z0_t (SubBytesIns_Inst_Sbox_12_L7), .Z0_f (new_AGEMA_signal_12734), .Z1_t (new_AGEMA_signal_12735), .Z1_f (new_AGEMA_signal_12736) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M51), .A0_f (new_AGEMA_signal_10853), .A1_t (new_AGEMA_signal_10854), .A1_f (new_AGEMA_signal_10855), .B0_t (SubBytesIns_Inst_Sbox_12_M59), .B0_f (new_AGEMA_signal_10862), .B1_t (new_AGEMA_signal_10863), .B1_f (new_AGEMA_signal_10864), .Z0_t (SubBytesIns_Inst_Sbox_12_L8), .Z0_f (new_AGEMA_signal_11582), .Z1_t (new_AGEMA_signal_11583), .Z1_f (new_AGEMA_signal_11584) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M52), .A0_f (new_AGEMA_signal_11561), .A1_t (new_AGEMA_signal_11562), .A1_f (new_AGEMA_signal_11563), .B0_t (SubBytesIns_Inst_Sbox_12_M53), .B0_f (new_AGEMA_signal_12176), .B1_t (new_AGEMA_signal_12177), .B1_f (new_AGEMA_signal_12178), .Z0_t (SubBytesIns_Inst_Sbox_12_L9), .Z0_f (new_AGEMA_signal_12737), .Z1_t (new_AGEMA_signal_12738), .Z1_f (new_AGEMA_signal_12739) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M53), .A0_f (new_AGEMA_signal_12176), .A1_t (new_AGEMA_signal_12177), .A1_f (new_AGEMA_signal_12178), .B0_t (SubBytesIns_Inst_Sbox_12_L4), .B0_f (new_AGEMA_signal_12188), .B1_t (new_AGEMA_signal_12189), .B1_f (new_AGEMA_signal_12190), .Z0_t (SubBytesIns_Inst_Sbox_12_L10), .Z0_f (new_AGEMA_signal_12740), .Z1_t (new_AGEMA_signal_12741), .Z1_f (new_AGEMA_signal_12742) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M60), .A0_f (new_AGEMA_signal_10865), .A1_t (new_AGEMA_signal_10866), .A1_f (new_AGEMA_signal_10867), .B0_t (SubBytesIns_Inst_Sbox_12_L2), .B0_f (new_AGEMA_signal_12182), .B1_t (new_AGEMA_signal_12183), .B1_f (new_AGEMA_signal_12184), .Z0_t (SubBytesIns_Inst_Sbox_12_L11), .Z0_f (new_AGEMA_signal_12743), .Z1_t (new_AGEMA_signal_12744), .Z1_f (new_AGEMA_signal_12745) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M48), .A0_f (new_AGEMA_signal_10847), .A1_t (new_AGEMA_signal_10848), .A1_f (new_AGEMA_signal_10849), .B0_t (SubBytesIns_Inst_Sbox_12_M51), .B0_f (new_AGEMA_signal_10853), .B1_t (new_AGEMA_signal_10854), .B1_f (new_AGEMA_signal_10855), .Z0_t (SubBytesIns_Inst_Sbox_12_L12), .Z0_f (new_AGEMA_signal_11585), .Z1_t (new_AGEMA_signal_11586), .Z1_f (new_AGEMA_signal_11587) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M50), .A0_f (new_AGEMA_signal_10850), .A1_t (new_AGEMA_signal_10851), .A1_f (new_AGEMA_signal_10852), .B0_t (SubBytesIns_Inst_Sbox_12_L0), .B0_f (new_AGEMA_signal_12728), .B1_t (new_AGEMA_signal_12729), .B1_f (new_AGEMA_signal_12730), .Z0_t (SubBytesIns_Inst_Sbox_12_L13), .Z0_f (new_AGEMA_signal_13364), .Z1_t (new_AGEMA_signal_13365), .Z1_f (new_AGEMA_signal_13366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M52), .A0_f (new_AGEMA_signal_11561), .A1_t (new_AGEMA_signal_11562), .A1_f (new_AGEMA_signal_11563), .B0_t (SubBytesIns_Inst_Sbox_12_M61), .B0_f (new_AGEMA_signal_11573), .B1_t (new_AGEMA_signal_11574), .B1_f (new_AGEMA_signal_11575), .Z0_t (SubBytesIns_Inst_Sbox_12_L14), .Z0_f (new_AGEMA_signal_12194), .Z1_t (new_AGEMA_signal_12195), .Z1_f (new_AGEMA_signal_12196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M55), .A0_f (new_AGEMA_signal_11567), .A1_t (new_AGEMA_signal_11568), .A1_f (new_AGEMA_signal_11569), .B0_t (SubBytesIns_Inst_Sbox_12_L1), .B0_f (new_AGEMA_signal_11579), .B1_t (new_AGEMA_signal_11580), .B1_f (new_AGEMA_signal_11581), .Z0_t (SubBytesIns_Inst_Sbox_12_L15), .Z0_f (new_AGEMA_signal_12197), .Z1_t (new_AGEMA_signal_12198), .Z1_f (new_AGEMA_signal_12199) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M56), .A0_f (new_AGEMA_signal_10856), .A1_t (new_AGEMA_signal_10857), .A1_f (new_AGEMA_signal_10858), .B0_t (SubBytesIns_Inst_Sbox_12_L0), .B0_f (new_AGEMA_signal_12728), .B1_t (new_AGEMA_signal_12729), .B1_f (new_AGEMA_signal_12730), .Z0_t (SubBytesIns_Inst_Sbox_12_L16), .Z0_f (new_AGEMA_signal_13367), .Z1_t (new_AGEMA_signal_13368), .Z1_f (new_AGEMA_signal_13369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M57), .A0_f (new_AGEMA_signal_10859), .A1_t (new_AGEMA_signal_10860), .A1_f (new_AGEMA_signal_10861), .B0_t (SubBytesIns_Inst_Sbox_12_L1), .B0_f (new_AGEMA_signal_11579), .B1_t (new_AGEMA_signal_11580), .B1_f (new_AGEMA_signal_11581), .Z0_t (SubBytesIns_Inst_Sbox_12_L17), .Z0_f (new_AGEMA_signal_12200), .Z1_t (new_AGEMA_signal_12201), .Z1_f (new_AGEMA_signal_12202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M58), .A0_f (new_AGEMA_signal_11570), .A1_t (new_AGEMA_signal_11571), .A1_f (new_AGEMA_signal_11572), .B0_t (SubBytesIns_Inst_Sbox_12_L8), .B0_f (new_AGEMA_signal_11582), .B1_t (new_AGEMA_signal_11583), .B1_f (new_AGEMA_signal_11584), .Z0_t (SubBytesIns_Inst_Sbox_12_L18), .Z0_f (new_AGEMA_signal_12203), .Z1_t (new_AGEMA_signal_12204), .Z1_f (new_AGEMA_signal_12205) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M63), .A0_f (new_AGEMA_signal_11576), .A1_t (new_AGEMA_signal_11577), .A1_f (new_AGEMA_signal_11578), .B0_t (SubBytesIns_Inst_Sbox_12_L4), .B0_f (new_AGEMA_signal_12188), .B1_t (new_AGEMA_signal_12189), .B1_f (new_AGEMA_signal_12190), .Z0_t (SubBytesIns_Inst_Sbox_12_L19), .Z0_f (new_AGEMA_signal_12746), .Z1_t (new_AGEMA_signal_12747), .Z1_f (new_AGEMA_signal_12748) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L0), .A0_f (new_AGEMA_signal_12728), .A1_t (new_AGEMA_signal_12729), .A1_f (new_AGEMA_signal_12730), .B0_t (SubBytesIns_Inst_Sbox_12_L1), .B0_f (new_AGEMA_signal_11579), .B1_t (new_AGEMA_signal_11580), .B1_f (new_AGEMA_signal_11581), .Z0_t (SubBytesIns_Inst_Sbox_12_L20), .Z0_f (new_AGEMA_signal_13370), .Z1_t (new_AGEMA_signal_13371), .Z1_f (new_AGEMA_signal_13372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L1), .A0_f (new_AGEMA_signal_11579), .A1_t (new_AGEMA_signal_11580), .A1_f (new_AGEMA_signal_11581), .B0_t (SubBytesIns_Inst_Sbox_12_L7), .B0_f (new_AGEMA_signal_12734), .B1_t (new_AGEMA_signal_12735), .B1_f (new_AGEMA_signal_12736), .Z0_t (SubBytesIns_Inst_Sbox_12_L21), .Z0_f (new_AGEMA_signal_13373), .Z1_t (new_AGEMA_signal_13374), .Z1_f (new_AGEMA_signal_13375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L3), .A0_f (new_AGEMA_signal_12185), .A1_t (new_AGEMA_signal_12186), .A1_f (new_AGEMA_signal_12187), .B0_t (SubBytesIns_Inst_Sbox_12_L12), .B0_f (new_AGEMA_signal_11585), .B1_t (new_AGEMA_signal_11586), .B1_f (new_AGEMA_signal_11587), .Z0_t (SubBytesIns_Inst_Sbox_12_L22), .Z0_f (new_AGEMA_signal_12749), .Z1_t (new_AGEMA_signal_12750), .Z1_f (new_AGEMA_signal_12751) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L18), .A0_f (new_AGEMA_signal_12203), .A1_t (new_AGEMA_signal_12204), .A1_f (new_AGEMA_signal_12205), .B0_t (SubBytesIns_Inst_Sbox_12_L2), .B0_f (new_AGEMA_signal_12182), .B1_t (new_AGEMA_signal_12183), .B1_f (new_AGEMA_signal_12184), .Z0_t (SubBytesIns_Inst_Sbox_12_L23), .Z0_f (new_AGEMA_signal_12752), .Z1_t (new_AGEMA_signal_12753), .Z1_f (new_AGEMA_signal_12754) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L15), .A0_f (new_AGEMA_signal_12197), .A1_t (new_AGEMA_signal_12198), .A1_f (new_AGEMA_signal_12199), .B0_t (SubBytesIns_Inst_Sbox_12_L9), .B0_f (new_AGEMA_signal_12737), .B1_t (new_AGEMA_signal_12738), .B1_f (new_AGEMA_signal_12739), .Z0_t (SubBytesIns_Inst_Sbox_12_L24), .Z0_f (new_AGEMA_signal_13376), .Z1_t (new_AGEMA_signal_13377), .Z1_f (new_AGEMA_signal_13378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L6), .A0_f (new_AGEMA_signal_12731), .A1_t (new_AGEMA_signal_12732), .A1_f (new_AGEMA_signal_12733), .B0_t (SubBytesIns_Inst_Sbox_12_L10), .B0_f (new_AGEMA_signal_12740), .B1_t (new_AGEMA_signal_12741), .B1_f (new_AGEMA_signal_12742), .Z0_t (SubBytesIns_Inst_Sbox_12_L25), .Z0_f (new_AGEMA_signal_13379), .Z1_t (new_AGEMA_signal_13380), .Z1_f (new_AGEMA_signal_13381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L7), .A0_f (new_AGEMA_signal_12734), .A1_t (new_AGEMA_signal_12735), .A1_f (new_AGEMA_signal_12736), .B0_t (SubBytesIns_Inst_Sbox_12_L9), .B0_f (new_AGEMA_signal_12737), .B1_t (new_AGEMA_signal_12738), .B1_f (new_AGEMA_signal_12739), .Z0_t (SubBytesIns_Inst_Sbox_12_L26), .Z0_f (new_AGEMA_signal_13382), .Z1_t (new_AGEMA_signal_13383), .Z1_f (new_AGEMA_signal_13384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L8), .A0_f (new_AGEMA_signal_11582), .A1_t (new_AGEMA_signal_11583), .A1_f (new_AGEMA_signal_11584), .B0_t (SubBytesIns_Inst_Sbox_12_L10), .B0_f (new_AGEMA_signal_12740), .B1_t (new_AGEMA_signal_12741), .B1_f (new_AGEMA_signal_12742), .Z0_t (SubBytesIns_Inst_Sbox_12_L27), .Z0_f (new_AGEMA_signal_13385), .Z1_t (new_AGEMA_signal_13386), .Z1_f (new_AGEMA_signal_13387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L11), .A0_f (new_AGEMA_signal_12743), .A1_t (new_AGEMA_signal_12744), .A1_f (new_AGEMA_signal_12745), .B0_t (SubBytesIns_Inst_Sbox_12_L14), .B0_f (new_AGEMA_signal_12194), .B1_t (new_AGEMA_signal_12195), .B1_f (new_AGEMA_signal_12196), .Z0_t (SubBytesIns_Inst_Sbox_12_L28), .Z0_f (new_AGEMA_signal_13388), .Z1_t (new_AGEMA_signal_13389), .Z1_f (new_AGEMA_signal_13390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L11), .A0_f (new_AGEMA_signal_12743), .A1_t (new_AGEMA_signal_12744), .A1_f (new_AGEMA_signal_12745), .B0_t (SubBytesIns_Inst_Sbox_12_L17), .B0_f (new_AGEMA_signal_12200), .B1_t (new_AGEMA_signal_12201), .B1_f (new_AGEMA_signal_12202), .Z0_t (SubBytesIns_Inst_Sbox_12_L29), .Z0_f (new_AGEMA_signal_13391), .Z1_t (new_AGEMA_signal_13392), .Z1_f (new_AGEMA_signal_13393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L6), .A0_f (new_AGEMA_signal_12731), .A1_t (new_AGEMA_signal_12732), .A1_f (new_AGEMA_signal_12733), .B0_t (SubBytesIns_Inst_Sbox_12_L24), .B0_f (new_AGEMA_signal_13376), .B1_t (new_AGEMA_signal_13377), .B1_f (new_AGEMA_signal_13378), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .Z0_f (new_AGEMA_signal_13892), .Z1_t (new_AGEMA_signal_13893), .Z1_f (new_AGEMA_signal_13894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L16), .A0_f (new_AGEMA_signal_13367), .A1_t (new_AGEMA_signal_13368), .A1_f (new_AGEMA_signal_13369), .B0_t (SubBytesIns_Inst_Sbox_12_L26), .B0_f (new_AGEMA_signal_13382), .B1_t (new_AGEMA_signal_13383), .B1_f (new_AGEMA_signal_13384), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .Z0_f (new_AGEMA_signal_13895), .Z1_t (new_AGEMA_signal_13896), .Z1_f (new_AGEMA_signal_13897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L19), .A0_f (new_AGEMA_signal_12746), .A1_t (new_AGEMA_signal_12747), .A1_f (new_AGEMA_signal_12748), .B0_t (SubBytesIns_Inst_Sbox_12_L28), .B0_f (new_AGEMA_signal_13388), .B1_t (new_AGEMA_signal_13389), .B1_f (new_AGEMA_signal_13390), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .Z0_f (new_AGEMA_signal_13898), .Z1_t (new_AGEMA_signal_13899), .Z1_f (new_AGEMA_signal_13900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L6), .A0_f (new_AGEMA_signal_12731), .A1_t (new_AGEMA_signal_12732), .A1_f (new_AGEMA_signal_12733), .B0_t (SubBytesIns_Inst_Sbox_12_L21), .B0_f (new_AGEMA_signal_13373), .B1_t (new_AGEMA_signal_13374), .B1_f (new_AGEMA_signal_13375), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .Z0_f (new_AGEMA_signal_13901), .Z1_t (new_AGEMA_signal_13902), .Z1_f (new_AGEMA_signal_13903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L20), .A0_f (new_AGEMA_signal_13370), .A1_t (new_AGEMA_signal_13371), .A1_f (new_AGEMA_signal_13372), .B0_t (SubBytesIns_Inst_Sbox_12_L22), .B0_f (new_AGEMA_signal_12749), .B1_t (new_AGEMA_signal_12750), .B1_f (new_AGEMA_signal_12751), .Z0_t (MixColumnsInput[67]), .Z0_f (new_AGEMA_signal_13904), .Z1_t (new_AGEMA_signal_13905), .Z1_f (new_AGEMA_signal_13906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L25), .A0_f (new_AGEMA_signal_13379), .A1_t (new_AGEMA_signal_13380), .A1_f (new_AGEMA_signal_13381), .B0_t (SubBytesIns_Inst_Sbox_12_L29), .B0_f (new_AGEMA_signal_13391), .B1_t (new_AGEMA_signal_13392), .B1_f (new_AGEMA_signal_13393), .Z0_t (MixColumnsInput[66]), .Z0_f (new_AGEMA_signal_13907), .Z1_t (new_AGEMA_signal_13908), .Z1_f (new_AGEMA_signal_13909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L13), .A0_f (new_AGEMA_signal_13364), .A1_t (new_AGEMA_signal_13365), .A1_f (new_AGEMA_signal_13366), .B0_t (SubBytesIns_Inst_Sbox_12_L27), .B0_f (new_AGEMA_signal_13385), .B1_t (new_AGEMA_signal_13386), .B1_f (new_AGEMA_signal_13387), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .Z0_f (new_AGEMA_signal_13910), .Z1_t (new_AGEMA_signal_13911), .Z1_f (new_AGEMA_signal_13912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L6), .A0_f (new_AGEMA_signal_12731), .A1_t (new_AGEMA_signal_12732), .A1_f (new_AGEMA_signal_12733), .B0_t (SubBytesIns_Inst_Sbox_12_L23), .B0_f (new_AGEMA_signal_12752), .B1_t (new_AGEMA_signal_12753), .B1_f (new_AGEMA_signal_12754), .Z0_t (MixColumnsInput[64]), .Z0_f (new_AGEMA_signal_13394), .Z1_t (new_AGEMA_signal_13395), .Z1_f (new_AGEMA_signal_13396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (ciphertext_s0_t[108]), .B0_f (ciphertext_s0_f[108]), .B1_t (ciphertext_s1_t[108]), .B1_f (ciphertext_s1_f[108]), .Z0_t (SubBytesIns_Inst_Sbox_13_T1), .Z0_f (new_AGEMA_signal_6736), .Z1_t (new_AGEMA_signal_6737), .Z1_f (new_AGEMA_signal_6738) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (ciphertext_s0_t[106]), .B0_f (ciphertext_s0_f[106]), .B1_t (ciphertext_s1_t[106]), .B1_f (ciphertext_s1_f[106]), .Z0_t (SubBytesIns_Inst_Sbox_13_T2), .Z0_f (new_AGEMA_signal_6739), .Z1_t (new_AGEMA_signal_6740), .Z1_f (new_AGEMA_signal_6741) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (ciphertext_s0_t[105]), .B0_f (ciphertext_s0_f[105]), .B1_t (ciphertext_s1_t[105]), .B1_f (ciphertext_s1_f[105]), .Z0_t (SubBytesIns_Inst_Sbox_13_T3), .Z0_f (new_AGEMA_signal_6742), .Z1_t (new_AGEMA_signal_6743), .Z1_f (new_AGEMA_signal_6744) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[108]), .A0_f (ciphertext_s0_f[108]), .A1_t (ciphertext_s1_t[108]), .A1_f (ciphertext_s1_f[108]), .B0_t (ciphertext_s0_t[106]), .B0_f (ciphertext_s0_f[106]), .B1_t (ciphertext_s1_t[106]), .B1_f (ciphertext_s1_f[106]), .Z0_t (SubBytesIns_Inst_Sbox_13_T4), .Z0_f (new_AGEMA_signal_6745), .Z1_t (new_AGEMA_signal_6746), .Z1_f (new_AGEMA_signal_6747) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[107]), .A0_f (ciphertext_s0_f[107]), .A1_t (ciphertext_s1_t[107]), .A1_f (ciphertext_s1_f[107]), .B0_t (ciphertext_s0_t[105]), .B0_f (ciphertext_s0_f[105]), .B1_t (ciphertext_s1_t[105]), .B1_f (ciphertext_s1_f[105]), .Z0_t (SubBytesIns_Inst_Sbox_13_T5), .Z0_f (new_AGEMA_signal_6748), .Z1_t (new_AGEMA_signal_6749), .Z1_f (new_AGEMA_signal_6750) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T1), .A0_f (new_AGEMA_signal_6736), .A1_t (new_AGEMA_signal_6737), .A1_f (new_AGEMA_signal_6738), .B0_t (SubBytesIns_Inst_Sbox_13_T5), .B0_f (new_AGEMA_signal_6748), .B1_t (new_AGEMA_signal_6749), .B1_f (new_AGEMA_signal_6750), .Z0_t (SubBytesIns_Inst_Sbox_13_T6), .Z0_f (new_AGEMA_signal_7240), .Z1_t (new_AGEMA_signal_7241), .Z1_f (new_AGEMA_signal_7242) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[110]), .A0_f (ciphertext_s0_f[110]), .A1_t (ciphertext_s1_t[110]), .A1_f (ciphertext_s1_f[110]), .B0_t (ciphertext_s0_t[109]), .B0_f (ciphertext_s0_f[109]), .B1_t (ciphertext_s1_t[109]), .B1_f (ciphertext_s1_f[109]), .Z0_t (SubBytesIns_Inst_Sbox_13_T7), .Z0_f (new_AGEMA_signal_6751), .Z1_t (new_AGEMA_signal_6752), .Z1_f (new_AGEMA_signal_6753) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[104]), .A0_f (ciphertext_s0_f[104]), .A1_t (ciphertext_s1_t[104]), .A1_f (ciphertext_s1_f[104]), .B0_t (SubBytesIns_Inst_Sbox_13_T6), .B0_f (new_AGEMA_signal_7240), .B1_t (new_AGEMA_signal_7241), .B1_f (new_AGEMA_signal_7242), .Z0_t (SubBytesIns_Inst_Sbox_13_T8), .Z0_f (new_AGEMA_signal_7979), .Z1_t (new_AGEMA_signal_7980), .Z1_f (new_AGEMA_signal_7981) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[104]), .A0_f (ciphertext_s0_f[104]), .A1_t (ciphertext_s1_t[104]), .A1_f (ciphertext_s1_f[104]), .B0_t (SubBytesIns_Inst_Sbox_13_T7), .B0_f (new_AGEMA_signal_6751), .B1_t (new_AGEMA_signal_6752), .B1_f (new_AGEMA_signal_6753), .Z0_t (SubBytesIns_Inst_Sbox_13_T9), .Z0_f (new_AGEMA_signal_7243), .Z1_t (new_AGEMA_signal_7244), .Z1_f (new_AGEMA_signal_7245) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T6), .A0_f (new_AGEMA_signal_7240), .A1_t (new_AGEMA_signal_7241), .A1_f (new_AGEMA_signal_7242), .B0_t (SubBytesIns_Inst_Sbox_13_T7), .B0_f (new_AGEMA_signal_6751), .B1_t (new_AGEMA_signal_6752), .B1_f (new_AGEMA_signal_6753), .Z0_t (SubBytesIns_Inst_Sbox_13_T10), .Z0_f (new_AGEMA_signal_7982), .Z1_t (new_AGEMA_signal_7983), .Z1_f (new_AGEMA_signal_7984) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[110]), .A0_f (ciphertext_s0_f[110]), .A1_t (ciphertext_s1_t[110]), .A1_f (ciphertext_s1_f[110]), .B0_t (ciphertext_s0_t[106]), .B0_f (ciphertext_s0_f[106]), .B1_t (ciphertext_s1_t[106]), .B1_f (ciphertext_s1_f[106]), .Z0_t (SubBytesIns_Inst_Sbox_13_T11), .Z0_f (new_AGEMA_signal_6754), .Z1_t (new_AGEMA_signal_6755), .Z1_f (new_AGEMA_signal_6756) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[109]), .A0_f (ciphertext_s0_f[109]), .A1_t (ciphertext_s1_t[109]), .A1_f (ciphertext_s1_f[109]), .B0_t (ciphertext_s0_t[106]), .B0_f (ciphertext_s0_f[106]), .B1_t (ciphertext_s1_t[106]), .B1_f (ciphertext_s1_f[106]), .Z0_t (SubBytesIns_Inst_Sbox_13_T12), .Z0_f (new_AGEMA_signal_6757), .Z1_t (new_AGEMA_signal_6758), .Z1_f (new_AGEMA_signal_6759) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T3), .A0_f (new_AGEMA_signal_6742), .A1_t (new_AGEMA_signal_6743), .A1_f (new_AGEMA_signal_6744), .B0_t (SubBytesIns_Inst_Sbox_13_T4), .B0_f (new_AGEMA_signal_6745), .B1_t (new_AGEMA_signal_6746), .B1_f (new_AGEMA_signal_6747), .Z0_t (SubBytesIns_Inst_Sbox_13_T13), .Z0_f (new_AGEMA_signal_7246), .Z1_t (new_AGEMA_signal_7247), .Z1_f (new_AGEMA_signal_7248) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T6), .A0_f (new_AGEMA_signal_7240), .A1_t (new_AGEMA_signal_7241), .A1_f (new_AGEMA_signal_7242), .B0_t (SubBytesIns_Inst_Sbox_13_T11), .B0_f (new_AGEMA_signal_6754), .B1_t (new_AGEMA_signal_6755), .B1_f (new_AGEMA_signal_6756), .Z0_t (SubBytesIns_Inst_Sbox_13_T14), .Z0_f (new_AGEMA_signal_7985), .Z1_t (new_AGEMA_signal_7986), .Z1_f (new_AGEMA_signal_7987) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T5), .A0_f (new_AGEMA_signal_6748), .A1_t (new_AGEMA_signal_6749), .A1_f (new_AGEMA_signal_6750), .B0_t (SubBytesIns_Inst_Sbox_13_T11), .B0_f (new_AGEMA_signal_6754), .B1_t (new_AGEMA_signal_6755), .B1_f (new_AGEMA_signal_6756), .Z0_t (SubBytesIns_Inst_Sbox_13_T15), .Z0_f (new_AGEMA_signal_7249), .Z1_t (new_AGEMA_signal_7250), .Z1_f (new_AGEMA_signal_7251) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T5), .A0_f (new_AGEMA_signal_6748), .A1_t (new_AGEMA_signal_6749), .A1_f (new_AGEMA_signal_6750), .B0_t (SubBytesIns_Inst_Sbox_13_T12), .B0_f (new_AGEMA_signal_6757), .B1_t (new_AGEMA_signal_6758), .B1_f (new_AGEMA_signal_6759), .Z0_t (SubBytesIns_Inst_Sbox_13_T16), .Z0_f (new_AGEMA_signal_7252), .Z1_t (new_AGEMA_signal_7253), .Z1_f (new_AGEMA_signal_7254) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T9), .A0_f (new_AGEMA_signal_7243), .A1_t (new_AGEMA_signal_7244), .A1_f (new_AGEMA_signal_7245), .B0_t (SubBytesIns_Inst_Sbox_13_T16), .B0_f (new_AGEMA_signal_7252), .B1_t (new_AGEMA_signal_7253), .B1_f (new_AGEMA_signal_7254), .Z0_t (SubBytesIns_Inst_Sbox_13_T17), .Z0_f (new_AGEMA_signal_7988), .Z1_t (new_AGEMA_signal_7989), .Z1_f (new_AGEMA_signal_7990) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[108]), .A0_f (ciphertext_s0_f[108]), .A1_t (ciphertext_s1_t[108]), .A1_f (ciphertext_s1_f[108]), .B0_t (ciphertext_s0_t[104]), .B0_f (ciphertext_s0_f[104]), .B1_t (ciphertext_s1_t[104]), .B1_f (ciphertext_s1_f[104]), .Z0_t (SubBytesIns_Inst_Sbox_13_T18), .Z0_f (new_AGEMA_signal_6760), .Z1_t (new_AGEMA_signal_6761), .Z1_f (new_AGEMA_signal_6762) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T7), .A0_f (new_AGEMA_signal_6751), .A1_t (new_AGEMA_signal_6752), .A1_f (new_AGEMA_signal_6753), .B0_t (SubBytesIns_Inst_Sbox_13_T18), .B0_f (new_AGEMA_signal_6760), .B1_t (new_AGEMA_signal_6761), .B1_f (new_AGEMA_signal_6762), .Z0_t (SubBytesIns_Inst_Sbox_13_T19), .Z0_f (new_AGEMA_signal_7255), .Z1_t (new_AGEMA_signal_7256), .Z1_f (new_AGEMA_signal_7257) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T1), .A0_f (new_AGEMA_signal_6736), .A1_t (new_AGEMA_signal_6737), .A1_f (new_AGEMA_signal_6738), .B0_t (SubBytesIns_Inst_Sbox_13_T19), .B0_f (new_AGEMA_signal_7255), .B1_t (new_AGEMA_signal_7256), .B1_f (new_AGEMA_signal_7257), .Z0_t (SubBytesIns_Inst_Sbox_13_T20), .Z0_f (new_AGEMA_signal_7991), .Z1_t (new_AGEMA_signal_7992), .Z1_f (new_AGEMA_signal_7993) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[105]), .A0_f (ciphertext_s0_f[105]), .A1_t (ciphertext_s1_t[105]), .A1_f (ciphertext_s1_f[105]), .B0_t (ciphertext_s0_t[104]), .B0_f (ciphertext_s0_f[104]), .B1_t (ciphertext_s1_t[104]), .B1_f (ciphertext_s1_f[104]), .Z0_t (SubBytesIns_Inst_Sbox_13_T21), .Z0_f (new_AGEMA_signal_6763), .Z1_t (new_AGEMA_signal_6764), .Z1_f (new_AGEMA_signal_6765) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T7), .A0_f (new_AGEMA_signal_6751), .A1_t (new_AGEMA_signal_6752), .A1_f (new_AGEMA_signal_6753), .B0_t (SubBytesIns_Inst_Sbox_13_T21), .B0_f (new_AGEMA_signal_6763), .B1_t (new_AGEMA_signal_6764), .B1_f (new_AGEMA_signal_6765), .Z0_t (SubBytesIns_Inst_Sbox_13_T22), .Z0_f (new_AGEMA_signal_7258), .Z1_t (new_AGEMA_signal_7259), .Z1_f (new_AGEMA_signal_7260) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T2), .A0_f (new_AGEMA_signal_6739), .A1_t (new_AGEMA_signal_6740), .A1_f (new_AGEMA_signal_6741), .B0_t (SubBytesIns_Inst_Sbox_13_T22), .B0_f (new_AGEMA_signal_7258), .B1_t (new_AGEMA_signal_7259), .B1_f (new_AGEMA_signal_7260), .Z0_t (SubBytesIns_Inst_Sbox_13_T23), .Z0_f (new_AGEMA_signal_7994), .Z1_t (new_AGEMA_signal_7995), .Z1_f (new_AGEMA_signal_7996) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T2), .A0_f (new_AGEMA_signal_6739), .A1_t (new_AGEMA_signal_6740), .A1_f (new_AGEMA_signal_6741), .B0_t (SubBytesIns_Inst_Sbox_13_T10), .B0_f (new_AGEMA_signal_7982), .B1_t (new_AGEMA_signal_7983), .B1_f (new_AGEMA_signal_7984), .Z0_t (SubBytesIns_Inst_Sbox_13_T24), .Z0_f (new_AGEMA_signal_8555), .Z1_t (new_AGEMA_signal_8556), .Z1_f (new_AGEMA_signal_8557) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T20), .A0_f (new_AGEMA_signal_7991), .A1_t (new_AGEMA_signal_7992), .A1_f (new_AGEMA_signal_7993), .B0_t (SubBytesIns_Inst_Sbox_13_T17), .B0_f (new_AGEMA_signal_7988), .B1_t (new_AGEMA_signal_7989), .B1_f (new_AGEMA_signal_7990), .Z0_t (SubBytesIns_Inst_Sbox_13_T25), .Z0_f (new_AGEMA_signal_8558), .Z1_t (new_AGEMA_signal_8559), .Z1_f (new_AGEMA_signal_8560) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T3), .A0_f (new_AGEMA_signal_6742), .A1_t (new_AGEMA_signal_6743), .A1_f (new_AGEMA_signal_6744), .B0_t (SubBytesIns_Inst_Sbox_13_T16), .B0_f (new_AGEMA_signal_7252), .B1_t (new_AGEMA_signal_7253), .B1_f (new_AGEMA_signal_7254), .Z0_t (SubBytesIns_Inst_Sbox_13_T26), .Z0_f (new_AGEMA_signal_7997), .Z1_t (new_AGEMA_signal_7998), .Z1_f (new_AGEMA_signal_7999) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T1), .A0_f (new_AGEMA_signal_6736), .A1_t (new_AGEMA_signal_6737), .A1_f (new_AGEMA_signal_6738), .B0_t (SubBytesIns_Inst_Sbox_13_T12), .B0_f (new_AGEMA_signal_6757), .B1_t (new_AGEMA_signal_6758), .B1_f (new_AGEMA_signal_6759), .Z0_t (SubBytesIns_Inst_Sbox_13_T27), .Z0_f (new_AGEMA_signal_7261), .Z1_t (new_AGEMA_signal_7262), .Z1_f (new_AGEMA_signal_7263) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T13), .A0_f (new_AGEMA_signal_7246), .A1_t (new_AGEMA_signal_7247), .A1_f (new_AGEMA_signal_7248), .B0_t (SubBytesIns_Inst_Sbox_13_T6), .B0_f (new_AGEMA_signal_7240), .B1_t (new_AGEMA_signal_7241), .B1_f (new_AGEMA_signal_7242), .Z0_t (SubBytesIns_Inst_Sbox_13_M1), .Z0_f (new_AGEMA_signal_8000), .Z1_t (new_AGEMA_signal_8001), .Z1_f (new_AGEMA_signal_8002) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T23), .A0_f (new_AGEMA_signal_7994), .A1_t (new_AGEMA_signal_7995), .A1_f (new_AGEMA_signal_7996), .B0_t (SubBytesIns_Inst_Sbox_13_T8), .B0_f (new_AGEMA_signal_7979), .B1_t (new_AGEMA_signal_7980), .B1_f (new_AGEMA_signal_7981), .Z0_t (SubBytesIns_Inst_Sbox_13_M2), .Z0_f (new_AGEMA_signal_8561), .Z1_t (new_AGEMA_signal_8562), .Z1_f (new_AGEMA_signal_8563) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T14), .A0_f (new_AGEMA_signal_7985), .A1_t (new_AGEMA_signal_7986), .A1_f (new_AGEMA_signal_7987), .B0_t (SubBytesIns_Inst_Sbox_13_M1), .B0_f (new_AGEMA_signal_8000), .B1_t (new_AGEMA_signal_8001), .B1_f (new_AGEMA_signal_8002), .Z0_t (SubBytesIns_Inst_Sbox_13_M3), .Z0_f (new_AGEMA_signal_8564), .Z1_t (new_AGEMA_signal_8565), .Z1_f (new_AGEMA_signal_8566) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T19), .A0_f (new_AGEMA_signal_7255), .A1_t (new_AGEMA_signal_7256), .A1_f (new_AGEMA_signal_7257), .B0_t (ciphertext_s0_t[104]), .B0_f (ciphertext_s0_f[104]), .B1_t (ciphertext_s1_t[104]), .B1_f (ciphertext_s1_f[104]), .Z0_t (SubBytesIns_Inst_Sbox_13_M4), .Z0_f (new_AGEMA_signal_8003), .Z1_t (new_AGEMA_signal_8004), .Z1_f (new_AGEMA_signal_8005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M4), .A0_f (new_AGEMA_signal_8003), .A1_t (new_AGEMA_signal_8004), .A1_f (new_AGEMA_signal_8005), .B0_t (SubBytesIns_Inst_Sbox_13_M1), .B0_f (new_AGEMA_signal_8000), .B1_t (new_AGEMA_signal_8001), .B1_f (new_AGEMA_signal_8002), .Z0_t (SubBytesIns_Inst_Sbox_13_M5), .Z0_f (new_AGEMA_signal_8567), .Z1_t (new_AGEMA_signal_8568), .Z1_f (new_AGEMA_signal_8569) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T3), .A0_f (new_AGEMA_signal_6742), .A1_t (new_AGEMA_signal_6743), .A1_f (new_AGEMA_signal_6744), .B0_t (SubBytesIns_Inst_Sbox_13_T16), .B0_f (new_AGEMA_signal_7252), .B1_t (new_AGEMA_signal_7253), .B1_f (new_AGEMA_signal_7254), .Z0_t (SubBytesIns_Inst_Sbox_13_M6), .Z0_f (new_AGEMA_signal_8006), .Z1_t (new_AGEMA_signal_8007), .Z1_f (new_AGEMA_signal_8008) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T22), .A0_f (new_AGEMA_signal_7258), .A1_t (new_AGEMA_signal_7259), .A1_f (new_AGEMA_signal_7260), .B0_t (SubBytesIns_Inst_Sbox_13_T9), .B0_f (new_AGEMA_signal_7243), .B1_t (new_AGEMA_signal_7244), .B1_f (new_AGEMA_signal_7245), .Z0_t (SubBytesIns_Inst_Sbox_13_M7), .Z0_f (new_AGEMA_signal_8009), .Z1_t (new_AGEMA_signal_8010), .Z1_f (new_AGEMA_signal_8011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T26), .A0_f (new_AGEMA_signal_7997), .A1_t (new_AGEMA_signal_7998), .A1_f (new_AGEMA_signal_7999), .B0_t (SubBytesIns_Inst_Sbox_13_M6), .B0_f (new_AGEMA_signal_8006), .B1_t (new_AGEMA_signal_8007), .B1_f (new_AGEMA_signal_8008), .Z0_t (SubBytesIns_Inst_Sbox_13_M8), .Z0_f (new_AGEMA_signal_8570), .Z1_t (new_AGEMA_signal_8571), .Z1_f (new_AGEMA_signal_8572) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T20), .A0_f (new_AGEMA_signal_7991), .A1_t (new_AGEMA_signal_7992), .A1_f (new_AGEMA_signal_7993), .B0_t (SubBytesIns_Inst_Sbox_13_T17), .B0_f (new_AGEMA_signal_7988), .B1_t (new_AGEMA_signal_7989), .B1_f (new_AGEMA_signal_7990), .Z0_t (SubBytesIns_Inst_Sbox_13_M9), .Z0_f (new_AGEMA_signal_8573), .Z1_t (new_AGEMA_signal_8574), .Z1_f (new_AGEMA_signal_8575) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M9), .A0_f (new_AGEMA_signal_8573), .A1_t (new_AGEMA_signal_8574), .A1_f (new_AGEMA_signal_8575), .B0_t (SubBytesIns_Inst_Sbox_13_M6), .B0_f (new_AGEMA_signal_8006), .B1_t (new_AGEMA_signal_8007), .B1_f (new_AGEMA_signal_8008), .Z0_t (SubBytesIns_Inst_Sbox_13_M10), .Z0_f (new_AGEMA_signal_8891), .Z1_t (new_AGEMA_signal_8892), .Z1_f (new_AGEMA_signal_8893) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T1), .A0_f (new_AGEMA_signal_6736), .A1_t (new_AGEMA_signal_6737), .A1_f (new_AGEMA_signal_6738), .B0_t (SubBytesIns_Inst_Sbox_13_T15), .B0_f (new_AGEMA_signal_7249), .B1_t (new_AGEMA_signal_7250), .B1_f (new_AGEMA_signal_7251), .Z0_t (SubBytesIns_Inst_Sbox_13_M11), .Z0_f (new_AGEMA_signal_8012), .Z1_t (new_AGEMA_signal_8013), .Z1_f (new_AGEMA_signal_8014) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T4), .A0_f (new_AGEMA_signal_6745), .A1_t (new_AGEMA_signal_6746), .A1_f (new_AGEMA_signal_6747), .B0_t (SubBytesIns_Inst_Sbox_13_T27), .B0_f (new_AGEMA_signal_7261), .B1_t (new_AGEMA_signal_7262), .B1_f (new_AGEMA_signal_7263), .Z0_t (SubBytesIns_Inst_Sbox_13_M12), .Z0_f (new_AGEMA_signal_8015), .Z1_t (new_AGEMA_signal_8016), .Z1_f (new_AGEMA_signal_8017) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M12), .A0_f (new_AGEMA_signal_8015), .A1_t (new_AGEMA_signal_8016), .A1_f (new_AGEMA_signal_8017), .B0_t (SubBytesIns_Inst_Sbox_13_M11), .B0_f (new_AGEMA_signal_8012), .B1_t (new_AGEMA_signal_8013), .B1_f (new_AGEMA_signal_8014), .Z0_t (SubBytesIns_Inst_Sbox_13_M13), .Z0_f (new_AGEMA_signal_8576), .Z1_t (new_AGEMA_signal_8577), .Z1_f (new_AGEMA_signal_8578) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T2), .A0_f (new_AGEMA_signal_6739), .A1_t (new_AGEMA_signal_6740), .A1_f (new_AGEMA_signal_6741), .B0_t (SubBytesIns_Inst_Sbox_13_T10), .B0_f (new_AGEMA_signal_7982), .B1_t (new_AGEMA_signal_7983), .B1_f (new_AGEMA_signal_7984), .Z0_t (SubBytesIns_Inst_Sbox_13_M14), .Z0_f (new_AGEMA_signal_8579), .Z1_t (new_AGEMA_signal_8580), .Z1_f (new_AGEMA_signal_8581) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M14), .A0_f (new_AGEMA_signal_8579), .A1_t (new_AGEMA_signal_8580), .A1_f (new_AGEMA_signal_8581), .B0_t (SubBytesIns_Inst_Sbox_13_M11), .B0_f (new_AGEMA_signal_8012), .B1_t (new_AGEMA_signal_8013), .B1_f (new_AGEMA_signal_8014), .Z0_t (SubBytesIns_Inst_Sbox_13_M15), .Z0_f (new_AGEMA_signal_8894), .Z1_t (new_AGEMA_signal_8895), .Z1_f (new_AGEMA_signal_8896) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M3), .A0_f (new_AGEMA_signal_8564), .A1_t (new_AGEMA_signal_8565), .A1_f (new_AGEMA_signal_8566), .B0_t (SubBytesIns_Inst_Sbox_13_M2), .B0_f (new_AGEMA_signal_8561), .B1_t (new_AGEMA_signal_8562), .B1_f (new_AGEMA_signal_8563), .Z0_t (SubBytesIns_Inst_Sbox_13_M16), .Z0_f (new_AGEMA_signal_8897), .Z1_t (new_AGEMA_signal_8898), .Z1_f (new_AGEMA_signal_8899) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M5), .A0_f (new_AGEMA_signal_8567), .A1_t (new_AGEMA_signal_8568), .A1_f (new_AGEMA_signal_8569), .B0_t (SubBytesIns_Inst_Sbox_13_T24), .B0_f (new_AGEMA_signal_8555), .B1_t (new_AGEMA_signal_8556), .B1_f (new_AGEMA_signal_8557), .Z0_t (SubBytesIns_Inst_Sbox_13_M17), .Z0_f (new_AGEMA_signal_8900), .Z1_t (new_AGEMA_signal_8901), .Z1_f (new_AGEMA_signal_8902) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M8), .A0_f (new_AGEMA_signal_8570), .A1_t (new_AGEMA_signal_8571), .A1_f (new_AGEMA_signal_8572), .B0_t (SubBytesIns_Inst_Sbox_13_M7), .B0_f (new_AGEMA_signal_8009), .B1_t (new_AGEMA_signal_8010), .B1_f (new_AGEMA_signal_8011), .Z0_t (SubBytesIns_Inst_Sbox_13_M18), .Z0_f (new_AGEMA_signal_8903), .Z1_t (new_AGEMA_signal_8904), .Z1_f (new_AGEMA_signal_8905) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M10), .A0_f (new_AGEMA_signal_8891), .A1_t (new_AGEMA_signal_8892), .A1_f (new_AGEMA_signal_8893), .B0_t (SubBytesIns_Inst_Sbox_13_M15), .B0_f (new_AGEMA_signal_8894), .B1_t (new_AGEMA_signal_8895), .B1_f (new_AGEMA_signal_8896), .Z0_t (SubBytesIns_Inst_Sbox_13_M19), .Z0_f (new_AGEMA_signal_9140), .Z1_t (new_AGEMA_signal_9141), .Z1_f (new_AGEMA_signal_9142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M16), .A0_f (new_AGEMA_signal_8897), .A1_t (new_AGEMA_signal_8898), .A1_f (new_AGEMA_signal_8899), .B0_t (SubBytesIns_Inst_Sbox_13_M13), .B0_f (new_AGEMA_signal_8576), .B1_t (new_AGEMA_signal_8577), .B1_f (new_AGEMA_signal_8578), .Z0_t (SubBytesIns_Inst_Sbox_13_M20), .Z0_f (new_AGEMA_signal_9143), .Z1_t (new_AGEMA_signal_9144), .Z1_f (new_AGEMA_signal_9145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M17), .A0_f (new_AGEMA_signal_8900), .A1_t (new_AGEMA_signal_8901), .A1_f (new_AGEMA_signal_8902), .B0_t (SubBytesIns_Inst_Sbox_13_M15), .B0_f (new_AGEMA_signal_8894), .B1_t (new_AGEMA_signal_8895), .B1_f (new_AGEMA_signal_8896), .Z0_t (SubBytesIns_Inst_Sbox_13_M21), .Z0_f (new_AGEMA_signal_9146), .Z1_t (new_AGEMA_signal_9147), .Z1_f (new_AGEMA_signal_9148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M18), .A0_f (new_AGEMA_signal_8903), .A1_t (new_AGEMA_signal_8904), .A1_f (new_AGEMA_signal_8905), .B0_t (SubBytesIns_Inst_Sbox_13_M13), .B0_f (new_AGEMA_signal_8576), .B1_t (new_AGEMA_signal_8577), .B1_f (new_AGEMA_signal_8578), .Z0_t (SubBytesIns_Inst_Sbox_13_M22), .Z0_f (new_AGEMA_signal_9149), .Z1_t (new_AGEMA_signal_9150), .Z1_f (new_AGEMA_signal_9151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M19), .A0_f (new_AGEMA_signal_9140), .A1_t (new_AGEMA_signal_9141), .A1_f (new_AGEMA_signal_9142), .B0_t (SubBytesIns_Inst_Sbox_13_T25), .B0_f (new_AGEMA_signal_8558), .B1_t (new_AGEMA_signal_8559), .B1_f (new_AGEMA_signal_8560), .Z0_t (SubBytesIns_Inst_Sbox_13_M23), .Z0_f (new_AGEMA_signal_9380), .Z1_t (new_AGEMA_signal_9381), .Z1_f (new_AGEMA_signal_9382) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M22), .A0_f (new_AGEMA_signal_9149), .A1_t (new_AGEMA_signal_9150), .A1_f (new_AGEMA_signal_9151), .B0_t (SubBytesIns_Inst_Sbox_13_M23), .B0_f (new_AGEMA_signal_9380), .B1_t (new_AGEMA_signal_9381), .B1_f (new_AGEMA_signal_9382), .Z0_t (SubBytesIns_Inst_Sbox_13_M24), .Z0_f (new_AGEMA_signal_9671), .Z1_t (new_AGEMA_signal_9672), .Z1_f (new_AGEMA_signal_9673) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M22), .A0_f (new_AGEMA_signal_9149), .A1_t (new_AGEMA_signal_9150), .A1_f (new_AGEMA_signal_9151), .B0_t (SubBytesIns_Inst_Sbox_13_M20), .B0_f (new_AGEMA_signal_9143), .B1_t (new_AGEMA_signal_9144), .B1_f (new_AGEMA_signal_9145), .Z0_t (SubBytesIns_Inst_Sbox_13_M25), .Z0_f (new_AGEMA_signal_9383), .Z1_t (new_AGEMA_signal_9384), .Z1_f (new_AGEMA_signal_9385) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M21), .A0_f (new_AGEMA_signal_9146), .A1_t (new_AGEMA_signal_9147), .A1_f (new_AGEMA_signal_9148), .B0_t (SubBytesIns_Inst_Sbox_13_M25), .B0_f (new_AGEMA_signal_9383), .B1_t (new_AGEMA_signal_9384), .B1_f (new_AGEMA_signal_9385), .Z0_t (SubBytesIns_Inst_Sbox_13_M26), .Z0_f (new_AGEMA_signal_9674), .Z1_t (new_AGEMA_signal_9675), .Z1_f (new_AGEMA_signal_9676) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M20), .A0_f (new_AGEMA_signal_9143), .A1_t (new_AGEMA_signal_9144), .A1_f (new_AGEMA_signal_9145), .B0_t (SubBytesIns_Inst_Sbox_13_M21), .B0_f (new_AGEMA_signal_9146), .B1_t (new_AGEMA_signal_9147), .B1_f (new_AGEMA_signal_9148), .Z0_t (SubBytesIns_Inst_Sbox_13_M27), .Z0_f (new_AGEMA_signal_9386), .Z1_t (new_AGEMA_signal_9387), .Z1_f (new_AGEMA_signal_9388) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M23), .A0_f (new_AGEMA_signal_9380), .A1_t (new_AGEMA_signal_9381), .A1_f (new_AGEMA_signal_9382), .B0_t (SubBytesIns_Inst_Sbox_13_M25), .B0_f (new_AGEMA_signal_9383), .B1_t (new_AGEMA_signal_9384), .B1_f (new_AGEMA_signal_9385), .Z0_t (SubBytesIns_Inst_Sbox_13_M28), .Z0_f (new_AGEMA_signal_9677), .Z1_t (new_AGEMA_signal_9678), .Z1_f (new_AGEMA_signal_9679) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M28), .A0_f (new_AGEMA_signal_9677), .A1_t (new_AGEMA_signal_9678), .A1_f (new_AGEMA_signal_9679), .B0_t (SubBytesIns_Inst_Sbox_13_M27), .B0_f (new_AGEMA_signal_9386), .B1_t (new_AGEMA_signal_9387), .B1_f (new_AGEMA_signal_9388), .Z0_t (SubBytesIns_Inst_Sbox_13_M29), .Z0_f (new_AGEMA_signal_9971), .Z1_t (new_AGEMA_signal_9972), .Z1_f (new_AGEMA_signal_9973) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M26), .A0_f (new_AGEMA_signal_9674), .A1_t (new_AGEMA_signal_9675), .A1_f (new_AGEMA_signal_9676), .B0_t (SubBytesIns_Inst_Sbox_13_M24), .B0_f (new_AGEMA_signal_9671), .B1_t (new_AGEMA_signal_9672), .B1_f (new_AGEMA_signal_9673), .Z0_t (SubBytesIns_Inst_Sbox_13_M30), .Z0_f (new_AGEMA_signal_9974), .Z1_t (new_AGEMA_signal_9975), .Z1_f (new_AGEMA_signal_9976) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M20), .A0_f (new_AGEMA_signal_9143), .A1_t (new_AGEMA_signal_9144), .A1_f (new_AGEMA_signal_9145), .B0_t (SubBytesIns_Inst_Sbox_13_M23), .B0_f (new_AGEMA_signal_9380), .B1_t (new_AGEMA_signal_9381), .B1_f (new_AGEMA_signal_9382), .Z0_t (SubBytesIns_Inst_Sbox_13_M31), .Z0_f (new_AGEMA_signal_9680), .Z1_t (new_AGEMA_signal_9681), .Z1_f (new_AGEMA_signal_9682) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M27), .A0_f (new_AGEMA_signal_9386), .A1_t (new_AGEMA_signal_9387), .A1_f (new_AGEMA_signal_9388), .B0_t (SubBytesIns_Inst_Sbox_13_M31), .B0_f (new_AGEMA_signal_9680), .B1_t (new_AGEMA_signal_9681), .B1_f (new_AGEMA_signal_9682), .Z0_t (SubBytesIns_Inst_Sbox_13_M32), .Z0_f (new_AGEMA_signal_9977), .Z1_t (new_AGEMA_signal_9978), .Z1_f (new_AGEMA_signal_9979) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M27), .A0_f (new_AGEMA_signal_9386), .A1_t (new_AGEMA_signal_9387), .A1_f (new_AGEMA_signal_9388), .B0_t (SubBytesIns_Inst_Sbox_13_M25), .B0_f (new_AGEMA_signal_9383), .B1_t (new_AGEMA_signal_9384), .B1_f (new_AGEMA_signal_9385), .Z0_t (SubBytesIns_Inst_Sbox_13_M33), .Z0_f (new_AGEMA_signal_9683), .Z1_t (new_AGEMA_signal_9684), .Z1_f (new_AGEMA_signal_9685) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M21), .A0_f (new_AGEMA_signal_9146), .A1_t (new_AGEMA_signal_9147), .A1_f (new_AGEMA_signal_9148), .B0_t (SubBytesIns_Inst_Sbox_13_M22), .B0_f (new_AGEMA_signal_9149), .B1_t (new_AGEMA_signal_9150), .B1_f (new_AGEMA_signal_9151), .Z0_t (SubBytesIns_Inst_Sbox_13_M34), .Z0_f (new_AGEMA_signal_9389), .Z1_t (new_AGEMA_signal_9390), .Z1_f (new_AGEMA_signal_9391) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M24), .A0_f (new_AGEMA_signal_9671), .A1_t (new_AGEMA_signal_9672), .A1_f (new_AGEMA_signal_9673), .B0_t (SubBytesIns_Inst_Sbox_13_M34), .B0_f (new_AGEMA_signal_9389), .B1_t (new_AGEMA_signal_9390), .B1_f (new_AGEMA_signal_9391), .Z0_t (SubBytesIns_Inst_Sbox_13_M35), .Z0_f (new_AGEMA_signal_9980), .Z1_t (new_AGEMA_signal_9981), .Z1_f (new_AGEMA_signal_9982) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M24), .A0_f (new_AGEMA_signal_9671), .A1_t (new_AGEMA_signal_9672), .A1_f (new_AGEMA_signal_9673), .B0_t (SubBytesIns_Inst_Sbox_13_M25), .B0_f (new_AGEMA_signal_9383), .B1_t (new_AGEMA_signal_9384), .B1_f (new_AGEMA_signal_9385), .Z0_t (SubBytesIns_Inst_Sbox_13_M36), .Z0_f (new_AGEMA_signal_9983), .Z1_t (new_AGEMA_signal_9984), .Z1_f (new_AGEMA_signal_9985) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M21), .A0_f (new_AGEMA_signal_9146), .A1_t (new_AGEMA_signal_9147), .A1_f (new_AGEMA_signal_9148), .B0_t (SubBytesIns_Inst_Sbox_13_M29), .B0_f (new_AGEMA_signal_9971), .B1_t (new_AGEMA_signal_9972), .B1_f (new_AGEMA_signal_9973), .Z0_t (SubBytesIns_Inst_Sbox_13_M37), .Z0_f (new_AGEMA_signal_10220), .Z1_t (new_AGEMA_signal_10221), .Z1_f (new_AGEMA_signal_10222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M32), .A0_f (new_AGEMA_signal_9977), .A1_t (new_AGEMA_signal_9978), .A1_f (new_AGEMA_signal_9979), .B0_t (SubBytesIns_Inst_Sbox_13_M33), .B0_f (new_AGEMA_signal_9683), .B1_t (new_AGEMA_signal_9684), .B1_f (new_AGEMA_signal_9685), .Z0_t (SubBytesIns_Inst_Sbox_13_M38), .Z0_f (new_AGEMA_signal_10223), .Z1_t (new_AGEMA_signal_10224), .Z1_f (new_AGEMA_signal_10225) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M23), .A0_f (new_AGEMA_signal_9380), .A1_t (new_AGEMA_signal_9381), .A1_f (new_AGEMA_signal_9382), .B0_t (SubBytesIns_Inst_Sbox_13_M30), .B0_f (new_AGEMA_signal_9974), .B1_t (new_AGEMA_signal_9975), .B1_f (new_AGEMA_signal_9976), .Z0_t (SubBytesIns_Inst_Sbox_13_M39), .Z0_f (new_AGEMA_signal_10226), .Z1_t (new_AGEMA_signal_10227), .Z1_f (new_AGEMA_signal_10228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M35), .A0_f (new_AGEMA_signal_9980), .A1_t (new_AGEMA_signal_9981), .A1_f (new_AGEMA_signal_9982), .B0_t (SubBytesIns_Inst_Sbox_13_M36), .B0_f (new_AGEMA_signal_9983), .B1_t (new_AGEMA_signal_9984), .B1_f (new_AGEMA_signal_9985), .Z0_t (SubBytesIns_Inst_Sbox_13_M40), .Z0_f (new_AGEMA_signal_10229), .Z1_t (new_AGEMA_signal_10230), .Z1_f (new_AGEMA_signal_10231) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M38), .A0_f (new_AGEMA_signal_10223), .A1_t (new_AGEMA_signal_10224), .A1_f (new_AGEMA_signal_10225), .B0_t (SubBytesIns_Inst_Sbox_13_M40), .B0_f (new_AGEMA_signal_10229), .B1_t (new_AGEMA_signal_10230), .B1_f (new_AGEMA_signal_10231), .Z0_t (SubBytesIns_Inst_Sbox_13_M41), .Z0_f (new_AGEMA_signal_10868), .Z1_t (new_AGEMA_signal_10869), .Z1_f (new_AGEMA_signal_10870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M37), .A0_f (new_AGEMA_signal_10220), .A1_t (new_AGEMA_signal_10221), .A1_f (new_AGEMA_signal_10222), .B0_t (SubBytesIns_Inst_Sbox_13_M39), .B0_f (new_AGEMA_signal_10226), .B1_t (new_AGEMA_signal_10227), .B1_f (new_AGEMA_signal_10228), .Z0_t (SubBytesIns_Inst_Sbox_13_M42), .Z0_f (new_AGEMA_signal_10871), .Z1_t (new_AGEMA_signal_10872), .Z1_f (new_AGEMA_signal_10873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M37), .A0_f (new_AGEMA_signal_10220), .A1_t (new_AGEMA_signal_10221), .A1_f (new_AGEMA_signal_10222), .B0_t (SubBytesIns_Inst_Sbox_13_M38), .B0_f (new_AGEMA_signal_10223), .B1_t (new_AGEMA_signal_10224), .B1_f (new_AGEMA_signal_10225), .Z0_t (SubBytesIns_Inst_Sbox_13_M43), .Z0_f (new_AGEMA_signal_10874), .Z1_t (new_AGEMA_signal_10875), .Z1_f (new_AGEMA_signal_10876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M39), .A0_f (new_AGEMA_signal_10226), .A1_t (new_AGEMA_signal_10227), .A1_f (new_AGEMA_signal_10228), .B0_t (SubBytesIns_Inst_Sbox_13_M40), .B0_f (new_AGEMA_signal_10229), .B1_t (new_AGEMA_signal_10230), .B1_f (new_AGEMA_signal_10231), .Z0_t (SubBytesIns_Inst_Sbox_13_M44), .Z0_f (new_AGEMA_signal_10877), .Z1_t (new_AGEMA_signal_10878), .Z1_f (new_AGEMA_signal_10879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M42), .A0_f (new_AGEMA_signal_10871), .A1_t (new_AGEMA_signal_10872), .A1_f (new_AGEMA_signal_10873), .B0_t (SubBytesIns_Inst_Sbox_13_M41), .B0_f (new_AGEMA_signal_10868), .B1_t (new_AGEMA_signal_10869), .B1_f (new_AGEMA_signal_10870), .Z0_t (SubBytesIns_Inst_Sbox_13_M45), .Z0_f (new_AGEMA_signal_11588), .Z1_t (new_AGEMA_signal_11589), .Z1_f (new_AGEMA_signal_11590) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M44), .A0_f (new_AGEMA_signal_10877), .A1_t (new_AGEMA_signal_10878), .A1_f (new_AGEMA_signal_10879), .B0_t (SubBytesIns_Inst_Sbox_13_T6), .B0_f (new_AGEMA_signal_7240), .B1_t (new_AGEMA_signal_7241), .B1_f (new_AGEMA_signal_7242), .Z0_t (SubBytesIns_Inst_Sbox_13_M46), .Z0_f (new_AGEMA_signal_11591), .Z1_t (new_AGEMA_signal_11592), .Z1_f (new_AGEMA_signal_11593) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M40), .A0_f (new_AGEMA_signal_10229), .A1_t (new_AGEMA_signal_10230), .A1_f (new_AGEMA_signal_10231), .B0_t (SubBytesIns_Inst_Sbox_13_T8), .B0_f (new_AGEMA_signal_7979), .B1_t (new_AGEMA_signal_7980), .B1_f (new_AGEMA_signal_7981), .Z0_t (SubBytesIns_Inst_Sbox_13_M47), .Z0_f (new_AGEMA_signal_10880), .Z1_t (new_AGEMA_signal_10881), .Z1_f (new_AGEMA_signal_10882) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M39), .A0_f (new_AGEMA_signal_10226), .A1_t (new_AGEMA_signal_10227), .A1_f (new_AGEMA_signal_10228), .B0_t (ciphertext_s0_t[104]), .B0_f (ciphertext_s0_f[104]), .B1_t (ciphertext_s1_t[104]), .B1_f (ciphertext_s1_f[104]), .Z0_t (SubBytesIns_Inst_Sbox_13_M48), .Z0_f (new_AGEMA_signal_10883), .Z1_t (new_AGEMA_signal_10884), .Z1_f (new_AGEMA_signal_10885) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M43), .A0_f (new_AGEMA_signal_10874), .A1_t (new_AGEMA_signal_10875), .A1_f (new_AGEMA_signal_10876), .B0_t (SubBytesIns_Inst_Sbox_13_T16), .B0_f (new_AGEMA_signal_7252), .B1_t (new_AGEMA_signal_7253), .B1_f (new_AGEMA_signal_7254), .Z0_t (SubBytesIns_Inst_Sbox_13_M49), .Z0_f (new_AGEMA_signal_11594), .Z1_t (new_AGEMA_signal_11595), .Z1_f (new_AGEMA_signal_11596) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M38), .A0_f (new_AGEMA_signal_10223), .A1_t (new_AGEMA_signal_10224), .A1_f (new_AGEMA_signal_10225), .B0_t (SubBytesIns_Inst_Sbox_13_T9), .B0_f (new_AGEMA_signal_7243), .B1_t (new_AGEMA_signal_7244), .B1_f (new_AGEMA_signal_7245), .Z0_t (SubBytesIns_Inst_Sbox_13_M50), .Z0_f (new_AGEMA_signal_10886), .Z1_t (new_AGEMA_signal_10887), .Z1_f (new_AGEMA_signal_10888) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M37), .A0_f (new_AGEMA_signal_10220), .A1_t (new_AGEMA_signal_10221), .A1_f (new_AGEMA_signal_10222), .B0_t (SubBytesIns_Inst_Sbox_13_T17), .B0_f (new_AGEMA_signal_7988), .B1_t (new_AGEMA_signal_7989), .B1_f (new_AGEMA_signal_7990), .Z0_t (SubBytesIns_Inst_Sbox_13_M51), .Z0_f (new_AGEMA_signal_10889), .Z1_t (new_AGEMA_signal_10890), .Z1_f (new_AGEMA_signal_10891) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M42), .A0_f (new_AGEMA_signal_10871), .A1_t (new_AGEMA_signal_10872), .A1_f (new_AGEMA_signal_10873), .B0_t (SubBytesIns_Inst_Sbox_13_T15), .B0_f (new_AGEMA_signal_7249), .B1_t (new_AGEMA_signal_7250), .B1_f (new_AGEMA_signal_7251), .Z0_t (SubBytesIns_Inst_Sbox_13_M52), .Z0_f (new_AGEMA_signal_11597), .Z1_t (new_AGEMA_signal_11598), .Z1_f (new_AGEMA_signal_11599) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M45), .A0_f (new_AGEMA_signal_11588), .A1_t (new_AGEMA_signal_11589), .A1_f (new_AGEMA_signal_11590), .B0_t (SubBytesIns_Inst_Sbox_13_T27), .B0_f (new_AGEMA_signal_7261), .B1_t (new_AGEMA_signal_7262), .B1_f (new_AGEMA_signal_7263), .Z0_t (SubBytesIns_Inst_Sbox_13_M53), .Z0_f (new_AGEMA_signal_12206), .Z1_t (new_AGEMA_signal_12207), .Z1_f (new_AGEMA_signal_12208) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M41), .A0_f (new_AGEMA_signal_10868), .A1_t (new_AGEMA_signal_10869), .A1_f (new_AGEMA_signal_10870), .B0_t (SubBytesIns_Inst_Sbox_13_T10), .B0_f (new_AGEMA_signal_7982), .B1_t (new_AGEMA_signal_7983), .B1_f (new_AGEMA_signal_7984), .Z0_t (SubBytesIns_Inst_Sbox_13_M54), .Z0_f (new_AGEMA_signal_11600), .Z1_t (new_AGEMA_signal_11601), .Z1_f (new_AGEMA_signal_11602) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M44), .A0_f (new_AGEMA_signal_10877), .A1_t (new_AGEMA_signal_10878), .A1_f (new_AGEMA_signal_10879), .B0_t (SubBytesIns_Inst_Sbox_13_T13), .B0_f (new_AGEMA_signal_7246), .B1_t (new_AGEMA_signal_7247), .B1_f (new_AGEMA_signal_7248), .Z0_t (SubBytesIns_Inst_Sbox_13_M55), .Z0_f (new_AGEMA_signal_11603), .Z1_t (new_AGEMA_signal_11604), .Z1_f (new_AGEMA_signal_11605) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M40), .A0_f (new_AGEMA_signal_10229), .A1_t (new_AGEMA_signal_10230), .A1_f (new_AGEMA_signal_10231), .B0_t (SubBytesIns_Inst_Sbox_13_T23), .B0_f (new_AGEMA_signal_7994), .B1_t (new_AGEMA_signal_7995), .B1_f (new_AGEMA_signal_7996), .Z0_t (SubBytesIns_Inst_Sbox_13_M56), .Z0_f (new_AGEMA_signal_10892), .Z1_t (new_AGEMA_signal_10893), .Z1_f (new_AGEMA_signal_10894) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M39), .A0_f (new_AGEMA_signal_10226), .A1_t (new_AGEMA_signal_10227), .A1_f (new_AGEMA_signal_10228), .B0_t (SubBytesIns_Inst_Sbox_13_T19), .B0_f (new_AGEMA_signal_7255), .B1_t (new_AGEMA_signal_7256), .B1_f (new_AGEMA_signal_7257), .Z0_t (SubBytesIns_Inst_Sbox_13_M57), .Z0_f (new_AGEMA_signal_10895), .Z1_t (new_AGEMA_signal_10896), .Z1_f (new_AGEMA_signal_10897) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M43), .A0_f (new_AGEMA_signal_10874), .A1_t (new_AGEMA_signal_10875), .A1_f (new_AGEMA_signal_10876), .B0_t (SubBytesIns_Inst_Sbox_13_T3), .B0_f (new_AGEMA_signal_6742), .B1_t (new_AGEMA_signal_6743), .B1_f (new_AGEMA_signal_6744), .Z0_t (SubBytesIns_Inst_Sbox_13_M58), .Z0_f (new_AGEMA_signal_11606), .Z1_t (new_AGEMA_signal_11607), .Z1_f (new_AGEMA_signal_11608) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M38), .A0_f (new_AGEMA_signal_10223), .A1_t (new_AGEMA_signal_10224), .A1_f (new_AGEMA_signal_10225), .B0_t (SubBytesIns_Inst_Sbox_13_T22), .B0_f (new_AGEMA_signal_7258), .B1_t (new_AGEMA_signal_7259), .B1_f (new_AGEMA_signal_7260), .Z0_t (SubBytesIns_Inst_Sbox_13_M59), .Z0_f (new_AGEMA_signal_10898), .Z1_t (new_AGEMA_signal_10899), .Z1_f (new_AGEMA_signal_10900) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M37), .A0_f (new_AGEMA_signal_10220), .A1_t (new_AGEMA_signal_10221), .A1_f (new_AGEMA_signal_10222), .B0_t (SubBytesIns_Inst_Sbox_13_T20), .B0_f (new_AGEMA_signal_7991), .B1_t (new_AGEMA_signal_7992), .B1_f (new_AGEMA_signal_7993), .Z0_t (SubBytesIns_Inst_Sbox_13_M60), .Z0_f (new_AGEMA_signal_10901), .Z1_t (new_AGEMA_signal_10902), .Z1_f (new_AGEMA_signal_10903) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M42), .A0_f (new_AGEMA_signal_10871), .A1_t (new_AGEMA_signal_10872), .A1_f (new_AGEMA_signal_10873), .B0_t (SubBytesIns_Inst_Sbox_13_T1), .B0_f (new_AGEMA_signal_6736), .B1_t (new_AGEMA_signal_6737), .B1_f (new_AGEMA_signal_6738), .Z0_t (SubBytesIns_Inst_Sbox_13_M61), .Z0_f (new_AGEMA_signal_11609), .Z1_t (new_AGEMA_signal_11610), .Z1_f (new_AGEMA_signal_11611) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M45), .A0_f (new_AGEMA_signal_11588), .A1_t (new_AGEMA_signal_11589), .A1_f (new_AGEMA_signal_11590), .B0_t (SubBytesIns_Inst_Sbox_13_T4), .B0_f (new_AGEMA_signal_6745), .B1_t (new_AGEMA_signal_6746), .B1_f (new_AGEMA_signal_6747), .Z0_t (SubBytesIns_Inst_Sbox_13_M62), .Z0_f (new_AGEMA_signal_12209), .Z1_t (new_AGEMA_signal_12210), .Z1_f (new_AGEMA_signal_12211) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M41), .A0_f (new_AGEMA_signal_10868), .A1_t (new_AGEMA_signal_10869), .A1_f (new_AGEMA_signal_10870), .B0_t (SubBytesIns_Inst_Sbox_13_T2), .B0_f (new_AGEMA_signal_6739), .B1_t (new_AGEMA_signal_6740), .B1_f (new_AGEMA_signal_6741), .Z0_t (SubBytesIns_Inst_Sbox_13_M63), .Z0_f (new_AGEMA_signal_11612), .Z1_t (new_AGEMA_signal_11613), .Z1_f (new_AGEMA_signal_11614) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M61), .A0_f (new_AGEMA_signal_11609), .A1_t (new_AGEMA_signal_11610), .A1_f (new_AGEMA_signal_11611), .B0_t (SubBytesIns_Inst_Sbox_13_M62), .B0_f (new_AGEMA_signal_12209), .B1_t (new_AGEMA_signal_12210), .B1_f (new_AGEMA_signal_12211), .Z0_t (SubBytesIns_Inst_Sbox_13_L0), .Z0_f (new_AGEMA_signal_12755), .Z1_t (new_AGEMA_signal_12756), .Z1_f (new_AGEMA_signal_12757) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M50), .A0_f (new_AGEMA_signal_10886), .A1_t (new_AGEMA_signal_10887), .A1_f (new_AGEMA_signal_10888), .B0_t (SubBytesIns_Inst_Sbox_13_M56), .B0_f (new_AGEMA_signal_10892), .B1_t (new_AGEMA_signal_10893), .B1_f (new_AGEMA_signal_10894), .Z0_t (SubBytesIns_Inst_Sbox_13_L1), .Z0_f (new_AGEMA_signal_11615), .Z1_t (new_AGEMA_signal_11616), .Z1_f (new_AGEMA_signal_11617) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M46), .A0_f (new_AGEMA_signal_11591), .A1_t (new_AGEMA_signal_11592), .A1_f (new_AGEMA_signal_11593), .B0_t (SubBytesIns_Inst_Sbox_13_M48), .B0_f (new_AGEMA_signal_10883), .B1_t (new_AGEMA_signal_10884), .B1_f (new_AGEMA_signal_10885), .Z0_t (SubBytesIns_Inst_Sbox_13_L2), .Z0_f (new_AGEMA_signal_12212), .Z1_t (new_AGEMA_signal_12213), .Z1_f (new_AGEMA_signal_12214) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M47), .A0_f (new_AGEMA_signal_10880), .A1_t (new_AGEMA_signal_10881), .A1_f (new_AGEMA_signal_10882), .B0_t (SubBytesIns_Inst_Sbox_13_M55), .B0_f (new_AGEMA_signal_11603), .B1_t (new_AGEMA_signal_11604), .B1_f (new_AGEMA_signal_11605), .Z0_t (SubBytesIns_Inst_Sbox_13_L3), .Z0_f (new_AGEMA_signal_12215), .Z1_t (new_AGEMA_signal_12216), .Z1_f (new_AGEMA_signal_12217) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M54), .A0_f (new_AGEMA_signal_11600), .A1_t (new_AGEMA_signal_11601), .A1_f (new_AGEMA_signal_11602), .B0_t (SubBytesIns_Inst_Sbox_13_M58), .B0_f (new_AGEMA_signal_11606), .B1_t (new_AGEMA_signal_11607), .B1_f (new_AGEMA_signal_11608), .Z0_t (SubBytesIns_Inst_Sbox_13_L4), .Z0_f (new_AGEMA_signal_12218), .Z1_t (new_AGEMA_signal_12219), .Z1_f (new_AGEMA_signal_12220) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M49), .A0_f (new_AGEMA_signal_11594), .A1_t (new_AGEMA_signal_11595), .A1_f (new_AGEMA_signal_11596), .B0_t (SubBytesIns_Inst_Sbox_13_M61), .B0_f (new_AGEMA_signal_11609), .B1_t (new_AGEMA_signal_11610), .B1_f (new_AGEMA_signal_11611), .Z0_t (SubBytesIns_Inst_Sbox_13_L5), .Z0_f (new_AGEMA_signal_12221), .Z1_t (new_AGEMA_signal_12222), .Z1_f (new_AGEMA_signal_12223) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M62), .A0_f (new_AGEMA_signal_12209), .A1_t (new_AGEMA_signal_12210), .A1_f (new_AGEMA_signal_12211), .B0_t (SubBytesIns_Inst_Sbox_13_L5), .B0_f (new_AGEMA_signal_12221), .B1_t (new_AGEMA_signal_12222), .B1_f (new_AGEMA_signal_12223), .Z0_t (SubBytesIns_Inst_Sbox_13_L6), .Z0_f (new_AGEMA_signal_12758), .Z1_t (new_AGEMA_signal_12759), .Z1_f (new_AGEMA_signal_12760) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M46), .A0_f (new_AGEMA_signal_11591), .A1_t (new_AGEMA_signal_11592), .A1_f (new_AGEMA_signal_11593), .B0_t (SubBytesIns_Inst_Sbox_13_L3), .B0_f (new_AGEMA_signal_12215), .B1_t (new_AGEMA_signal_12216), .B1_f (new_AGEMA_signal_12217), .Z0_t (SubBytesIns_Inst_Sbox_13_L7), .Z0_f (new_AGEMA_signal_12761), .Z1_t (new_AGEMA_signal_12762), .Z1_f (new_AGEMA_signal_12763) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M51), .A0_f (new_AGEMA_signal_10889), .A1_t (new_AGEMA_signal_10890), .A1_f (new_AGEMA_signal_10891), .B0_t (SubBytesIns_Inst_Sbox_13_M59), .B0_f (new_AGEMA_signal_10898), .B1_t (new_AGEMA_signal_10899), .B1_f (new_AGEMA_signal_10900), .Z0_t (SubBytesIns_Inst_Sbox_13_L8), .Z0_f (new_AGEMA_signal_11618), .Z1_t (new_AGEMA_signal_11619), .Z1_f (new_AGEMA_signal_11620) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M52), .A0_f (new_AGEMA_signal_11597), .A1_t (new_AGEMA_signal_11598), .A1_f (new_AGEMA_signal_11599), .B0_t (SubBytesIns_Inst_Sbox_13_M53), .B0_f (new_AGEMA_signal_12206), .B1_t (new_AGEMA_signal_12207), .B1_f (new_AGEMA_signal_12208), .Z0_t (SubBytesIns_Inst_Sbox_13_L9), .Z0_f (new_AGEMA_signal_12764), .Z1_t (new_AGEMA_signal_12765), .Z1_f (new_AGEMA_signal_12766) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M53), .A0_f (new_AGEMA_signal_12206), .A1_t (new_AGEMA_signal_12207), .A1_f (new_AGEMA_signal_12208), .B0_t (SubBytesIns_Inst_Sbox_13_L4), .B0_f (new_AGEMA_signal_12218), .B1_t (new_AGEMA_signal_12219), .B1_f (new_AGEMA_signal_12220), .Z0_t (SubBytesIns_Inst_Sbox_13_L10), .Z0_f (new_AGEMA_signal_12767), .Z1_t (new_AGEMA_signal_12768), .Z1_f (new_AGEMA_signal_12769) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M60), .A0_f (new_AGEMA_signal_10901), .A1_t (new_AGEMA_signal_10902), .A1_f (new_AGEMA_signal_10903), .B0_t (SubBytesIns_Inst_Sbox_13_L2), .B0_f (new_AGEMA_signal_12212), .B1_t (new_AGEMA_signal_12213), .B1_f (new_AGEMA_signal_12214), .Z0_t (SubBytesIns_Inst_Sbox_13_L11), .Z0_f (new_AGEMA_signal_12770), .Z1_t (new_AGEMA_signal_12771), .Z1_f (new_AGEMA_signal_12772) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M48), .A0_f (new_AGEMA_signal_10883), .A1_t (new_AGEMA_signal_10884), .A1_f (new_AGEMA_signal_10885), .B0_t (SubBytesIns_Inst_Sbox_13_M51), .B0_f (new_AGEMA_signal_10889), .B1_t (new_AGEMA_signal_10890), .B1_f (new_AGEMA_signal_10891), .Z0_t (SubBytesIns_Inst_Sbox_13_L12), .Z0_f (new_AGEMA_signal_11621), .Z1_t (new_AGEMA_signal_11622), .Z1_f (new_AGEMA_signal_11623) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M50), .A0_f (new_AGEMA_signal_10886), .A1_t (new_AGEMA_signal_10887), .A1_f (new_AGEMA_signal_10888), .B0_t (SubBytesIns_Inst_Sbox_13_L0), .B0_f (new_AGEMA_signal_12755), .B1_t (new_AGEMA_signal_12756), .B1_f (new_AGEMA_signal_12757), .Z0_t (SubBytesIns_Inst_Sbox_13_L13), .Z0_f (new_AGEMA_signal_13397), .Z1_t (new_AGEMA_signal_13398), .Z1_f (new_AGEMA_signal_13399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M52), .A0_f (new_AGEMA_signal_11597), .A1_t (new_AGEMA_signal_11598), .A1_f (new_AGEMA_signal_11599), .B0_t (SubBytesIns_Inst_Sbox_13_M61), .B0_f (new_AGEMA_signal_11609), .B1_t (new_AGEMA_signal_11610), .B1_f (new_AGEMA_signal_11611), .Z0_t (SubBytesIns_Inst_Sbox_13_L14), .Z0_f (new_AGEMA_signal_12224), .Z1_t (new_AGEMA_signal_12225), .Z1_f (new_AGEMA_signal_12226) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M55), .A0_f (new_AGEMA_signal_11603), .A1_t (new_AGEMA_signal_11604), .A1_f (new_AGEMA_signal_11605), .B0_t (SubBytesIns_Inst_Sbox_13_L1), .B0_f (new_AGEMA_signal_11615), .B1_t (new_AGEMA_signal_11616), .B1_f (new_AGEMA_signal_11617), .Z0_t (SubBytesIns_Inst_Sbox_13_L15), .Z0_f (new_AGEMA_signal_12227), .Z1_t (new_AGEMA_signal_12228), .Z1_f (new_AGEMA_signal_12229) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M56), .A0_f (new_AGEMA_signal_10892), .A1_t (new_AGEMA_signal_10893), .A1_f (new_AGEMA_signal_10894), .B0_t (SubBytesIns_Inst_Sbox_13_L0), .B0_f (new_AGEMA_signal_12755), .B1_t (new_AGEMA_signal_12756), .B1_f (new_AGEMA_signal_12757), .Z0_t (SubBytesIns_Inst_Sbox_13_L16), .Z0_f (new_AGEMA_signal_13400), .Z1_t (new_AGEMA_signal_13401), .Z1_f (new_AGEMA_signal_13402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M57), .A0_f (new_AGEMA_signal_10895), .A1_t (new_AGEMA_signal_10896), .A1_f (new_AGEMA_signal_10897), .B0_t (SubBytesIns_Inst_Sbox_13_L1), .B0_f (new_AGEMA_signal_11615), .B1_t (new_AGEMA_signal_11616), .B1_f (new_AGEMA_signal_11617), .Z0_t (SubBytesIns_Inst_Sbox_13_L17), .Z0_f (new_AGEMA_signal_12230), .Z1_t (new_AGEMA_signal_12231), .Z1_f (new_AGEMA_signal_12232) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M58), .A0_f (new_AGEMA_signal_11606), .A1_t (new_AGEMA_signal_11607), .A1_f (new_AGEMA_signal_11608), .B0_t (SubBytesIns_Inst_Sbox_13_L8), .B0_f (new_AGEMA_signal_11618), .B1_t (new_AGEMA_signal_11619), .B1_f (new_AGEMA_signal_11620), .Z0_t (SubBytesIns_Inst_Sbox_13_L18), .Z0_f (new_AGEMA_signal_12233), .Z1_t (new_AGEMA_signal_12234), .Z1_f (new_AGEMA_signal_12235) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M63), .A0_f (new_AGEMA_signal_11612), .A1_t (new_AGEMA_signal_11613), .A1_f (new_AGEMA_signal_11614), .B0_t (SubBytesIns_Inst_Sbox_13_L4), .B0_f (new_AGEMA_signal_12218), .B1_t (new_AGEMA_signal_12219), .B1_f (new_AGEMA_signal_12220), .Z0_t (SubBytesIns_Inst_Sbox_13_L19), .Z0_f (new_AGEMA_signal_12773), .Z1_t (new_AGEMA_signal_12774), .Z1_f (new_AGEMA_signal_12775) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L0), .A0_f (new_AGEMA_signal_12755), .A1_t (new_AGEMA_signal_12756), .A1_f (new_AGEMA_signal_12757), .B0_t (SubBytesIns_Inst_Sbox_13_L1), .B0_f (new_AGEMA_signal_11615), .B1_t (new_AGEMA_signal_11616), .B1_f (new_AGEMA_signal_11617), .Z0_t (SubBytesIns_Inst_Sbox_13_L20), .Z0_f (new_AGEMA_signal_13403), .Z1_t (new_AGEMA_signal_13404), .Z1_f (new_AGEMA_signal_13405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L1), .A0_f (new_AGEMA_signal_11615), .A1_t (new_AGEMA_signal_11616), .A1_f (new_AGEMA_signal_11617), .B0_t (SubBytesIns_Inst_Sbox_13_L7), .B0_f (new_AGEMA_signal_12761), .B1_t (new_AGEMA_signal_12762), .B1_f (new_AGEMA_signal_12763), .Z0_t (SubBytesIns_Inst_Sbox_13_L21), .Z0_f (new_AGEMA_signal_13406), .Z1_t (new_AGEMA_signal_13407), .Z1_f (new_AGEMA_signal_13408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L3), .A0_f (new_AGEMA_signal_12215), .A1_t (new_AGEMA_signal_12216), .A1_f (new_AGEMA_signal_12217), .B0_t (SubBytesIns_Inst_Sbox_13_L12), .B0_f (new_AGEMA_signal_11621), .B1_t (new_AGEMA_signal_11622), .B1_f (new_AGEMA_signal_11623), .Z0_t (SubBytesIns_Inst_Sbox_13_L22), .Z0_f (new_AGEMA_signal_12776), .Z1_t (new_AGEMA_signal_12777), .Z1_f (new_AGEMA_signal_12778) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L18), .A0_f (new_AGEMA_signal_12233), .A1_t (new_AGEMA_signal_12234), .A1_f (new_AGEMA_signal_12235), .B0_t (SubBytesIns_Inst_Sbox_13_L2), .B0_f (new_AGEMA_signal_12212), .B1_t (new_AGEMA_signal_12213), .B1_f (new_AGEMA_signal_12214), .Z0_t (SubBytesIns_Inst_Sbox_13_L23), .Z0_f (new_AGEMA_signal_12779), .Z1_t (new_AGEMA_signal_12780), .Z1_f (new_AGEMA_signal_12781) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L15), .A0_f (new_AGEMA_signal_12227), .A1_t (new_AGEMA_signal_12228), .A1_f (new_AGEMA_signal_12229), .B0_t (SubBytesIns_Inst_Sbox_13_L9), .B0_f (new_AGEMA_signal_12764), .B1_t (new_AGEMA_signal_12765), .B1_f (new_AGEMA_signal_12766), .Z0_t (SubBytesIns_Inst_Sbox_13_L24), .Z0_f (new_AGEMA_signal_13409), .Z1_t (new_AGEMA_signal_13410), .Z1_f (new_AGEMA_signal_13411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L6), .A0_f (new_AGEMA_signal_12758), .A1_t (new_AGEMA_signal_12759), .A1_f (new_AGEMA_signal_12760), .B0_t (SubBytesIns_Inst_Sbox_13_L10), .B0_f (new_AGEMA_signal_12767), .B1_t (new_AGEMA_signal_12768), .B1_f (new_AGEMA_signal_12769), .Z0_t (SubBytesIns_Inst_Sbox_13_L25), .Z0_f (new_AGEMA_signal_13412), .Z1_t (new_AGEMA_signal_13413), .Z1_f (new_AGEMA_signal_13414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L7), .A0_f (new_AGEMA_signal_12761), .A1_t (new_AGEMA_signal_12762), .A1_f (new_AGEMA_signal_12763), .B0_t (SubBytesIns_Inst_Sbox_13_L9), .B0_f (new_AGEMA_signal_12764), .B1_t (new_AGEMA_signal_12765), .B1_f (new_AGEMA_signal_12766), .Z0_t (SubBytesIns_Inst_Sbox_13_L26), .Z0_f (new_AGEMA_signal_13415), .Z1_t (new_AGEMA_signal_13416), .Z1_f (new_AGEMA_signal_13417) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L8), .A0_f (new_AGEMA_signal_11618), .A1_t (new_AGEMA_signal_11619), .A1_f (new_AGEMA_signal_11620), .B0_t (SubBytesIns_Inst_Sbox_13_L10), .B0_f (new_AGEMA_signal_12767), .B1_t (new_AGEMA_signal_12768), .B1_f (new_AGEMA_signal_12769), .Z0_t (SubBytesIns_Inst_Sbox_13_L27), .Z0_f (new_AGEMA_signal_13418), .Z1_t (new_AGEMA_signal_13419), .Z1_f (new_AGEMA_signal_13420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L11), .A0_f (new_AGEMA_signal_12770), .A1_t (new_AGEMA_signal_12771), .A1_f (new_AGEMA_signal_12772), .B0_t (SubBytesIns_Inst_Sbox_13_L14), .B0_f (new_AGEMA_signal_12224), .B1_t (new_AGEMA_signal_12225), .B1_f (new_AGEMA_signal_12226), .Z0_t (SubBytesIns_Inst_Sbox_13_L28), .Z0_f (new_AGEMA_signal_13421), .Z1_t (new_AGEMA_signal_13422), .Z1_f (new_AGEMA_signal_13423) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L11), .A0_f (new_AGEMA_signal_12770), .A1_t (new_AGEMA_signal_12771), .A1_f (new_AGEMA_signal_12772), .B0_t (SubBytesIns_Inst_Sbox_13_L17), .B0_f (new_AGEMA_signal_12230), .B1_t (new_AGEMA_signal_12231), .B1_f (new_AGEMA_signal_12232), .Z0_t (SubBytesIns_Inst_Sbox_13_L29), .Z0_f (new_AGEMA_signal_13424), .Z1_t (new_AGEMA_signal_13425), .Z1_f (new_AGEMA_signal_13426) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L6), .A0_f (new_AGEMA_signal_12758), .A1_t (new_AGEMA_signal_12759), .A1_f (new_AGEMA_signal_12760), .B0_t (SubBytesIns_Inst_Sbox_13_L24), .B0_f (new_AGEMA_signal_13409), .B1_t (new_AGEMA_signal_13410), .B1_f (new_AGEMA_signal_13411), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .Z0_f (new_AGEMA_signal_13913), .Z1_t (new_AGEMA_signal_13914), .Z1_f (new_AGEMA_signal_13915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L16), .A0_f (new_AGEMA_signal_13400), .A1_t (new_AGEMA_signal_13401), .A1_f (new_AGEMA_signal_13402), .B0_t (SubBytesIns_Inst_Sbox_13_L26), .B0_f (new_AGEMA_signal_13415), .B1_t (new_AGEMA_signal_13416), .B1_f (new_AGEMA_signal_13417), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .Z0_f (new_AGEMA_signal_13916), .Z1_t (new_AGEMA_signal_13917), .Z1_f (new_AGEMA_signal_13918) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L19), .A0_f (new_AGEMA_signal_12773), .A1_t (new_AGEMA_signal_12774), .A1_f (new_AGEMA_signal_12775), .B0_t (SubBytesIns_Inst_Sbox_13_L28), .B0_f (new_AGEMA_signal_13421), .B1_t (new_AGEMA_signal_13422), .B1_f (new_AGEMA_signal_13423), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .Z0_f (new_AGEMA_signal_13919), .Z1_t (new_AGEMA_signal_13920), .Z1_f (new_AGEMA_signal_13921) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L6), .A0_f (new_AGEMA_signal_12758), .A1_t (new_AGEMA_signal_12759), .A1_f (new_AGEMA_signal_12760), .B0_t (SubBytesIns_Inst_Sbox_13_L21), .B0_f (new_AGEMA_signal_13406), .B1_t (new_AGEMA_signal_13407), .B1_f (new_AGEMA_signal_13408), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .Z0_f (new_AGEMA_signal_13922), .Z1_t (new_AGEMA_signal_13923), .Z1_f (new_AGEMA_signal_13924) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L20), .A0_f (new_AGEMA_signal_13403), .A1_t (new_AGEMA_signal_13404), .A1_f (new_AGEMA_signal_13405), .B0_t (SubBytesIns_Inst_Sbox_13_L22), .B0_f (new_AGEMA_signal_12776), .B1_t (new_AGEMA_signal_12777), .B1_f (new_AGEMA_signal_12778), .Z0_t (MixColumnsInput[43]), .Z0_f (new_AGEMA_signal_13925), .Z1_t (new_AGEMA_signal_13926), .Z1_f (new_AGEMA_signal_13927) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L25), .A0_f (new_AGEMA_signal_13412), .A1_t (new_AGEMA_signal_13413), .A1_f (new_AGEMA_signal_13414), .B0_t (SubBytesIns_Inst_Sbox_13_L29), .B0_f (new_AGEMA_signal_13424), .B1_t (new_AGEMA_signal_13425), .B1_f (new_AGEMA_signal_13426), .Z0_t (MixColumnsInput[42]), .Z0_f (new_AGEMA_signal_13928), .Z1_t (new_AGEMA_signal_13929), .Z1_f (new_AGEMA_signal_13930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L13), .A0_f (new_AGEMA_signal_13397), .A1_t (new_AGEMA_signal_13398), .A1_f (new_AGEMA_signal_13399), .B0_t (SubBytesIns_Inst_Sbox_13_L27), .B0_f (new_AGEMA_signal_13418), .B1_t (new_AGEMA_signal_13419), .B1_f (new_AGEMA_signal_13420), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .Z0_f (new_AGEMA_signal_13931), .Z1_t (new_AGEMA_signal_13932), .Z1_f (new_AGEMA_signal_13933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L6), .A0_f (new_AGEMA_signal_12758), .A1_t (new_AGEMA_signal_12759), .A1_f (new_AGEMA_signal_12760), .B0_t (SubBytesIns_Inst_Sbox_13_L23), .B0_f (new_AGEMA_signal_12779), .B1_t (new_AGEMA_signal_12780), .B1_f (new_AGEMA_signal_12781), .Z0_t (MixColumnsInput[40]), .Z0_f (new_AGEMA_signal_13427), .Z1_t (new_AGEMA_signal_13428), .Z1_f (new_AGEMA_signal_13429) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (ciphertext_s0_t[116]), .B0_f (ciphertext_s0_f[116]), .B1_t (ciphertext_s1_t[116]), .B1_f (ciphertext_s1_f[116]), .Z0_t (SubBytesIns_Inst_Sbox_14_T1), .Z0_f (new_AGEMA_signal_6766), .Z1_t (new_AGEMA_signal_6767), .Z1_f (new_AGEMA_signal_6768) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (ciphertext_s0_t[114]), .B0_f (ciphertext_s0_f[114]), .B1_t (ciphertext_s1_t[114]), .B1_f (ciphertext_s1_f[114]), .Z0_t (SubBytesIns_Inst_Sbox_14_T2), .Z0_f (new_AGEMA_signal_6769), .Z1_t (new_AGEMA_signal_6770), .Z1_f (new_AGEMA_signal_6771) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (ciphertext_s0_t[113]), .B0_f (ciphertext_s0_f[113]), .B1_t (ciphertext_s1_t[113]), .B1_f (ciphertext_s1_f[113]), .Z0_t (SubBytesIns_Inst_Sbox_14_T3), .Z0_f (new_AGEMA_signal_6772), .Z1_t (new_AGEMA_signal_6773), .Z1_f (new_AGEMA_signal_6774) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[116]), .A0_f (ciphertext_s0_f[116]), .A1_t (ciphertext_s1_t[116]), .A1_f (ciphertext_s1_f[116]), .B0_t (ciphertext_s0_t[114]), .B0_f (ciphertext_s0_f[114]), .B1_t (ciphertext_s1_t[114]), .B1_f (ciphertext_s1_f[114]), .Z0_t (SubBytesIns_Inst_Sbox_14_T4), .Z0_f (new_AGEMA_signal_6775), .Z1_t (new_AGEMA_signal_6776), .Z1_f (new_AGEMA_signal_6777) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[115]), .A0_f (ciphertext_s0_f[115]), .A1_t (ciphertext_s1_t[115]), .A1_f (ciphertext_s1_f[115]), .B0_t (ciphertext_s0_t[113]), .B0_f (ciphertext_s0_f[113]), .B1_t (ciphertext_s1_t[113]), .B1_f (ciphertext_s1_f[113]), .Z0_t (SubBytesIns_Inst_Sbox_14_T5), .Z0_f (new_AGEMA_signal_6778), .Z1_t (new_AGEMA_signal_6779), .Z1_f (new_AGEMA_signal_6780) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T1), .A0_f (new_AGEMA_signal_6766), .A1_t (new_AGEMA_signal_6767), .A1_f (new_AGEMA_signal_6768), .B0_t (SubBytesIns_Inst_Sbox_14_T5), .B0_f (new_AGEMA_signal_6778), .B1_t (new_AGEMA_signal_6779), .B1_f (new_AGEMA_signal_6780), .Z0_t (SubBytesIns_Inst_Sbox_14_T6), .Z0_f (new_AGEMA_signal_7264), .Z1_t (new_AGEMA_signal_7265), .Z1_f (new_AGEMA_signal_7266) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[118]), .A0_f (ciphertext_s0_f[118]), .A1_t (ciphertext_s1_t[118]), .A1_f (ciphertext_s1_f[118]), .B0_t (ciphertext_s0_t[117]), .B0_f (ciphertext_s0_f[117]), .B1_t (ciphertext_s1_t[117]), .B1_f (ciphertext_s1_f[117]), .Z0_t (SubBytesIns_Inst_Sbox_14_T7), .Z0_f (new_AGEMA_signal_6781), .Z1_t (new_AGEMA_signal_6782), .Z1_f (new_AGEMA_signal_6783) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[112]), .A0_f (ciphertext_s0_f[112]), .A1_t (ciphertext_s1_t[112]), .A1_f (ciphertext_s1_f[112]), .B0_t (SubBytesIns_Inst_Sbox_14_T6), .B0_f (new_AGEMA_signal_7264), .B1_t (new_AGEMA_signal_7265), .B1_f (new_AGEMA_signal_7266), .Z0_t (SubBytesIns_Inst_Sbox_14_T8), .Z0_f (new_AGEMA_signal_8018), .Z1_t (new_AGEMA_signal_8019), .Z1_f (new_AGEMA_signal_8020) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[112]), .A0_f (ciphertext_s0_f[112]), .A1_t (ciphertext_s1_t[112]), .A1_f (ciphertext_s1_f[112]), .B0_t (SubBytesIns_Inst_Sbox_14_T7), .B0_f (new_AGEMA_signal_6781), .B1_t (new_AGEMA_signal_6782), .B1_f (new_AGEMA_signal_6783), .Z0_t (SubBytesIns_Inst_Sbox_14_T9), .Z0_f (new_AGEMA_signal_7267), .Z1_t (new_AGEMA_signal_7268), .Z1_f (new_AGEMA_signal_7269) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T6), .A0_f (new_AGEMA_signal_7264), .A1_t (new_AGEMA_signal_7265), .A1_f (new_AGEMA_signal_7266), .B0_t (SubBytesIns_Inst_Sbox_14_T7), .B0_f (new_AGEMA_signal_6781), .B1_t (new_AGEMA_signal_6782), .B1_f (new_AGEMA_signal_6783), .Z0_t (SubBytesIns_Inst_Sbox_14_T10), .Z0_f (new_AGEMA_signal_8021), .Z1_t (new_AGEMA_signal_8022), .Z1_f (new_AGEMA_signal_8023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[118]), .A0_f (ciphertext_s0_f[118]), .A1_t (ciphertext_s1_t[118]), .A1_f (ciphertext_s1_f[118]), .B0_t (ciphertext_s0_t[114]), .B0_f (ciphertext_s0_f[114]), .B1_t (ciphertext_s1_t[114]), .B1_f (ciphertext_s1_f[114]), .Z0_t (SubBytesIns_Inst_Sbox_14_T11), .Z0_f (new_AGEMA_signal_6784), .Z1_t (new_AGEMA_signal_6785), .Z1_f (new_AGEMA_signal_6786) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[117]), .A0_f (ciphertext_s0_f[117]), .A1_t (ciphertext_s1_t[117]), .A1_f (ciphertext_s1_f[117]), .B0_t (ciphertext_s0_t[114]), .B0_f (ciphertext_s0_f[114]), .B1_t (ciphertext_s1_t[114]), .B1_f (ciphertext_s1_f[114]), .Z0_t (SubBytesIns_Inst_Sbox_14_T12), .Z0_f (new_AGEMA_signal_6787), .Z1_t (new_AGEMA_signal_6788), .Z1_f (new_AGEMA_signal_6789) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T3), .A0_f (new_AGEMA_signal_6772), .A1_t (new_AGEMA_signal_6773), .A1_f (new_AGEMA_signal_6774), .B0_t (SubBytesIns_Inst_Sbox_14_T4), .B0_f (new_AGEMA_signal_6775), .B1_t (new_AGEMA_signal_6776), .B1_f (new_AGEMA_signal_6777), .Z0_t (SubBytesIns_Inst_Sbox_14_T13), .Z0_f (new_AGEMA_signal_7270), .Z1_t (new_AGEMA_signal_7271), .Z1_f (new_AGEMA_signal_7272) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T6), .A0_f (new_AGEMA_signal_7264), .A1_t (new_AGEMA_signal_7265), .A1_f (new_AGEMA_signal_7266), .B0_t (SubBytesIns_Inst_Sbox_14_T11), .B0_f (new_AGEMA_signal_6784), .B1_t (new_AGEMA_signal_6785), .B1_f (new_AGEMA_signal_6786), .Z0_t (SubBytesIns_Inst_Sbox_14_T14), .Z0_f (new_AGEMA_signal_8024), .Z1_t (new_AGEMA_signal_8025), .Z1_f (new_AGEMA_signal_8026) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T5), .A0_f (new_AGEMA_signal_6778), .A1_t (new_AGEMA_signal_6779), .A1_f (new_AGEMA_signal_6780), .B0_t (SubBytesIns_Inst_Sbox_14_T11), .B0_f (new_AGEMA_signal_6784), .B1_t (new_AGEMA_signal_6785), .B1_f (new_AGEMA_signal_6786), .Z0_t (SubBytesIns_Inst_Sbox_14_T15), .Z0_f (new_AGEMA_signal_7273), .Z1_t (new_AGEMA_signal_7274), .Z1_f (new_AGEMA_signal_7275) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T5), .A0_f (new_AGEMA_signal_6778), .A1_t (new_AGEMA_signal_6779), .A1_f (new_AGEMA_signal_6780), .B0_t (SubBytesIns_Inst_Sbox_14_T12), .B0_f (new_AGEMA_signal_6787), .B1_t (new_AGEMA_signal_6788), .B1_f (new_AGEMA_signal_6789), .Z0_t (SubBytesIns_Inst_Sbox_14_T16), .Z0_f (new_AGEMA_signal_7276), .Z1_t (new_AGEMA_signal_7277), .Z1_f (new_AGEMA_signal_7278) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T9), .A0_f (new_AGEMA_signal_7267), .A1_t (new_AGEMA_signal_7268), .A1_f (new_AGEMA_signal_7269), .B0_t (SubBytesIns_Inst_Sbox_14_T16), .B0_f (new_AGEMA_signal_7276), .B1_t (new_AGEMA_signal_7277), .B1_f (new_AGEMA_signal_7278), .Z0_t (SubBytesIns_Inst_Sbox_14_T17), .Z0_f (new_AGEMA_signal_8027), .Z1_t (new_AGEMA_signal_8028), .Z1_f (new_AGEMA_signal_8029) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[116]), .A0_f (ciphertext_s0_f[116]), .A1_t (ciphertext_s1_t[116]), .A1_f (ciphertext_s1_f[116]), .B0_t (ciphertext_s0_t[112]), .B0_f (ciphertext_s0_f[112]), .B1_t (ciphertext_s1_t[112]), .B1_f (ciphertext_s1_f[112]), .Z0_t (SubBytesIns_Inst_Sbox_14_T18), .Z0_f (new_AGEMA_signal_6790), .Z1_t (new_AGEMA_signal_6791), .Z1_f (new_AGEMA_signal_6792) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T7), .A0_f (new_AGEMA_signal_6781), .A1_t (new_AGEMA_signal_6782), .A1_f (new_AGEMA_signal_6783), .B0_t (SubBytesIns_Inst_Sbox_14_T18), .B0_f (new_AGEMA_signal_6790), .B1_t (new_AGEMA_signal_6791), .B1_f (new_AGEMA_signal_6792), .Z0_t (SubBytesIns_Inst_Sbox_14_T19), .Z0_f (new_AGEMA_signal_7279), .Z1_t (new_AGEMA_signal_7280), .Z1_f (new_AGEMA_signal_7281) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T1), .A0_f (new_AGEMA_signal_6766), .A1_t (new_AGEMA_signal_6767), .A1_f (new_AGEMA_signal_6768), .B0_t (SubBytesIns_Inst_Sbox_14_T19), .B0_f (new_AGEMA_signal_7279), .B1_t (new_AGEMA_signal_7280), .B1_f (new_AGEMA_signal_7281), .Z0_t (SubBytesIns_Inst_Sbox_14_T20), .Z0_f (new_AGEMA_signal_8030), .Z1_t (new_AGEMA_signal_8031), .Z1_f (new_AGEMA_signal_8032) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[113]), .A0_f (ciphertext_s0_f[113]), .A1_t (ciphertext_s1_t[113]), .A1_f (ciphertext_s1_f[113]), .B0_t (ciphertext_s0_t[112]), .B0_f (ciphertext_s0_f[112]), .B1_t (ciphertext_s1_t[112]), .B1_f (ciphertext_s1_f[112]), .Z0_t (SubBytesIns_Inst_Sbox_14_T21), .Z0_f (new_AGEMA_signal_6793), .Z1_t (new_AGEMA_signal_6794), .Z1_f (new_AGEMA_signal_6795) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T7), .A0_f (new_AGEMA_signal_6781), .A1_t (new_AGEMA_signal_6782), .A1_f (new_AGEMA_signal_6783), .B0_t (SubBytesIns_Inst_Sbox_14_T21), .B0_f (new_AGEMA_signal_6793), .B1_t (new_AGEMA_signal_6794), .B1_f (new_AGEMA_signal_6795), .Z0_t (SubBytesIns_Inst_Sbox_14_T22), .Z0_f (new_AGEMA_signal_7282), .Z1_t (new_AGEMA_signal_7283), .Z1_f (new_AGEMA_signal_7284) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T2), .A0_f (new_AGEMA_signal_6769), .A1_t (new_AGEMA_signal_6770), .A1_f (new_AGEMA_signal_6771), .B0_t (SubBytesIns_Inst_Sbox_14_T22), .B0_f (new_AGEMA_signal_7282), .B1_t (new_AGEMA_signal_7283), .B1_f (new_AGEMA_signal_7284), .Z0_t (SubBytesIns_Inst_Sbox_14_T23), .Z0_f (new_AGEMA_signal_8033), .Z1_t (new_AGEMA_signal_8034), .Z1_f (new_AGEMA_signal_8035) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T2), .A0_f (new_AGEMA_signal_6769), .A1_t (new_AGEMA_signal_6770), .A1_f (new_AGEMA_signal_6771), .B0_t (SubBytesIns_Inst_Sbox_14_T10), .B0_f (new_AGEMA_signal_8021), .B1_t (new_AGEMA_signal_8022), .B1_f (new_AGEMA_signal_8023), .Z0_t (SubBytesIns_Inst_Sbox_14_T24), .Z0_f (new_AGEMA_signal_8582), .Z1_t (new_AGEMA_signal_8583), .Z1_f (new_AGEMA_signal_8584) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T20), .A0_f (new_AGEMA_signal_8030), .A1_t (new_AGEMA_signal_8031), .A1_f (new_AGEMA_signal_8032), .B0_t (SubBytesIns_Inst_Sbox_14_T17), .B0_f (new_AGEMA_signal_8027), .B1_t (new_AGEMA_signal_8028), .B1_f (new_AGEMA_signal_8029), .Z0_t (SubBytesIns_Inst_Sbox_14_T25), .Z0_f (new_AGEMA_signal_8585), .Z1_t (new_AGEMA_signal_8586), .Z1_f (new_AGEMA_signal_8587) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T3), .A0_f (new_AGEMA_signal_6772), .A1_t (new_AGEMA_signal_6773), .A1_f (new_AGEMA_signal_6774), .B0_t (SubBytesIns_Inst_Sbox_14_T16), .B0_f (new_AGEMA_signal_7276), .B1_t (new_AGEMA_signal_7277), .B1_f (new_AGEMA_signal_7278), .Z0_t (SubBytesIns_Inst_Sbox_14_T26), .Z0_f (new_AGEMA_signal_8036), .Z1_t (new_AGEMA_signal_8037), .Z1_f (new_AGEMA_signal_8038) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T1), .A0_f (new_AGEMA_signal_6766), .A1_t (new_AGEMA_signal_6767), .A1_f (new_AGEMA_signal_6768), .B0_t (SubBytesIns_Inst_Sbox_14_T12), .B0_f (new_AGEMA_signal_6787), .B1_t (new_AGEMA_signal_6788), .B1_f (new_AGEMA_signal_6789), .Z0_t (SubBytesIns_Inst_Sbox_14_T27), .Z0_f (new_AGEMA_signal_7285), .Z1_t (new_AGEMA_signal_7286), .Z1_f (new_AGEMA_signal_7287) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T13), .A0_f (new_AGEMA_signal_7270), .A1_t (new_AGEMA_signal_7271), .A1_f (new_AGEMA_signal_7272), .B0_t (SubBytesIns_Inst_Sbox_14_T6), .B0_f (new_AGEMA_signal_7264), .B1_t (new_AGEMA_signal_7265), .B1_f (new_AGEMA_signal_7266), .Z0_t (SubBytesIns_Inst_Sbox_14_M1), .Z0_f (new_AGEMA_signal_8039), .Z1_t (new_AGEMA_signal_8040), .Z1_f (new_AGEMA_signal_8041) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T23), .A0_f (new_AGEMA_signal_8033), .A1_t (new_AGEMA_signal_8034), .A1_f (new_AGEMA_signal_8035), .B0_t (SubBytesIns_Inst_Sbox_14_T8), .B0_f (new_AGEMA_signal_8018), .B1_t (new_AGEMA_signal_8019), .B1_f (new_AGEMA_signal_8020), .Z0_t (SubBytesIns_Inst_Sbox_14_M2), .Z0_f (new_AGEMA_signal_8588), .Z1_t (new_AGEMA_signal_8589), .Z1_f (new_AGEMA_signal_8590) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T14), .A0_f (new_AGEMA_signal_8024), .A1_t (new_AGEMA_signal_8025), .A1_f (new_AGEMA_signal_8026), .B0_t (SubBytesIns_Inst_Sbox_14_M1), .B0_f (new_AGEMA_signal_8039), .B1_t (new_AGEMA_signal_8040), .B1_f (new_AGEMA_signal_8041), .Z0_t (SubBytesIns_Inst_Sbox_14_M3), .Z0_f (new_AGEMA_signal_8591), .Z1_t (new_AGEMA_signal_8592), .Z1_f (new_AGEMA_signal_8593) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T19), .A0_f (new_AGEMA_signal_7279), .A1_t (new_AGEMA_signal_7280), .A1_f (new_AGEMA_signal_7281), .B0_t (ciphertext_s0_t[112]), .B0_f (ciphertext_s0_f[112]), .B1_t (ciphertext_s1_t[112]), .B1_f (ciphertext_s1_f[112]), .Z0_t (SubBytesIns_Inst_Sbox_14_M4), .Z0_f (new_AGEMA_signal_8042), .Z1_t (new_AGEMA_signal_8043), .Z1_f (new_AGEMA_signal_8044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M4), .A0_f (new_AGEMA_signal_8042), .A1_t (new_AGEMA_signal_8043), .A1_f (new_AGEMA_signal_8044), .B0_t (SubBytesIns_Inst_Sbox_14_M1), .B0_f (new_AGEMA_signal_8039), .B1_t (new_AGEMA_signal_8040), .B1_f (new_AGEMA_signal_8041), .Z0_t (SubBytesIns_Inst_Sbox_14_M5), .Z0_f (new_AGEMA_signal_8594), .Z1_t (new_AGEMA_signal_8595), .Z1_f (new_AGEMA_signal_8596) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T3), .A0_f (new_AGEMA_signal_6772), .A1_t (new_AGEMA_signal_6773), .A1_f (new_AGEMA_signal_6774), .B0_t (SubBytesIns_Inst_Sbox_14_T16), .B0_f (new_AGEMA_signal_7276), .B1_t (new_AGEMA_signal_7277), .B1_f (new_AGEMA_signal_7278), .Z0_t (SubBytesIns_Inst_Sbox_14_M6), .Z0_f (new_AGEMA_signal_8045), .Z1_t (new_AGEMA_signal_8046), .Z1_f (new_AGEMA_signal_8047) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T22), .A0_f (new_AGEMA_signal_7282), .A1_t (new_AGEMA_signal_7283), .A1_f (new_AGEMA_signal_7284), .B0_t (SubBytesIns_Inst_Sbox_14_T9), .B0_f (new_AGEMA_signal_7267), .B1_t (new_AGEMA_signal_7268), .B1_f (new_AGEMA_signal_7269), .Z0_t (SubBytesIns_Inst_Sbox_14_M7), .Z0_f (new_AGEMA_signal_8048), .Z1_t (new_AGEMA_signal_8049), .Z1_f (new_AGEMA_signal_8050) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T26), .A0_f (new_AGEMA_signal_8036), .A1_t (new_AGEMA_signal_8037), .A1_f (new_AGEMA_signal_8038), .B0_t (SubBytesIns_Inst_Sbox_14_M6), .B0_f (new_AGEMA_signal_8045), .B1_t (new_AGEMA_signal_8046), .B1_f (new_AGEMA_signal_8047), .Z0_t (SubBytesIns_Inst_Sbox_14_M8), .Z0_f (new_AGEMA_signal_8597), .Z1_t (new_AGEMA_signal_8598), .Z1_f (new_AGEMA_signal_8599) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T20), .A0_f (new_AGEMA_signal_8030), .A1_t (new_AGEMA_signal_8031), .A1_f (new_AGEMA_signal_8032), .B0_t (SubBytesIns_Inst_Sbox_14_T17), .B0_f (new_AGEMA_signal_8027), .B1_t (new_AGEMA_signal_8028), .B1_f (new_AGEMA_signal_8029), .Z0_t (SubBytesIns_Inst_Sbox_14_M9), .Z0_f (new_AGEMA_signal_8600), .Z1_t (new_AGEMA_signal_8601), .Z1_f (new_AGEMA_signal_8602) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M9), .A0_f (new_AGEMA_signal_8600), .A1_t (new_AGEMA_signal_8601), .A1_f (new_AGEMA_signal_8602), .B0_t (SubBytesIns_Inst_Sbox_14_M6), .B0_f (new_AGEMA_signal_8045), .B1_t (new_AGEMA_signal_8046), .B1_f (new_AGEMA_signal_8047), .Z0_t (SubBytesIns_Inst_Sbox_14_M10), .Z0_f (new_AGEMA_signal_8906), .Z1_t (new_AGEMA_signal_8907), .Z1_f (new_AGEMA_signal_8908) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T1), .A0_f (new_AGEMA_signal_6766), .A1_t (new_AGEMA_signal_6767), .A1_f (new_AGEMA_signal_6768), .B0_t (SubBytesIns_Inst_Sbox_14_T15), .B0_f (new_AGEMA_signal_7273), .B1_t (new_AGEMA_signal_7274), .B1_f (new_AGEMA_signal_7275), .Z0_t (SubBytesIns_Inst_Sbox_14_M11), .Z0_f (new_AGEMA_signal_8051), .Z1_t (new_AGEMA_signal_8052), .Z1_f (new_AGEMA_signal_8053) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T4), .A0_f (new_AGEMA_signal_6775), .A1_t (new_AGEMA_signal_6776), .A1_f (new_AGEMA_signal_6777), .B0_t (SubBytesIns_Inst_Sbox_14_T27), .B0_f (new_AGEMA_signal_7285), .B1_t (new_AGEMA_signal_7286), .B1_f (new_AGEMA_signal_7287), .Z0_t (SubBytesIns_Inst_Sbox_14_M12), .Z0_f (new_AGEMA_signal_8054), .Z1_t (new_AGEMA_signal_8055), .Z1_f (new_AGEMA_signal_8056) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M12), .A0_f (new_AGEMA_signal_8054), .A1_t (new_AGEMA_signal_8055), .A1_f (new_AGEMA_signal_8056), .B0_t (SubBytesIns_Inst_Sbox_14_M11), .B0_f (new_AGEMA_signal_8051), .B1_t (new_AGEMA_signal_8052), .B1_f (new_AGEMA_signal_8053), .Z0_t (SubBytesIns_Inst_Sbox_14_M13), .Z0_f (new_AGEMA_signal_8603), .Z1_t (new_AGEMA_signal_8604), .Z1_f (new_AGEMA_signal_8605) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T2), .A0_f (new_AGEMA_signal_6769), .A1_t (new_AGEMA_signal_6770), .A1_f (new_AGEMA_signal_6771), .B0_t (SubBytesIns_Inst_Sbox_14_T10), .B0_f (new_AGEMA_signal_8021), .B1_t (new_AGEMA_signal_8022), .B1_f (new_AGEMA_signal_8023), .Z0_t (SubBytesIns_Inst_Sbox_14_M14), .Z0_f (new_AGEMA_signal_8606), .Z1_t (new_AGEMA_signal_8607), .Z1_f (new_AGEMA_signal_8608) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M14), .A0_f (new_AGEMA_signal_8606), .A1_t (new_AGEMA_signal_8607), .A1_f (new_AGEMA_signal_8608), .B0_t (SubBytesIns_Inst_Sbox_14_M11), .B0_f (new_AGEMA_signal_8051), .B1_t (new_AGEMA_signal_8052), .B1_f (new_AGEMA_signal_8053), .Z0_t (SubBytesIns_Inst_Sbox_14_M15), .Z0_f (new_AGEMA_signal_8909), .Z1_t (new_AGEMA_signal_8910), .Z1_f (new_AGEMA_signal_8911) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M3), .A0_f (new_AGEMA_signal_8591), .A1_t (new_AGEMA_signal_8592), .A1_f (new_AGEMA_signal_8593), .B0_t (SubBytesIns_Inst_Sbox_14_M2), .B0_f (new_AGEMA_signal_8588), .B1_t (new_AGEMA_signal_8589), .B1_f (new_AGEMA_signal_8590), .Z0_t (SubBytesIns_Inst_Sbox_14_M16), .Z0_f (new_AGEMA_signal_8912), .Z1_t (new_AGEMA_signal_8913), .Z1_f (new_AGEMA_signal_8914) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M5), .A0_f (new_AGEMA_signal_8594), .A1_t (new_AGEMA_signal_8595), .A1_f (new_AGEMA_signal_8596), .B0_t (SubBytesIns_Inst_Sbox_14_T24), .B0_f (new_AGEMA_signal_8582), .B1_t (new_AGEMA_signal_8583), .B1_f (new_AGEMA_signal_8584), .Z0_t (SubBytesIns_Inst_Sbox_14_M17), .Z0_f (new_AGEMA_signal_8915), .Z1_t (new_AGEMA_signal_8916), .Z1_f (new_AGEMA_signal_8917) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M8), .A0_f (new_AGEMA_signal_8597), .A1_t (new_AGEMA_signal_8598), .A1_f (new_AGEMA_signal_8599), .B0_t (SubBytesIns_Inst_Sbox_14_M7), .B0_f (new_AGEMA_signal_8048), .B1_t (new_AGEMA_signal_8049), .B1_f (new_AGEMA_signal_8050), .Z0_t (SubBytesIns_Inst_Sbox_14_M18), .Z0_f (new_AGEMA_signal_8918), .Z1_t (new_AGEMA_signal_8919), .Z1_f (new_AGEMA_signal_8920) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M10), .A0_f (new_AGEMA_signal_8906), .A1_t (new_AGEMA_signal_8907), .A1_f (new_AGEMA_signal_8908), .B0_t (SubBytesIns_Inst_Sbox_14_M15), .B0_f (new_AGEMA_signal_8909), .B1_t (new_AGEMA_signal_8910), .B1_f (new_AGEMA_signal_8911), .Z0_t (SubBytesIns_Inst_Sbox_14_M19), .Z0_f (new_AGEMA_signal_9152), .Z1_t (new_AGEMA_signal_9153), .Z1_f (new_AGEMA_signal_9154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M16), .A0_f (new_AGEMA_signal_8912), .A1_t (new_AGEMA_signal_8913), .A1_f (new_AGEMA_signal_8914), .B0_t (SubBytesIns_Inst_Sbox_14_M13), .B0_f (new_AGEMA_signal_8603), .B1_t (new_AGEMA_signal_8604), .B1_f (new_AGEMA_signal_8605), .Z0_t (SubBytesIns_Inst_Sbox_14_M20), .Z0_f (new_AGEMA_signal_9155), .Z1_t (new_AGEMA_signal_9156), .Z1_f (new_AGEMA_signal_9157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M17), .A0_f (new_AGEMA_signal_8915), .A1_t (new_AGEMA_signal_8916), .A1_f (new_AGEMA_signal_8917), .B0_t (SubBytesIns_Inst_Sbox_14_M15), .B0_f (new_AGEMA_signal_8909), .B1_t (new_AGEMA_signal_8910), .B1_f (new_AGEMA_signal_8911), .Z0_t (SubBytesIns_Inst_Sbox_14_M21), .Z0_f (new_AGEMA_signal_9158), .Z1_t (new_AGEMA_signal_9159), .Z1_f (new_AGEMA_signal_9160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M18), .A0_f (new_AGEMA_signal_8918), .A1_t (new_AGEMA_signal_8919), .A1_f (new_AGEMA_signal_8920), .B0_t (SubBytesIns_Inst_Sbox_14_M13), .B0_f (new_AGEMA_signal_8603), .B1_t (new_AGEMA_signal_8604), .B1_f (new_AGEMA_signal_8605), .Z0_t (SubBytesIns_Inst_Sbox_14_M22), .Z0_f (new_AGEMA_signal_9161), .Z1_t (new_AGEMA_signal_9162), .Z1_f (new_AGEMA_signal_9163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M19), .A0_f (new_AGEMA_signal_9152), .A1_t (new_AGEMA_signal_9153), .A1_f (new_AGEMA_signal_9154), .B0_t (SubBytesIns_Inst_Sbox_14_T25), .B0_f (new_AGEMA_signal_8585), .B1_t (new_AGEMA_signal_8586), .B1_f (new_AGEMA_signal_8587), .Z0_t (SubBytesIns_Inst_Sbox_14_M23), .Z0_f (new_AGEMA_signal_9392), .Z1_t (new_AGEMA_signal_9393), .Z1_f (new_AGEMA_signal_9394) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M22), .A0_f (new_AGEMA_signal_9161), .A1_t (new_AGEMA_signal_9162), .A1_f (new_AGEMA_signal_9163), .B0_t (SubBytesIns_Inst_Sbox_14_M23), .B0_f (new_AGEMA_signal_9392), .B1_t (new_AGEMA_signal_9393), .B1_f (new_AGEMA_signal_9394), .Z0_t (SubBytesIns_Inst_Sbox_14_M24), .Z0_f (new_AGEMA_signal_9686), .Z1_t (new_AGEMA_signal_9687), .Z1_f (new_AGEMA_signal_9688) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M22), .A0_f (new_AGEMA_signal_9161), .A1_t (new_AGEMA_signal_9162), .A1_f (new_AGEMA_signal_9163), .B0_t (SubBytesIns_Inst_Sbox_14_M20), .B0_f (new_AGEMA_signal_9155), .B1_t (new_AGEMA_signal_9156), .B1_f (new_AGEMA_signal_9157), .Z0_t (SubBytesIns_Inst_Sbox_14_M25), .Z0_f (new_AGEMA_signal_9395), .Z1_t (new_AGEMA_signal_9396), .Z1_f (new_AGEMA_signal_9397) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M21), .A0_f (new_AGEMA_signal_9158), .A1_t (new_AGEMA_signal_9159), .A1_f (new_AGEMA_signal_9160), .B0_t (SubBytesIns_Inst_Sbox_14_M25), .B0_f (new_AGEMA_signal_9395), .B1_t (new_AGEMA_signal_9396), .B1_f (new_AGEMA_signal_9397), .Z0_t (SubBytesIns_Inst_Sbox_14_M26), .Z0_f (new_AGEMA_signal_9689), .Z1_t (new_AGEMA_signal_9690), .Z1_f (new_AGEMA_signal_9691) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M20), .A0_f (new_AGEMA_signal_9155), .A1_t (new_AGEMA_signal_9156), .A1_f (new_AGEMA_signal_9157), .B0_t (SubBytesIns_Inst_Sbox_14_M21), .B0_f (new_AGEMA_signal_9158), .B1_t (new_AGEMA_signal_9159), .B1_f (new_AGEMA_signal_9160), .Z0_t (SubBytesIns_Inst_Sbox_14_M27), .Z0_f (new_AGEMA_signal_9398), .Z1_t (new_AGEMA_signal_9399), .Z1_f (new_AGEMA_signal_9400) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M23), .A0_f (new_AGEMA_signal_9392), .A1_t (new_AGEMA_signal_9393), .A1_f (new_AGEMA_signal_9394), .B0_t (SubBytesIns_Inst_Sbox_14_M25), .B0_f (new_AGEMA_signal_9395), .B1_t (new_AGEMA_signal_9396), .B1_f (new_AGEMA_signal_9397), .Z0_t (SubBytesIns_Inst_Sbox_14_M28), .Z0_f (new_AGEMA_signal_9692), .Z1_t (new_AGEMA_signal_9693), .Z1_f (new_AGEMA_signal_9694) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M28), .A0_f (new_AGEMA_signal_9692), .A1_t (new_AGEMA_signal_9693), .A1_f (new_AGEMA_signal_9694), .B0_t (SubBytesIns_Inst_Sbox_14_M27), .B0_f (new_AGEMA_signal_9398), .B1_t (new_AGEMA_signal_9399), .B1_f (new_AGEMA_signal_9400), .Z0_t (SubBytesIns_Inst_Sbox_14_M29), .Z0_f (new_AGEMA_signal_9986), .Z1_t (new_AGEMA_signal_9987), .Z1_f (new_AGEMA_signal_9988) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M26), .A0_f (new_AGEMA_signal_9689), .A1_t (new_AGEMA_signal_9690), .A1_f (new_AGEMA_signal_9691), .B0_t (SubBytesIns_Inst_Sbox_14_M24), .B0_f (new_AGEMA_signal_9686), .B1_t (new_AGEMA_signal_9687), .B1_f (new_AGEMA_signal_9688), .Z0_t (SubBytesIns_Inst_Sbox_14_M30), .Z0_f (new_AGEMA_signal_9989), .Z1_t (new_AGEMA_signal_9990), .Z1_f (new_AGEMA_signal_9991) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M20), .A0_f (new_AGEMA_signal_9155), .A1_t (new_AGEMA_signal_9156), .A1_f (new_AGEMA_signal_9157), .B0_t (SubBytesIns_Inst_Sbox_14_M23), .B0_f (new_AGEMA_signal_9392), .B1_t (new_AGEMA_signal_9393), .B1_f (new_AGEMA_signal_9394), .Z0_t (SubBytesIns_Inst_Sbox_14_M31), .Z0_f (new_AGEMA_signal_9695), .Z1_t (new_AGEMA_signal_9696), .Z1_f (new_AGEMA_signal_9697) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M27), .A0_f (new_AGEMA_signal_9398), .A1_t (new_AGEMA_signal_9399), .A1_f (new_AGEMA_signal_9400), .B0_t (SubBytesIns_Inst_Sbox_14_M31), .B0_f (new_AGEMA_signal_9695), .B1_t (new_AGEMA_signal_9696), .B1_f (new_AGEMA_signal_9697), .Z0_t (SubBytesIns_Inst_Sbox_14_M32), .Z0_f (new_AGEMA_signal_9992), .Z1_t (new_AGEMA_signal_9993), .Z1_f (new_AGEMA_signal_9994) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M27), .A0_f (new_AGEMA_signal_9398), .A1_t (new_AGEMA_signal_9399), .A1_f (new_AGEMA_signal_9400), .B0_t (SubBytesIns_Inst_Sbox_14_M25), .B0_f (new_AGEMA_signal_9395), .B1_t (new_AGEMA_signal_9396), .B1_f (new_AGEMA_signal_9397), .Z0_t (SubBytesIns_Inst_Sbox_14_M33), .Z0_f (new_AGEMA_signal_9698), .Z1_t (new_AGEMA_signal_9699), .Z1_f (new_AGEMA_signal_9700) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M21), .A0_f (new_AGEMA_signal_9158), .A1_t (new_AGEMA_signal_9159), .A1_f (new_AGEMA_signal_9160), .B0_t (SubBytesIns_Inst_Sbox_14_M22), .B0_f (new_AGEMA_signal_9161), .B1_t (new_AGEMA_signal_9162), .B1_f (new_AGEMA_signal_9163), .Z0_t (SubBytesIns_Inst_Sbox_14_M34), .Z0_f (new_AGEMA_signal_9401), .Z1_t (new_AGEMA_signal_9402), .Z1_f (new_AGEMA_signal_9403) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M24), .A0_f (new_AGEMA_signal_9686), .A1_t (new_AGEMA_signal_9687), .A1_f (new_AGEMA_signal_9688), .B0_t (SubBytesIns_Inst_Sbox_14_M34), .B0_f (new_AGEMA_signal_9401), .B1_t (new_AGEMA_signal_9402), .B1_f (new_AGEMA_signal_9403), .Z0_t (SubBytesIns_Inst_Sbox_14_M35), .Z0_f (new_AGEMA_signal_9995), .Z1_t (new_AGEMA_signal_9996), .Z1_f (new_AGEMA_signal_9997) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M24), .A0_f (new_AGEMA_signal_9686), .A1_t (new_AGEMA_signal_9687), .A1_f (new_AGEMA_signal_9688), .B0_t (SubBytesIns_Inst_Sbox_14_M25), .B0_f (new_AGEMA_signal_9395), .B1_t (new_AGEMA_signal_9396), .B1_f (new_AGEMA_signal_9397), .Z0_t (SubBytesIns_Inst_Sbox_14_M36), .Z0_f (new_AGEMA_signal_9998), .Z1_t (new_AGEMA_signal_9999), .Z1_f (new_AGEMA_signal_10000) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M21), .A0_f (new_AGEMA_signal_9158), .A1_t (new_AGEMA_signal_9159), .A1_f (new_AGEMA_signal_9160), .B0_t (SubBytesIns_Inst_Sbox_14_M29), .B0_f (new_AGEMA_signal_9986), .B1_t (new_AGEMA_signal_9987), .B1_f (new_AGEMA_signal_9988), .Z0_t (SubBytesIns_Inst_Sbox_14_M37), .Z0_f (new_AGEMA_signal_10232), .Z1_t (new_AGEMA_signal_10233), .Z1_f (new_AGEMA_signal_10234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M32), .A0_f (new_AGEMA_signal_9992), .A1_t (new_AGEMA_signal_9993), .A1_f (new_AGEMA_signal_9994), .B0_t (SubBytesIns_Inst_Sbox_14_M33), .B0_f (new_AGEMA_signal_9698), .B1_t (new_AGEMA_signal_9699), .B1_f (new_AGEMA_signal_9700), .Z0_t (SubBytesIns_Inst_Sbox_14_M38), .Z0_f (new_AGEMA_signal_10235), .Z1_t (new_AGEMA_signal_10236), .Z1_f (new_AGEMA_signal_10237) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M23), .A0_f (new_AGEMA_signal_9392), .A1_t (new_AGEMA_signal_9393), .A1_f (new_AGEMA_signal_9394), .B0_t (SubBytesIns_Inst_Sbox_14_M30), .B0_f (new_AGEMA_signal_9989), .B1_t (new_AGEMA_signal_9990), .B1_f (new_AGEMA_signal_9991), .Z0_t (SubBytesIns_Inst_Sbox_14_M39), .Z0_f (new_AGEMA_signal_10238), .Z1_t (new_AGEMA_signal_10239), .Z1_f (new_AGEMA_signal_10240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M35), .A0_f (new_AGEMA_signal_9995), .A1_t (new_AGEMA_signal_9996), .A1_f (new_AGEMA_signal_9997), .B0_t (SubBytesIns_Inst_Sbox_14_M36), .B0_f (new_AGEMA_signal_9998), .B1_t (new_AGEMA_signal_9999), .B1_f (new_AGEMA_signal_10000), .Z0_t (SubBytesIns_Inst_Sbox_14_M40), .Z0_f (new_AGEMA_signal_10241), .Z1_t (new_AGEMA_signal_10242), .Z1_f (new_AGEMA_signal_10243) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M38), .A0_f (new_AGEMA_signal_10235), .A1_t (new_AGEMA_signal_10236), .A1_f (new_AGEMA_signal_10237), .B0_t (SubBytesIns_Inst_Sbox_14_M40), .B0_f (new_AGEMA_signal_10241), .B1_t (new_AGEMA_signal_10242), .B1_f (new_AGEMA_signal_10243), .Z0_t (SubBytesIns_Inst_Sbox_14_M41), .Z0_f (new_AGEMA_signal_10904), .Z1_t (new_AGEMA_signal_10905), .Z1_f (new_AGEMA_signal_10906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M37), .A0_f (new_AGEMA_signal_10232), .A1_t (new_AGEMA_signal_10233), .A1_f (new_AGEMA_signal_10234), .B0_t (SubBytesIns_Inst_Sbox_14_M39), .B0_f (new_AGEMA_signal_10238), .B1_t (new_AGEMA_signal_10239), .B1_f (new_AGEMA_signal_10240), .Z0_t (SubBytesIns_Inst_Sbox_14_M42), .Z0_f (new_AGEMA_signal_10907), .Z1_t (new_AGEMA_signal_10908), .Z1_f (new_AGEMA_signal_10909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M37), .A0_f (new_AGEMA_signal_10232), .A1_t (new_AGEMA_signal_10233), .A1_f (new_AGEMA_signal_10234), .B0_t (SubBytesIns_Inst_Sbox_14_M38), .B0_f (new_AGEMA_signal_10235), .B1_t (new_AGEMA_signal_10236), .B1_f (new_AGEMA_signal_10237), .Z0_t (SubBytesIns_Inst_Sbox_14_M43), .Z0_f (new_AGEMA_signal_10910), .Z1_t (new_AGEMA_signal_10911), .Z1_f (new_AGEMA_signal_10912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M39), .A0_f (new_AGEMA_signal_10238), .A1_t (new_AGEMA_signal_10239), .A1_f (new_AGEMA_signal_10240), .B0_t (SubBytesIns_Inst_Sbox_14_M40), .B0_f (new_AGEMA_signal_10241), .B1_t (new_AGEMA_signal_10242), .B1_f (new_AGEMA_signal_10243), .Z0_t (SubBytesIns_Inst_Sbox_14_M44), .Z0_f (new_AGEMA_signal_10913), .Z1_t (new_AGEMA_signal_10914), .Z1_f (new_AGEMA_signal_10915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M42), .A0_f (new_AGEMA_signal_10907), .A1_t (new_AGEMA_signal_10908), .A1_f (new_AGEMA_signal_10909), .B0_t (SubBytesIns_Inst_Sbox_14_M41), .B0_f (new_AGEMA_signal_10904), .B1_t (new_AGEMA_signal_10905), .B1_f (new_AGEMA_signal_10906), .Z0_t (SubBytesIns_Inst_Sbox_14_M45), .Z0_f (new_AGEMA_signal_11624), .Z1_t (new_AGEMA_signal_11625), .Z1_f (new_AGEMA_signal_11626) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M44), .A0_f (new_AGEMA_signal_10913), .A1_t (new_AGEMA_signal_10914), .A1_f (new_AGEMA_signal_10915), .B0_t (SubBytesIns_Inst_Sbox_14_T6), .B0_f (new_AGEMA_signal_7264), .B1_t (new_AGEMA_signal_7265), .B1_f (new_AGEMA_signal_7266), .Z0_t (SubBytesIns_Inst_Sbox_14_M46), .Z0_f (new_AGEMA_signal_11627), .Z1_t (new_AGEMA_signal_11628), .Z1_f (new_AGEMA_signal_11629) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M40), .A0_f (new_AGEMA_signal_10241), .A1_t (new_AGEMA_signal_10242), .A1_f (new_AGEMA_signal_10243), .B0_t (SubBytesIns_Inst_Sbox_14_T8), .B0_f (new_AGEMA_signal_8018), .B1_t (new_AGEMA_signal_8019), .B1_f (new_AGEMA_signal_8020), .Z0_t (SubBytesIns_Inst_Sbox_14_M47), .Z0_f (new_AGEMA_signal_10916), .Z1_t (new_AGEMA_signal_10917), .Z1_f (new_AGEMA_signal_10918) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M39), .A0_f (new_AGEMA_signal_10238), .A1_t (new_AGEMA_signal_10239), .A1_f (new_AGEMA_signal_10240), .B0_t (ciphertext_s0_t[112]), .B0_f (ciphertext_s0_f[112]), .B1_t (ciphertext_s1_t[112]), .B1_f (ciphertext_s1_f[112]), .Z0_t (SubBytesIns_Inst_Sbox_14_M48), .Z0_f (new_AGEMA_signal_10919), .Z1_t (new_AGEMA_signal_10920), .Z1_f (new_AGEMA_signal_10921) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M43), .A0_f (new_AGEMA_signal_10910), .A1_t (new_AGEMA_signal_10911), .A1_f (new_AGEMA_signal_10912), .B0_t (SubBytesIns_Inst_Sbox_14_T16), .B0_f (new_AGEMA_signal_7276), .B1_t (new_AGEMA_signal_7277), .B1_f (new_AGEMA_signal_7278), .Z0_t (SubBytesIns_Inst_Sbox_14_M49), .Z0_f (new_AGEMA_signal_11630), .Z1_t (new_AGEMA_signal_11631), .Z1_f (new_AGEMA_signal_11632) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M38), .A0_f (new_AGEMA_signal_10235), .A1_t (new_AGEMA_signal_10236), .A1_f (new_AGEMA_signal_10237), .B0_t (SubBytesIns_Inst_Sbox_14_T9), .B0_f (new_AGEMA_signal_7267), .B1_t (new_AGEMA_signal_7268), .B1_f (new_AGEMA_signal_7269), .Z0_t (SubBytesIns_Inst_Sbox_14_M50), .Z0_f (new_AGEMA_signal_10922), .Z1_t (new_AGEMA_signal_10923), .Z1_f (new_AGEMA_signal_10924) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M37), .A0_f (new_AGEMA_signal_10232), .A1_t (new_AGEMA_signal_10233), .A1_f (new_AGEMA_signal_10234), .B0_t (SubBytesIns_Inst_Sbox_14_T17), .B0_f (new_AGEMA_signal_8027), .B1_t (new_AGEMA_signal_8028), .B1_f (new_AGEMA_signal_8029), .Z0_t (SubBytesIns_Inst_Sbox_14_M51), .Z0_f (new_AGEMA_signal_10925), .Z1_t (new_AGEMA_signal_10926), .Z1_f (new_AGEMA_signal_10927) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M42), .A0_f (new_AGEMA_signal_10907), .A1_t (new_AGEMA_signal_10908), .A1_f (new_AGEMA_signal_10909), .B0_t (SubBytesIns_Inst_Sbox_14_T15), .B0_f (new_AGEMA_signal_7273), .B1_t (new_AGEMA_signal_7274), .B1_f (new_AGEMA_signal_7275), .Z0_t (SubBytesIns_Inst_Sbox_14_M52), .Z0_f (new_AGEMA_signal_11633), .Z1_t (new_AGEMA_signal_11634), .Z1_f (new_AGEMA_signal_11635) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M45), .A0_f (new_AGEMA_signal_11624), .A1_t (new_AGEMA_signal_11625), .A1_f (new_AGEMA_signal_11626), .B0_t (SubBytesIns_Inst_Sbox_14_T27), .B0_f (new_AGEMA_signal_7285), .B1_t (new_AGEMA_signal_7286), .B1_f (new_AGEMA_signal_7287), .Z0_t (SubBytesIns_Inst_Sbox_14_M53), .Z0_f (new_AGEMA_signal_12236), .Z1_t (new_AGEMA_signal_12237), .Z1_f (new_AGEMA_signal_12238) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M41), .A0_f (new_AGEMA_signal_10904), .A1_t (new_AGEMA_signal_10905), .A1_f (new_AGEMA_signal_10906), .B0_t (SubBytesIns_Inst_Sbox_14_T10), .B0_f (new_AGEMA_signal_8021), .B1_t (new_AGEMA_signal_8022), .B1_f (new_AGEMA_signal_8023), .Z0_t (SubBytesIns_Inst_Sbox_14_M54), .Z0_f (new_AGEMA_signal_11636), .Z1_t (new_AGEMA_signal_11637), .Z1_f (new_AGEMA_signal_11638) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M44), .A0_f (new_AGEMA_signal_10913), .A1_t (new_AGEMA_signal_10914), .A1_f (new_AGEMA_signal_10915), .B0_t (SubBytesIns_Inst_Sbox_14_T13), .B0_f (new_AGEMA_signal_7270), .B1_t (new_AGEMA_signal_7271), .B1_f (new_AGEMA_signal_7272), .Z0_t (SubBytesIns_Inst_Sbox_14_M55), .Z0_f (new_AGEMA_signal_11639), .Z1_t (new_AGEMA_signal_11640), .Z1_f (new_AGEMA_signal_11641) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M40), .A0_f (new_AGEMA_signal_10241), .A1_t (new_AGEMA_signal_10242), .A1_f (new_AGEMA_signal_10243), .B0_t (SubBytesIns_Inst_Sbox_14_T23), .B0_f (new_AGEMA_signal_8033), .B1_t (new_AGEMA_signal_8034), .B1_f (new_AGEMA_signal_8035), .Z0_t (SubBytesIns_Inst_Sbox_14_M56), .Z0_f (new_AGEMA_signal_10928), .Z1_t (new_AGEMA_signal_10929), .Z1_f (new_AGEMA_signal_10930) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M39), .A0_f (new_AGEMA_signal_10238), .A1_t (new_AGEMA_signal_10239), .A1_f (new_AGEMA_signal_10240), .B0_t (SubBytesIns_Inst_Sbox_14_T19), .B0_f (new_AGEMA_signal_7279), .B1_t (new_AGEMA_signal_7280), .B1_f (new_AGEMA_signal_7281), .Z0_t (SubBytesIns_Inst_Sbox_14_M57), .Z0_f (new_AGEMA_signal_10931), .Z1_t (new_AGEMA_signal_10932), .Z1_f (new_AGEMA_signal_10933) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M43), .A0_f (new_AGEMA_signal_10910), .A1_t (new_AGEMA_signal_10911), .A1_f (new_AGEMA_signal_10912), .B0_t (SubBytesIns_Inst_Sbox_14_T3), .B0_f (new_AGEMA_signal_6772), .B1_t (new_AGEMA_signal_6773), .B1_f (new_AGEMA_signal_6774), .Z0_t (SubBytesIns_Inst_Sbox_14_M58), .Z0_f (new_AGEMA_signal_11642), .Z1_t (new_AGEMA_signal_11643), .Z1_f (new_AGEMA_signal_11644) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M38), .A0_f (new_AGEMA_signal_10235), .A1_t (new_AGEMA_signal_10236), .A1_f (new_AGEMA_signal_10237), .B0_t (SubBytesIns_Inst_Sbox_14_T22), .B0_f (new_AGEMA_signal_7282), .B1_t (new_AGEMA_signal_7283), .B1_f (new_AGEMA_signal_7284), .Z0_t (SubBytesIns_Inst_Sbox_14_M59), .Z0_f (new_AGEMA_signal_10934), .Z1_t (new_AGEMA_signal_10935), .Z1_f (new_AGEMA_signal_10936) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M37), .A0_f (new_AGEMA_signal_10232), .A1_t (new_AGEMA_signal_10233), .A1_f (new_AGEMA_signal_10234), .B0_t (SubBytesIns_Inst_Sbox_14_T20), .B0_f (new_AGEMA_signal_8030), .B1_t (new_AGEMA_signal_8031), .B1_f (new_AGEMA_signal_8032), .Z0_t (SubBytesIns_Inst_Sbox_14_M60), .Z0_f (new_AGEMA_signal_10937), .Z1_t (new_AGEMA_signal_10938), .Z1_f (new_AGEMA_signal_10939) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M42), .A0_f (new_AGEMA_signal_10907), .A1_t (new_AGEMA_signal_10908), .A1_f (new_AGEMA_signal_10909), .B0_t (SubBytesIns_Inst_Sbox_14_T1), .B0_f (new_AGEMA_signal_6766), .B1_t (new_AGEMA_signal_6767), .B1_f (new_AGEMA_signal_6768), .Z0_t (SubBytesIns_Inst_Sbox_14_M61), .Z0_f (new_AGEMA_signal_11645), .Z1_t (new_AGEMA_signal_11646), .Z1_f (new_AGEMA_signal_11647) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M45), .A0_f (new_AGEMA_signal_11624), .A1_t (new_AGEMA_signal_11625), .A1_f (new_AGEMA_signal_11626), .B0_t (SubBytesIns_Inst_Sbox_14_T4), .B0_f (new_AGEMA_signal_6775), .B1_t (new_AGEMA_signal_6776), .B1_f (new_AGEMA_signal_6777), .Z0_t (SubBytesIns_Inst_Sbox_14_M62), .Z0_f (new_AGEMA_signal_12239), .Z1_t (new_AGEMA_signal_12240), .Z1_f (new_AGEMA_signal_12241) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M41), .A0_f (new_AGEMA_signal_10904), .A1_t (new_AGEMA_signal_10905), .A1_f (new_AGEMA_signal_10906), .B0_t (SubBytesIns_Inst_Sbox_14_T2), .B0_f (new_AGEMA_signal_6769), .B1_t (new_AGEMA_signal_6770), .B1_f (new_AGEMA_signal_6771), .Z0_t (SubBytesIns_Inst_Sbox_14_M63), .Z0_f (new_AGEMA_signal_11648), .Z1_t (new_AGEMA_signal_11649), .Z1_f (new_AGEMA_signal_11650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M61), .A0_f (new_AGEMA_signal_11645), .A1_t (new_AGEMA_signal_11646), .A1_f (new_AGEMA_signal_11647), .B0_t (SubBytesIns_Inst_Sbox_14_M62), .B0_f (new_AGEMA_signal_12239), .B1_t (new_AGEMA_signal_12240), .B1_f (new_AGEMA_signal_12241), .Z0_t (SubBytesIns_Inst_Sbox_14_L0), .Z0_f (new_AGEMA_signal_12782), .Z1_t (new_AGEMA_signal_12783), .Z1_f (new_AGEMA_signal_12784) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M50), .A0_f (new_AGEMA_signal_10922), .A1_t (new_AGEMA_signal_10923), .A1_f (new_AGEMA_signal_10924), .B0_t (SubBytesIns_Inst_Sbox_14_M56), .B0_f (new_AGEMA_signal_10928), .B1_t (new_AGEMA_signal_10929), .B1_f (new_AGEMA_signal_10930), .Z0_t (SubBytesIns_Inst_Sbox_14_L1), .Z0_f (new_AGEMA_signal_11651), .Z1_t (new_AGEMA_signal_11652), .Z1_f (new_AGEMA_signal_11653) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M46), .A0_f (new_AGEMA_signal_11627), .A1_t (new_AGEMA_signal_11628), .A1_f (new_AGEMA_signal_11629), .B0_t (SubBytesIns_Inst_Sbox_14_M48), .B0_f (new_AGEMA_signal_10919), .B1_t (new_AGEMA_signal_10920), .B1_f (new_AGEMA_signal_10921), .Z0_t (SubBytesIns_Inst_Sbox_14_L2), .Z0_f (new_AGEMA_signal_12242), .Z1_t (new_AGEMA_signal_12243), .Z1_f (new_AGEMA_signal_12244) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M47), .A0_f (new_AGEMA_signal_10916), .A1_t (new_AGEMA_signal_10917), .A1_f (new_AGEMA_signal_10918), .B0_t (SubBytesIns_Inst_Sbox_14_M55), .B0_f (new_AGEMA_signal_11639), .B1_t (new_AGEMA_signal_11640), .B1_f (new_AGEMA_signal_11641), .Z0_t (SubBytesIns_Inst_Sbox_14_L3), .Z0_f (new_AGEMA_signal_12245), .Z1_t (new_AGEMA_signal_12246), .Z1_f (new_AGEMA_signal_12247) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M54), .A0_f (new_AGEMA_signal_11636), .A1_t (new_AGEMA_signal_11637), .A1_f (new_AGEMA_signal_11638), .B0_t (SubBytesIns_Inst_Sbox_14_M58), .B0_f (new_AGEMA_signal_11642), .B1_t (new_AGEMA_signal_11643), .B1_f (new_AGEMA_signal_11644), .Z0_t (SubBytesIns_Inst_Sbox_14_L4), .Z0_f (new_AGEMA_signal_12248), .Z1_t (new_AGEMA_signal_12249), .Z1_f (new_AGEMA_signal_12250) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M49), .A0_f (new_AGEMA_signal_11630), .A1_t (new_AGEMA_signal_11631), .A1_f (new_AGEMA_signal_11632), .B0_t (SubBytesIns_Inst_Sbox_14_M61), .B0_f (new_AGEMA_signal_11645), .B1_t (new_AGEMA_signal_11646), .B1_f (new_AGEMA_signal_11647), .Z0_t (SubBytesIns_Inst_Sbox_14_L5), .Z0_f (new_AGEMA_signal_12251), .Z1_t (new_AGEMA_signal_12252), .Z1_f (new_AGEMA_signal_12253) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M62), .A0_f (new_AGEMA_signal_12239), .A1_t (new_AGEMA_signal_12240), .A1_f (new_AGEMA_signal_12241), .B0_t (SubBytesIns_Inst_Sbox_14_L5), .B0_f (new_AGEMA_signal_12251), .B1_t (new_AGEMA_signal_12252), .B1_f (new_AGEMA_signal_12253), .Z0_t (SubBytesIns_Inst_Sbox_14_L6), .Z0_f (new_AGEMA_signal_12785), .Z1_t (new_AGEMA_signal_12786), .Z1_f (new_AGEMA_signal_12787) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M46), .A0_f (new_AGEMA_signal_11627), .A1_t (new_AGEMA_signal_11628), .A1_f (new_AGEMA_signal_11629), .B0_t (SubBytesIns_Inst_Sbox_14_L3), .B0_f (new_AGEMA_signal_12245), .B1_t (new_AGEMA_signal_12246), .B1_f (new_AGEMA_signal_12247), .Z0_t (SubBytesIns_Inst_Sbox_14_L7), .Z0_f (new_AGEMA_signal_12788), .Z1_t (new_AGEMA_signal_12789), .Z1_f (new_AGEMA_signal_12790) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M51), .A0_f (new_AGEMA_signal_10925), .A1_t (new_AGEMA_signal_10926), .A1_f (new_AGEMA_signal_10927), .B0_t (SubBytesIns_Inst_Sbox_14_M59), .B0_f (new_AGEMA_signal_10934), .B1_t (new_AGEMA_signal_10935), .B1_f (new_AGEMA_signal_10936), .Z0_t (SubBytesIns_Inst_Sbox_14_L8), .Z0_f (new_AGEMA_signal_11654), .Z1_t (new_AGEMA_signal_11655), .Z1_f (new_AGEMA_signal_11656) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M52), .A0_f (new_AGEMA_signal_11633), .A1_t (new_AGEMA_signal_11634), .A1_f (new_AGEMA_signal_11635), .B0_t (SubBytesIns_Inst_Sbox_14_M53), .B0_f (new_AGEMA_signal_12236), .B1_t (new_AGEMA_signal_12237), .B1_f (new_AGEMA_signal_12238), .Z0_t (SubBytesIns_Inst_Sbox_14_L9), .Z0_f (new_AGEMA_signal_12791), .Z1_t (new_AGEMA_signal_12792), .Z1_f (new_AGEMA_signal_12793) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M53), .A0_f (new_AGEMA_signal_12236), .A1_t (new_AGEMA_signal_12237), .A1_f (new_AGEMA_signal_12238), .B0_t (SubBytesIns_Inst_Sbox_14_L4), .B0_f (new_AGEMA_signal_12248), .B1_t (new_AGEMA_signal_12249), .B1_f (new_AGEMA_signal_12250), .Z0_t (SubBytesIns_Inst_Sbox_14_L10), .Z0_f (new_AGEMA_signal_12794), .Z1_t (new_AGEMA_signal_12795), .Z1_f (new_AGEMA_signal_12796) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M60), .A0_f (new_AGEMA_signal_10937), .A1_t (new_AGEMA_signal_10938), .A1_f (new_AGEMA_signal_10939), .B0_t (SubBytesIns_Inst_Sbox_14_L2), .B0_f (new_AGEMA_signal_12242), .B1_t (new_AGEMA_signal_12243), .B1_f (new_AGEMA_signal_12244), .Z0_t (SubBytesIns_Inst_Sbox_14_L11), .Z0_f (new_AGEMA_signal_12797), .Z1_t (new_AGEMA_signal_12798), .Z1_f (new_AGEMA_signal_12799) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M48), .A0_f (new_AGEMA_signal_10919), .A1_t (new_AGEMA_signal_10920), .A1_f (new_AGEMA_signal_10921), .B0_t (SubBytesIns_Inst_Sbox_14_M51), .B0_f (new_AGEMA_signal_10925), .B1_t (new_AGEMA_signal_10926), .B1_f (new_AGEMA_signal_10927), .Z0_t (SubBytesIns_Inst_Sbox_14_L12), .Z0_f (new_AGEMA_signal_11657), .Z1_t (new_AGEMA_signal_11658), .Z1_f (new_AGEMA_signal_11659) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M50), .A0_f (new_AGEMA_signal_10922), .A1_t (new_AGEMA_signal_10923), .A1_f (new_AGEMA_signal_10924), .B0_t (SubBytesIns_Inst_Sbox_14_L0), .B0_f (new_AGEMA_signal_12782), .B1_t (new_AGEMA_signal_12783), .B1_f (new_AGEMA_signal_12784), .Z0_t (SubBytesIns_Inst_Sbox_14_L13), .Z0_f (new_AGEMA_signal_13430), .Z1_t (new_AGEMA_signal_13431), .Z1_f (new_AGEMA_signal_13432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M52), .A0_f (new_AGEMA_signal_11633), .A1_t (new_AGEMA_signal_11634), .A1_f (new_AGEMA_signal_11635), .B0_t (SubBytesIns_Inst_Sbox_14_M61), .B0_f (new_AGEMA_signal_11645), .B1_t (new_AGEMA_signal_11646), .B1_f (new_AGEMA_signal_11647), .Z0_t (SubBytesIns_Inst_Sbox_14_L14), .Z0_f (new_AGEMA_signal_12254), .Z1_t (new_AGEMA_signal_12255), .Z1_f (new_AGEMA_signal_12256) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M55), .A0_f (new_AGEMA_signal_11639), .A1_t (new_AGEMA_signal_11640), .A1_f (new_AGEMA_signal_11641), .B0_t (SubBytesIns_Inst_Sbox_14_L1), .B0_f (new_AGEMA_signal_11651), .B1_t (new_AGEMA_signal_11652), .B1_f (new_AGEMA_signal_11653), .Z0_t (SubBytesIns_Inst_Sbox_14_L15), .Z0_f (new_AGEMA_signal_12257), .Z1_t (new_AGEMA_signal_12258), .Z1_f (new_AGEMA_signal_12259) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M56), .A0_f (new_AGEMA_signal_10928), .A1_t (new_AGEMA_signal_10929), .A1_f (new_AGEMA_signal_10930), .B0_t (SubBytesIns_Inst_Sbox_14_L0), .B0_f (new_AGEMA_signal_12782), .B1_t (new_AGEMA_signal_12783), .B1_f (new_AGEMA_signal_12784), .Z0_t (SubBytesIns_Inst_Sbox_14_L16), .Z0_f (new_AGEMA_signal_13433), .Z1_t (new_AGEMA_signal_13434), .Z1_f (new_AGEMA_signal_13435) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M57), .A0_f (new_AGEMA_signal_10931), .A1_t (new_AGEMA_signal_10932), .A1_f (new_AGEMA_signal_10933), .B0_t (SubBytesIns_Inst_Sbox_14_L1), .B0_f (new_AGEMA_signal_11651), .B1_t (new_AGEMA_signal_11652), .B1_f (new_AGEMA_signal_11653), .Z0_t (SubBytesIns_Inst_Sbox_14_L17), .Z0_f (new_AGEMA_signal_12260), .Z1_t (new_AGEMA_signal_12261), .Z1_f (new_AGEMA_signal_12262) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M58), .A0_f (new_AGEMA_signal_11642), .A1_t (new_AGEMA_signal_11643), .A1_f (new_AGEMA_signal_11644), .B0_t (SubBytesIns_Inst_Sbox_14_L8), .B0_f (new_AGEMA_signal_11654), .B1_t (new_AGEMA_signal_11655), .B1_f (new_AGEMA_signal_11656), .Z0_t (SubBytesIns_Inst_Sbox_14_L18), .Z0_f (new_AGEMA_signal_12263), .Z1_t (new_AGEMA_signal_12264), .Z1_f (new_AGEMA_signal_12265) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M63), .A0_f (new_AGEMA_signal_11648), .A1_t (new_AGEMA_signal_11649), .A1_f (new_AGEMA_signal_11650), .B0_t (SubBytesIns_Inst_Sbox_14_L4), .B0_f (new_AGEMA_signal_12248), .B1_t (new_AGEMA_signal_12249), .B1_f (new_AGEMA_signal_12250), .Z0_t (SubBytesIns_Inst_Sbox_14_L19), .Z0_f (new_AGEMA_signal_12800), .Z1_t (new_AGEMA_signal_12801), .Z1_f (new_AGEMA_signal_12802) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L0), .A0_f (new_AGEMA_signal_12782), .A1_t (new_AGEMA_signal_12783), .A1_f (new_AGEMA_signal_12784), .B0_t (SubBytesIns_Inst_Sbox_14_L1), .B0_f (new_AGEMA_signal_11651), .B1_t (new_AGEMA_signal_11652), .B1_f (new_AGEMA_signal_11653), .Z0_t (SubBytesIns_Inst_Sbox_14_L20), .Z0_f (new_AGEMA_signal_13436), .Z1_t (new_AGEMA_signal_13437), .Z1_f (new_AGEMA_signal_13438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L1), .A0_f (new_AGEMA_signal_11651), .A1_t (new_AGEMA_signal_11652), .A1_f (new_AGEMA_signal_11653), .B0_t (SubBytesIns_Inst_Sbox_14_L7), .B0_f (new_AGEMA_signal_12788), .B1_t (new_AGEMA_signal_12789), .B1_f (new_AGEMA_signal_12790), .Z0_t (SubBytesIns_Inst_Sbox_14_L21), .Z0_f (new_AGEMA_signal_13439), .Z1_t (new_AGEMA_signal_13440), .Z1_f (new_AGEMA_signal_13441) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L3), .A0_f (new_AGEMA_signal_12245), .A1_t (new_AGEMA_signal_12246), .A1_f (new_AGEMA_signal_12247), .B0_t (SubBytesIns_Inst_Sbox_14_L12), .B0_f (new_AGEMA_signal_11657), .B1_t (new_AGEMA_signal_11658), .B1_f (new_AGEMA_signal_11659), .Z0_t (SubBytesIns_Inst_Sbox_14_L22), .Z0_f (new_AGEMA_signal_12803), .Z1_t (new_AGEMA_signal_12804), .Z1_f (new_AGEMA_signal_12805) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L18), .A0_f (new_AGEMA_signal_12263), .A1_t (new_AGEMA_signal_12264), .A1_f (new_AGEMA_signal_12265), .B0_t (SubBytesIns_Inst_Sbox_14_L2), .B0_f (new_AGEMA_signal_12242), .B1_t (new_AGEMA_signal_12243), .B1_f (new_AGEMA_signal_12244), .Z0_t (SubBytesIns_Inst_Sbox_14_L23), .Z0_f (new_AGEMA_signal_12806), .Z1_t (new_AGEMA_signal_12807), .Z1_f (new_AGEMA_signal_12808) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L15), .A0_f (new_AGEMA_signal_12257), .A1_t (new_AGEMA_signal_12258), .A1_f (new_AGEMA_signal_12259), .B0_t (SubBytesIns_Inst_Sbox_14_L9), .B0_f (new_AGEMA_signal_12791), .B1_t (new_AGEMA_signal_12792), .B1_f (new_AGEMA_signal_12793), .Z0_t (SubBytesIns_Inst_Sbox_14_L24), .Z0_f (new_AGEMA_signal_13442), .Z1_t (new_AGEMA_signal_13443), .Z1_f (new_AGEMA_signal_13444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L6), .A0_f (new_AGEMA_signal_12785), .A1_t (new_AGEMA_signal_12786), .A1_f (new_AGEMA_signal_12787), .B0_t (SubBytesIns_Inst_Sbox_14_L10), .B0_f (new_AGEMA_signal_12794), .B1_t (new_AGEMA_signal_12795), .B1_f (new_AGEMA_signal_12796), .Z0_t (SubBytesIns_Inst_Sbox_14_L25), .Z0_f (new_AGEMA_signal_13445), .Z1_t (new_AGEMA_signal_13446), .Z1_f (new_AGEMA_signal_13447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L7), .A0_f (new_AGEMA_signal_12788), .A1_t (new_AGEMA_signal_12789), .A1_f (new_AGEMA_signal_12790), .B0_t (SubBytesIns_Inst_Sbox_14_L9), .B0_f (new_AGEMA_signal_12791), .B1_t (new_AGEMA_signal_12792), .B1_f (new_AGEMA_signal_12793), .Z0_t (SubBytesIns_Inst_Sbox_14_L26), .Z0_f (new_AGEMA_signal_13448), .Z1_t (new_AGEMA_signal_13449), .Z1_f (new_AGEMA_signal_13450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L8), .A0_f (new_AGEMA_signal_11654), .A1_t (new_AGEMA_signal_11655), .A1_f (new_AGEMA_signal_11656), .B0_t (SubBytesIns_Inst_Sbox_14_L10), .B0_f (new_AGEMA_signal_12794), .B1_t (new_AGEMA_signal_12795), .B1_f (new_AGEMA_signal_12796), .Z0_t (SubBytesIns_Inst_Sbox_14_L27), .Z0_f (new_AGEMA_signal_13451), .Z1_t (new_AGEMA_signal_13452), .Z1_f (new_AGEMA_signal_13453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L11), .A0_f (new_AGEMA_signal_12797), .A1_t (new_AGEMA_signal_12798), .A1_f (new_AGEMA_signal_12799), .B0_t (SubBytesIns_Inst_Sbox_14_L14), .B0_f (new_AGEMA_signal_12254), .B1_t (new_AGEMA_signal_12255), .B1_f (new_AGEMA_signal_12256), .Z0_t (SubBytesIns_Inst_Sbox_14_L28), .Z0_f (new_AGEMA_signal_13454), .Z1_t (new_AGEMA_signal_13455), .Z1_f (new_AGEMA_signal_13456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L11), .A0_f (new_AGEMA_signal_12797), .A1_t (new_AGEMA_signal_12798), .A1_f (new_AGEMA_signal_12799), .B0_t (SubBytesIns_Inst_Sbox_14_L17), .B0_f (new_AGEMA_signal_12260), .B1_t (new_AGEMA_signal_12261), .B1_f (new_AGEMA_signal_12262), .Z0_t (SubBytesIns_Inst_Sbox_14_L29), .Z0_f (new_AGEMA_signal_13457), .Z1_t (new_AGEMA_signal_13458), .Z1_f (new_AGEMA_signal_13459) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L6), .A0_f (new_AGEMA_signal_12785), .A1_t (new_AGEMA_signal_12786), .A1_f (new_AGEMA_signal_12787), .B0_t (SubBytesIns_Inst_Sbox_14_L24), .B0_f (new_AGEMA_signal_13442), .B1_t (new_AGEMA_signal_13443), .B1_f (new_AGEMA_signal_13444), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .Z0_f (new_AGEMA_signal_13934), .Z1_t (new_AGEMA_signal_13935), .Z1_f (new_AGEMA_signal_13936) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L16), .A0_f (new_AGEMA_signal_13433), .A1_t (new_AGEMA_signal_13434), .A1_f (new_AGEMA_signal_13435), .B0_t (SubBytesIns_Inst_Sbox_14_L26), .B0_f (new_AGEMA_signal_13448), .B1_t (new_AGEMA_signal_13449), .B1_f (new_AGEMA_signal_13450), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .Z0_f (new_AGEMA_signal_13937), .Z1_t (new_AGEMA_signal_13938), .Z1_f (new_AGEMA_signal_13939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L19), .A0_f (new_AGEMA_signal_12800), .A1_t (new_AGEMA_signal_12801), .A1_f (new_AGEMA_signal_12802), .B0_t (SubBytesIns_Inst_Sbox_14_L28), .B0_f (new_AGEMA_signal_13454), .B1_t (new_AGEMA_signal_13455), .B1_f (new_AGEMA_signal_13456), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .Z0_f (new_AGEMA_signal_13940), .Z1_t (new_AGEMA_signal_13941), .Z1_f (new_AGEMA_signal_13942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L6), .A0_f (new_AGEMA_signal_12785), .A1_t (new_AGEMA_signal_12786), .A1_f (new_AGEMA_signal_12787), .B0_t (SubBytesIns_Inst_Sbox_14_L21), .B0_f (new_AGEMA_signal_13439), .B1_t (new_AGEMA_signal_13440), .B1_f (new_AGEMA_signal_13441), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .Z0_f (new_AGEMA_signal_13943), .Z1_t (new_AGEMA_signal_13944), .Z1_f (new_AGEMA_signal_13945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L20), .A0_f (new_AGEMA_signal_13436), .A1_t (new_AGEMA_signal_13437), .A1_f (new_AGEMA_signal_13438), .B0_t (SubBytesIns_Inst_Sbox_14_L22), .B0_f (new_AGEMA_signal_12803), .B1_t (new_AGEMA_signal_12804), .B1_f (new_AGEMA_signal_12805), .Z0_t (MixColumnsInput[19]), .Z0_f (new_AGEMA_signal_13946), .Z1_t (new_AGEMA_signal_13947), .Z1_f (new_AGEMA_signal_13948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L25), .A0_f (new_AGEMA_signal_13445), .A1_t (new_AGEMA_signal_13446), .A1_f (new_AGEMA_signal_13447), .B0_t (SubBytesIns_Inst_Sbox_14_L29), .B0_f (new_AGEMA_signal_13457), .B1_t (new_AGEMA_signal_13458), .B1_f (new_AGEMA_signal_13459), .Z0_t (MixColumnsInput[18]), .Z0_f (new_AGEMA_signal_13949), .Z1_t (new_AGEMA_signal_13950), .Z1_f (new_AGEMA_signal_13951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L13), .A0_f (new_AGEMA_signal_13430), .A1_t (new_AGEMA_signal_13431), .A1_f (new_AGEMA_signal_13432), .B0_t (SubBytesIns_Inst_Sbox_14_L27), .B0_f (new_AGEMA_signal_13451), .B1_t (new_AGEMA_signal_13452), .B1_f (new_AGEMA_signal_13453), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .Z0_f (new_AGEMA_signal_13952), .Z1_t (new_AGEMA_signal_13953), .Z1_f (new_AGEMA_signal_13954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L6), .A0_f (new_AGEMA_signal_12785), .A1_t (new_AGEMA_signal_12786), .A1_f (new_AGEMA_signal_12787), .B0_t (SubBytesIns_Inst_Sbox_14_L23), .B0_f (new_AGEMA_signal_12806), .B1_t (new_AGEMA_signal_12807), .B1_f (new_AGEMA_signal_12808), .Z0_t (MixColumnsInput[16]), .Z0_f (new_AGEMA_signal_13460), .Z1_t (new_AGEMA_signal_13461), .Z1_f (new_AGEMA_signal_13462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T1_U1 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (ciphertext_s0_t[124]), .B0_f (ciphertext_s0_f[124]), .B1_t (ciphertext_s1_t[124]), .B1_f (ciphertext_s1_f[124]), .Z0_t (SubBytesIns_Inst_Sbox_15_T1), .Z0_f (new_AGEMA_signal_6796), .Z1_t (new_AGEMA_signal_6797), .Z1_f (new_AGEMA_signal_6798) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T2_U1 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (ciphertext_s0_t[122]), .B0_f (ciphertext_s0_f[122]), .B1_t (ciphertext_s1_t[122]), .B1_f (ciphertext_s1_f[122]), .Z0_t (SubBytesIns_Inst_Sbox_15_T2), .Z0_f (new_AGEMA_signal_6799), .Z1_t (new_AGEMA_signal_6800), .Z1_f (new_AGEMA_signal_6801) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T3_U1 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (ciphertext_s0_t[121]), .B0_f (ciphertext_s0_f[121]), .B1_t (ciphertext_s1_t[121]), .B1_f (ciphertext_s1_f[121]), .Z0_t (SubBytesIns_Inst_Sbox_15_T3), .Z0_f (new_AGEMA_signal_6802), .Z1_t (new_AGEMA_signal_6803), .Z1_f (new_AGEMA_signal_6804) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T4_U1 ( .A0_t (ciphertext_s0_t[124]), .A0_f (ciphertext_s0_f[124]), .A1_t (ciphertext_s1_t[124]), .A1_f (ciphertext_s1_f[124]), .B0_t (ciphertext_s0_t[122]), .B0_f (ciphertext_s0_f[122]), .B1_t (ciphertext_s1_t[122]), .B1_f (ciphertext_s1_f[122]), .Z0_t (SubBytesIns_Inst_Sbox_15_T4), .Z0_f (new_AGEMA_signal_6805), .Z1_t (new_AGEMA_signal_6806), .Z1_f (new_AGEMA_signal_6807) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T5_U1 ( .A0_t (ciphertext_s0_t[123]), .A0_f (ciphertext_s0_f[123]), .A1_t (ciphertext_s1_t[123]), .A1_f (ciphertext_s1_f[123]), .B0_t (ciphertext_s0_t[121]), .B0_f (ciphertext_s0_f[121]), .B1_t (ciphertext_s1_t[121]), .B1_f (ciphertext_s1_f[121]), .Z0_t (SubBytesIns_Inst_Sbox_15_T5), .Z0_f (new_AGEMA_signal_6808), .Z1_t (new_AGEMA_signal_6809), .Z1_f (new_AGEMA_signal_6810) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T1), .A0_f (new_AGEMA_signal_6796), .A1_t (new_AGEMA_signal_6797), .A1_f (new_AGEMA_signal_6798), .B0_t (SubBytesIns_Inst_Sbox_15_T5), .B0_f (new_AGEMA_signal_6808), .B1_t (new_AGEMA_signal_6809), .B1_f (new_AGEMA_signal_6810), .Z0_t (SubBytesIns_Inst_Sbox_15_T6), .Z0_f (new_AGEMA_signal_7288), .Z1_t (new_AGEMA_signal_7289), .Z1_f (new_AGEMA_signal_7290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T7_U1 ( .A0_t (ciphertext_s0_t[126]), .A0_f (ciphertext_s0_f[126]), .A1_t (ciphertext_s1_t[126]), .A1_f (ciphertext_s1_f[126]), .B0_t (ciphertext_s0_t[125]), .B0_f (ciphertext_s0_f[125]), .B1_t (ciphertext_s1_t[125]), .B1_f (ciphertext_s1_f[125]), .Z0_t (SubBytesIns_Inst_Sbox_15_T7), .Z0_f (new_AGEMA_signal_6811), .Z1_t (new_AGEMA_signal_6812), .Z1_f (new_AGEMA_signal_6813) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T8_U1 ( .A0_t (ciphertext_s0_t[120]), .A0_f (ciphertext_s0_f[120]), .A1_t (ciphertext_s1_t[120]), .A1_f (ciphertext_s1_f[120]), .B0_t (SubBytesIns_Inst_Sbox_15_T6), .B0_f (new_AGEMA_signal_7288), .B1_t (new_AGEMA_signal_7289), .B1_f (new_AGEMA_signal_7290), .Z0_t (SubBytesIns_Inst_Sbox_15_T8), .Z0_f (new_AGEMA_signal_8057), .Z1_t (new_AGEMA_signal_8058), .Z1_f (new_AGEMA_signal_8059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T9_U1 ( .A0_t (ciphertext_s0_t[120]), .A0_f (ciphertext_s0_f[120]), .A1_t (ciphertext_s1_t[120]), .A1_f (ciphertext_s1_f[120]), .B0_t (SubBytesIns_Inst_Sbox_15_T7), .B0_f (new_AGEMA_signal_6811), .B1_t (new_AGEMA_signal_6812), .B1_f (new_AGEMA_signal_6813), .Z0_t (SubBytesIns_Inst_Sbox_15_T9), .Z0_f (new_AGEMA_signal_7291), .Z1_t (new_AGEMA_signal_7292), .Z1_f (new_AGEMA_signal_7293) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T6), .A0_f (new_AGEMA_signal_7288), .A1_t (new_AGEMA_signal_7289), .A1_f (new_AGEMA_signal_7290), .B0_t (SubBytesIns_Inst_Sbox_15_T7), .B0_f (new_AGEMA_signal_6811), .B1_t (new_AGEMA_signal_6812), .B1_f (new_AGEMA_signal_6813), .Z0_t (SubBytesIns_Inst_Sbox_15_T10), .Z0_f (new_AGEMA_signal_8060), .Z1_t (new_AGEMA_signal_8061), .Z1_f (new_AGEMA_signal_8062) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T11_U1 ( .A0_t (ciphertext_s0_t[126]), .A0_f (ciphertext_s0_f[126]), .A1_t (ciphertext_s1_t[126]), .A1_f (ciphertext_s1_f[126]), .B0_t (ciphertext_s0_t[122]), .B0_f (ciphertext_s0_f[122]), .B1_t (ciphertext_s1_t[122]), .B1_f (ciphertext_s1_f[122]), .Z0_t (SubBytesIns_Inst_Sbox_15_T11), .Z0_f (new_AGEMA_signal_6814), .Z1_t (new_AGEMA_signal_6815), .Z1_f (new_AGEMA_signal_6816) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T12_U1 ( .A0_t (ciphertext_s0_t[125]), .A0_f (ciphertext_s0_f[125]), .A1_t (ciphertext_s1_t[125]), .A1_f (ciphertext_s1_f[125]), .B0_t (ciphertext_s0_t[122]), .B0_f (ciphertext_s0_f[122]), .B1_t (ciphertext_s1_t[122]), .B1_f (ciphertext_s1_f[122]), .Z0_t (SubBytesIns_Inst_Sbox_15_T12), .Z0_f (new_AGEMA_signal_6817), .Z1_t (new_AGEMA_signal_6818), .Z1_f (new_AGEMA_signal_6819) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T3), .A0_f (new_AGEMA_signal_6802), .A1_t (new_AGEMA_signal_6803), .A1_f (new_AGEMA_signal_6804), .B0_t (SubBytesIns_Inst_Sbox_15_T4), .B0_f (new_AGEMA_signal_6805), .B1_t (new_AGEMA_signal_6806), .B1_f (new_AGEMA_signal_6807), .Z0_t (SubBytesIns_Inst_Sbox_15_T13), .Z0_f (new_AGEMA_signal_7294), .Z1_t (new_AGEMA_signal_7295), .Z1_f (new_AGEMA_signal_7296) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T6), .A0_f (new_AGEMA_signal_7288), .A1_t (new_AGEMA_signal_7289), .A1_f (new_AGEMA_signal_7290), .B0_t (SubBytesIns_Inst_Sbox_15_T11), .B0_f (new_AGEMA_signal_6814), .B1_t (new_AGEMA_signal_6815), .B1_f (new_AGEMA_signal_6816), .Z0_t (SubBytesIns_Inst_Sbox_15_T14), .Z0_f (new_AGEMA_signal_8063), .Z1_t (new_AGEMA_signal_8064), .Z1_f (new_AGEMA_signal_8065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T5), .A0_f (new_AGEMA_signal_6808), .A1_t (new_AGEMA_signal_6809), .A1_f (new_AGEMA_signal_6810), .B0_t (SubBytesIns_Inst_Sbox_15_T11), .B0_f (new_AGEMA_signal_6814), .B1_t (new_AGEMA_signal_6815), .B1_f (new_AGEMA_signal_6816), .Z0_t (SubBytesIns_Inst_Sbox_15_T15), .Z0_f (new_AGEMA_signal_7297), .Z1_t (new_AGEMA_signal_7298), .Z1_f (new_AGEMA_signal_7299) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T5), .A0_f (new_AGEMA_signal_6808), .A1_t (new_AGEMA_signal_6809), .A1_f (new_AGEMA_signal_6810), .B0_t (SubBytesIns_Inst_Sbox_15_T12), .B0_f (new_AGEMA_signal_6817), .B1_t (new_AGEMA_signal_6818), .B1_f (new_AGEMA_signal_6819), .Z0_t (SubBytesIns_Inst_Sbox_15_T16), .Z0_f (new_AGEMA_signal_7300), .Z1_t (new_AGEMA_signal_7301), .Z1_f (new_AGEMA_signal_7302) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T9), .A0_f (new_AGEMA_signal_7291), .A1_t (new_AGEMA_signal_7292), .A1_f (new_AGEMA_signal_7293), .B0_t (SubBytesIns_Inst_Sbox_15_T16), .B0_f (new_AGEMA_signal_7300), .B1_t (new_AGEMA_signal_7301), .B1_f (new_AGEMA_signal_7302), .Z0_t (SubBytesIns_Inst_Sbox_15_T17), .Z0_f (new_AGEMA_signal_8066), .Z1_t (new_AGEMA_signal_8067), .Z1_f (new_AGEMA_signal_8068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T18_U1 ( .A0_t (ciphertext_s0_t[124]), .A0_f (ciphertext_s0_f[124]), .A1_t (ciphertext_s1_t[124]), .A1_f (ciphertext_s1_f[124]), .B0_t (ciphertext_s0_t[120]), .B0_f (ciphertext_s0_f[120]), .B1_t (ciphertext_s1_t[120]), .B1_f (ciphertext_s1_f[120]), .Z0_t (SubBytesIns_Inst_Sbox_15_T18), .Z0_f (new_AGEMA_signal_6820), .Z1_t (new_AGEMA_signal_6821), .Z1_f (new_AGEMA_signal_6822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T7), .A0_f (new_AGEMA_signal_6811), .A1_t (new_AGEMA_signal_6812), .A1_f (new_AGEMA_signal_6813), .B0_t (SubBytesIns_Inst_Sbox_15_T18), .B0_f (new_AGEMA_signal_6820), .B1_t (new_AGEMA_signal_6821), .B1_f (new_AGEMA_signal_6822), .Z0_t (SubBytesIns_Inst_Sbox_15_T19), .Z0_f (new_AGEMA_signal_7303), .Z1_t (new_AGEMA_signal_7304), .Z1_f (new_AGEMA_signal_7305) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T1), .A0_f (new_AGEMA_signal_6796), .A1_t (new_AGEMA_signal_6797), .A1_f (new_AGEMA_signal_6798), .B0_t (SubBytesIns_Inst_Sbox_15_T19), .B0_f (new_AGEMA_signal_7303), .B1_t (new_AGEMA_signal_7304), .B1_f (new_AGEMA_signal_7305), .Z0_t (SubBytesIns_Inst_Sbox_15_T20), .Z0_f (new_AGEMA_signal_8069), .Z1_t (new_AGEMA_signal_8070), .Z1_f (new_AGEMA_signal_8071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T21_U1 ( .A0_t (ciphertext_s0_t[121]), .A0_f (ciphertext_s0_f[121]), .A1_t (ciphertext_s1_t[121]), .A1_f (ciphertext_s1_f[121]), .B0_t (ciphertext_s0_t[120]), .B0_f (ciphertext_s0_f[120]), .B1_t (ciphertext_s1_t[120]), .B1_f (ciphertext_s1_f[120]), .Z0_t (SubBytesIns_Inst_Sbox_15_T21), .Z0_f (new_AGEMA_signal_6823), .Z1_t (new_AGEMA_signal_6824), .Z1_f (new_AGEMA_signal_6825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T7), .A0_f (new_AGEMA_signal_6811), .A1_t (new_AGEMA_signal_6812), .A1_f (new_AGEMA_signal_6813), .B0_t (SubBytesIns_Inst_Sbox_15_T21), .B0_f (new_AGEMA_signal_6823), .B1_t (new_AGEMA_signal_6824), .B1_f (new_AGEMA_signal_6825), .Z0_t (SubBytesIns_Inst_Sbox_15_T22), .Z0_f (new_AGEMA_signal_7306), .Z1_t (new_AGEMA_signal_7307), .Z1_f (new_AGEMA_signal_7308) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T2), .A0_f (new_AGEMA_signal_6799), .A1_t (new_AGEMA_signal_6800), .A1_f (new_AGEMA_signal_6801), .B0_t (SubBytesIns_Inst_Sbox_15_T22), .B0_f (new_AGEMA_signal_7306), .B1_t (new_AGEMA_signal_7307), .B1_f (new_AGEMA_signal_7308), .Z0_t (SubBytesIns_Inst_Sbox_15_T23), .Z0_f (new_AGEMA_signal_8072), .Z1_t (new_AGEMA_signal_8073), .Z1_f (new_AGEMA_signal_8074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T2), .A0_f (new_AGEMA_signal_6799), .A1_t (new_AGEMA_signal_6800), .A1_f (new_AGEMA_signal_6801), .B0_t (SubBytesIns_Inst_Sbox_15_T10), .B0_f (new_AGEMA_signal_8060), .B1_t (new_AGEMA_signal_8061), .B1_f (new_AGEMA_signal_8062), .Z0_t (SubBytesIns_Inst_Sbox_15_T24), .Z0_f (new_AGEMA_signal_8609), .Z1_t (new_AGEMA_signal_8610), .Z1_f (new_AGEMA_signal_8611) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T20), .A0_f (new_AGEMA_signal_8069), .A1_t (new_AGEMA_signal_8070), .A1_f (new_AGEMA_signal_8071), .B0_t (SubBytesIns_Inst_Sbox_15_T17), .B0_f (new_AGEMA_signal_8066), .B1_t (new_AGEMA_signal_8067), .B1_f (new_AGEMA_signal_8068), .Z0_t (SubBytesIns_Inst_Sbox_15_T25), .Z0_f (new_AGEMA_signal_8612), .Z1_t (new_AGEMA_signal_8613), .Z1_f (new_AGEMA_signal_8614) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T3), .A0_f (new_AGEMA_signal_6802), .A1_t (new_AGEMA_signal_6803), .A1_f (new_AGEMA_signal_6804), .B0_t (SubBytesIns_Inst_Sbox_15_T16), .B0_f (new_AGEMA_signal_7300), .B1_t (new_AGEMA_signal_7301), .B1_f (new_AGEMA_signal_7302), .Z0_t (SubBytesIns_Inst_Sbox_15_T26), .Z0_f (new_AGEMA_signal_8075), .Z1_t (new_AGEMA_signal_8076), .Z1_f (new_AGEMA_signal_8077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T1), .A0_f (new_AGEMA_signal_6796), .A1_t (new_AGEMA_signal_6797), .A1_f (new_AGEMA_signal_6798), .B0_t (SubBytesIns_Inst_Sbox_15_T12), .B0_f (new_AGEMA_signal_6817), .B1_t (new_AGEMA_signal_6818), .B1_f (new_AGEMA_signal_6819), .Z0_t (SubBytesIns_Inst_Sbox_15_T27), .Z0_f (new_AGEMA_signal_7309), .Z1_t (new_AGEMA_signal_7310), .Z1_f (new_AGEMA_signal_7311) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T13), .A0_f (new_AGEMA_signal_7294), .A1_t (new_AGEMA_signal_7295), .A1_f (new_AGEMA_signal_7296), .B0_t (SubBytesIns_Inst_Sbox_15_T6), .B0_f (new_AGEMA_signal_7288), .B1_t (new_AGEMA_signal_7289), .B1_f (new_AGEMA_signal_7290), .Z0_t (SubBytesIns_Inst_Sbox_15_M1), .Z0_f (new_AGEMA_signal_8078), .Z1_t (new_AGEMA_signal_8079), .Z1_f (new_AGEMA_signal_8080) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T23), .A0_f (new_AGEMA_signal_8072), .A1_t (new_AGEMA_signal_8073), .A1_f (new_AGEMA_signal_8074), .B0_t (SubBytesIns_Inst_Sbox_15_T8), .B0_f (new_AGEMA_signal_8057), .B1_t (new_AGEMA_signal_8058), .B1_f (new_AGEMA_signal_8059), .Z0_t (SubBytesIns_Inst_Sbox_15_M2), .Z0_f (new_AGEMA_signal_8615), .Z1_t (new_AGEMA_signal_8616), .Z1_f (new_AGEMA_signal_8617) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T14), .A0_f (new_AGEMA_signal_8063), .A1_t (new_AGEMA_signal_8064), .A1_f (new_AGEMA_signal_8065), .B0_t (SubBytesIns_Inst_Sbox_15_M1), .B0_f (new_AGEMA_signal_8078), .B1_t (new_AGEMA_signal_8079), .B1_f (new_AGEMA_signal_8080), .Z0_t (SubBytesIns_Inst_Sbox_15_M3), .Z0_f (new_AGEMA_signal_8618), .Z1_t (new_AGEMA_signal_8619), .Z1_f (new_AGEMA_signal_8620) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T19), .A0_f (new_AGEMA_signal_7303), .A1_t (new_AGEMA_signal_7304), .A1_f (new_AGEMA_signal_7305), .B0_t (ciphertext_s0_t[120]), .B0_f (ciphertext_s0_f[120]), .B1_t (ciphertext_s1_t[120]), .B1_f (ciphertext_s1_f[120]), .Z0_t (SubBytesIns_Inst_Sbox_15_M4), .Z0_f (new_AGEMA_signal_8081), .Z1_t (new_AGEMA_signal_8082), .Z1_f (new_AGEMA_signal_8083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M4), .A0_f (new_AGEMA_signal_8081), .A1_t (new_AGEMA_signal_8082), .A1_f (new_AGEMA_signal_8083), .B0_t (SubBytesIns_Inst_Sbox_15_M1), .B0_f (new_AGEMA_signal_8078), .B1_t (new_AGEMA_signal_8079), .B1_f (new_AGEMA_signal_8080), .Z0_t (SubBytesIns_Inst_Sbox_15_M5), .Z0_f (new_AGEMA_signal_8621), .Z1_t (new_AGEMA_signal_8622), .Z1_f (new_AGEMA_signal_8623) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T3), .A0_f (new_AGEMA_signal_6802), .A1_t (new_AGEMA_signal_6803), .A1_f (new_AGEMA_signal_6804), .B0_t (SubBytesIns_Inst_Sbox_15_T16), .B0_f (new_AGEMA_signal_7300), .B1_t (new_AGEMA_signal_7301), .B1_f (new_AGEMA_signal_7302), .Z0_t (SubBytesIns_Inst_Sbox_15_M6), .Z0_f (new_AGEMA_signal_8084), .Z1_t (new_AGEMA_signal_8085), .Z1_f (new_AGEMA_signal_8086) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T22), .A0_f (new_AGEMA_signal_7306), .A1_t (new_AGEMA_signal_7307), .A1_f (new_AGEMA_signal_7308), .B0_t (SubBytesIns_Inst_Sbox_15_T9), .B0_f (new_AGEMA_signal_7291), .B1_t (new_AGEMA_signal_7292), .B1_f (new_AGEMA_signal_7293), .Z0_t (SubBytesIns_Inst_Sbox_15_M7), .Z0_f (new_AGEMA_signal_8087), .Z1_t (new_AGEMA_signal_8088), .Z1_f (new_AGEMA_signal_8089) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T26), .A0_f (new_AGEMA_signal_8075), .A1_t (new_AGEMA_signal_8076), .A1_f (new_AGEMA_signal_8077), .B0_t (SubBytesIns_Inst_Sbox_15_M6), .B0_f (new_AGEMA_signal_8084), .B1_t (new_AGEMA_signal_8085), .B1_f (new_AGEMA_signal_8086), .Z0_t (SubBytesIns_Inst_Sbox_15_M8), .Z0_f (new_AGEMA_signal_8624), .Z1_t (new_AGEMA_signal_8625), .Z1_f (new_AGEMA_signal_8626) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T20), .A0_f (new_AGEMA_signal_8069), .A1_t (new_AGEMA_signal_8070), .A1_f (new_AGEMA_signal_8071), .B0_t (SubBytesIns_Inst_Sbox_15_T17), .B0_f (new_AGEMA_signal_8066), .B1_t (new_AGEMA_signal_8067), .B1_f (new_AGEMA_signal_8068), .Z0_t (SubBytesIns_Inst_Sbox_15_M9), .Z0_f (new_AGEMA_signal_8627), .Z1_t (new_AGEMA_signal_8628), .Z1_f (new_AGEMA_signal_8629) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M9), .A0_f (new_AGEMA_signal_8627), .A1_t (new_AGEMA_signal_8628), .A1_f (new_AGEMA_signal_8629), .B0_t (SubBytesIns_Inst_Sbox_15_M6), .B0_f (new_AGEMA_signal_8084), .B1_t (new_AGEMA_signal_8085), .B1_f (new_AGEMA_signal_8086), .Z0_t (SubBytesIns_Inst_Sbox_15_M10), .Z0_f (new_AGEMA_signal_8921), .Z1_t (new_AGEMA_signal_8922), .Z1_f (new_AGEMA_signal_8923) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T1), .A0_f (new_AGEMA_signal_6796), .A1_t (new_AGEMA_signal_6797), .A1_f (new_AGEMA_signal_6798), .B0_t (SubBytesIns_Inst_Sbox_15_T15), .B0_f (new_AGEMA_signal_7297), .B1_t (new_AGEMA_signal_7298), .B1_f (new_AGEMA_signal_7299), .Z0_t (SubBytesIns_Inst_Sbox_15_M11), .Z0_f (new_AGEMA_signal_8090), .Z1_t (new_AGEMA_signal_8091), .Z1_f (new_AGEMA_signal_8092) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T4), .A0_f (new_AGEMA_signal_6805), .A1_t (new_AGEMA_signal_6806), .A1_f (new_AGEMA_signal_6807), .B0_t (SubBytesIns_Inst_Sbox_15_T27), .B0_f (new_AGEMA_signal_7309), .B1_t (new_AGEMA_signal_7310), .B1_f (new_AGEMA_signal_7311), .Z0_t (SubBytesIns_Inst_Sbox_15_M12), .Z0_f (new_AGEMA_signal_8093), .Z1_t (new_AGEMA_signal_8094), .Z1_f (new_AGEMA_signal_8095) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M12), .A0_f (new_AGEMA_signal_8093), .A1_t (new_AGEMA_signal_8094), .A1_f (new_AGEMA_signal_8095), .B0_t (SubBytesIns_Inst_Sbox_15_M11), .B0_f (new_AGEMA_signal_8090), .B1_t (new_AGEMA_signal_8091), .B1_f (new_AGEMA_signal_8092), .Z0_t (SubBytesIns_Inst_Sbox_15_M13), .Z0_f (new_AGEMA_signal_8630), .Z1_t (new_AGEMA_signal_8631), .Z1_f (new_AGEMA_signal_8632) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T2), .A0_f (new_AGEMA_signal_6799), .A1_t (new_AGEMA_signal_6800), .A1_f (new_AGEMA_signal_6801), .B0_t (SubBytesIns_Inst_Sbox_15_T10), .B0_f (new_AGEMA_signal_8060), .B1_t (new_AGEMA_signal_8061), .B1_f (new_AGEMA_signal_8062), .Z0_t (SubBytesIns_Inst_Sbox_15_M14), .Z0_f (new_AGEMA_signal_8633), .Z1_t (new_AGEMA_signal_8634), .Z1_f (new_AGEMA_signal_8635) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M14), .A0_f (new_AGEMA_signal_8633), .A1_t (new_AGEMA_signal_8634), .A1_f (new_AGEMA_signal_8635), .B0_t (SubBytesIns_Inst_Sbox_15_M11), .B0_f (new_AGEMA_signal_8090), .B1_t (new_AGEMA_signal_8091), .B1_f (new_AGEMA_signal_8092), .Z0_t (SubBytesIns_Inst_Sbox_15_M15), .Z0_f (new_AGEMA_signal_8924), .Z1_t (new_AGEMA_signal_8925), .Z1_f (new_AGEMA_signal_8926) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M3), .A0_f (new_AGEMA_signal_8618), .A1_t (new_AGEMA_signal_8619), .A1_f (new_AGEMA_signal_8620), .B0_t (SubBytesIns_Inst_Sbox_15_M2), .B0_f (new_AGEMA_signal_8615), .B1_t (new_AGEMA_signal_8616), .B1_f (new_AGEMA_signal_8617), .Z0_t (SubBytesIns_Inst_Sbox_15_M16), .Z0_f (new_AGEMA_signal_8927), .Z1_t (new_AGEMA_signal_8928), .Z1_f (new_AGEMA_signal_8929) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M5), .A0_f (new_AGEMA_signal_8621), .A1_t (new_AGEMA_signal_8622), .A1_f (new_AGEMA_signal_8623), .B0_t (SubBytesIns_Inst_Sbox_15_T24), .B0_f (new_AGEMA_signal_8609), .B1_t (new_AGEMA_signal_8610), .B1_f (new_AGEMA_signal_8611), .Z0_t (SubBytesIns_Inst_Sbox_15_M17), .Z0_f (new_AGEMA_signal_8930), .Z1_t (new_AGEMA_signal_8931), .Z1_f (new_AGEMA_signal_8932) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M8), .A0_f (new_AGEMA_signal_8624), .A1_t (new_AGEMA_signal_8625), .A1_f (new_AGEMA_signal_8626), .B0_t (SubBytesIns_Inst_Sbox_15_M7), .B0_f (new_AGEMA_signal_8087), .B1_t (new_AGEMA_signal_8088), .B1_f (new_AGEMA_signal_8089), .Z0_t (SubBytesIns_Inst_Sbox_15_M18), .Z0_f (new_AGEMA_signal_8933), .Z1_t (new_AGEMA_signal_8934), .Z1_f (new_AGEMA_signal_8935) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M10), .A0_f (new_AGEMA_signal_8921), .A1_t (new_AGEMA_signal_8922), .A1_f (new_AGEMA_signal_8923), .B0_t (SubBytesIns_Inst_Sbox_15_M15), .B0_f (new_AGEMA_signal_8924), .B1_t (new_AGEMA_signal_8925), .B1_f (new_AGEMA_signal_8926), .Z0_t (SubBytesIns_Inst_Sbox_15_M19), .Z0_f (new_AGEMA_signal_9164), .Z1_t (new_AGEMA_signal_9165), .Z1_f (new_AGEMA_signal_9166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M16), .A0_f (new_AGEMA_signal_8927), .A1_t (new_AGEMA_signal_8928), .A1_f (new_AGEMA_signal_8929), .B0_t (SubBytesIns_Inst_Sbox_15_M13), .B0_f (new_AGEMA_signal_8630), .B1_t (new_AGEMA_signal_8631), .B1_f (new_AGEMA_signal_8632), .Z0_t (SubBytesIns_Inst_Sbox_15_M20), .Z0_f (new_AGEMA_signal_9167), .Z1_t (new_AGEMA_signal_9168), .Z1_f (new_AGEMA_signal_9169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M17), .A0_f (new_AGEMA_signal_8930), .A1_t (new_AGEMA_signal_8931), .A1_f (new_AGEMA_signal_8932), .B0_t (SubBytesIns_Inst_Sbox_15_M15), .B0_f (new_AGEMA_signal_8924), .B1_t (new_AGEMA_signal_8925), .B1_f (new_AGEMA_signal_8926), .Z0_t (SubBytesIns_Inst_Sbox_15_M21), .Z0_f (new_AGEMA_signal_9170), .Z1_t (new_AGEMA_signal_9171), .Z1_f (new_AGEMA_signal_9172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M18), .A0_f (new_AGEMA_signal_8933), .A1_t (new_AGEMA_signal_8934), .A1_f (new_AGEMA_signal_8935), .B0_t (SubBytesIns_Inst_Sbox_15_M13), .B0_f (new_AGEMA_signal_8630), .B1_t (new_AGEMA_signal_8631), .B1_f (new_AGEMA_signal_8632), .Z0_t (SubBytesIns_Inst_Sbox_15_M22), .Z0_f (new_AGEMA_signal_9173), .Z1_t (new_AGEMA_signal_9174), .Z1_f (new_AGEMA_signal_9175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M19), .A0_f (new_AGEMA_signal_9164), .A1_t (new_AGEMA_signal_9165), .A1_f (new_AGEMA_signal_9166), .B0_t (SubBytesIns_Inst_Sbox_15_T25), .B0_f (new_AGEMA_signal_8612), .B1_t (new_AGEMA_signal_8613), .B1_f (new_AGEMA_signal_8614), .Z0_t (SubBytesIns_Inst_Sbox_15_M23), .Z0_f (new_AGEMA_signal_9404), .Z1_t (new_AGEMA_signal_9405), .Z1_f (new_AGEMA_signal_9406) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M22), .A0_f (new_AGEMA_signal_9173), .A1_t (new_AGEMA_signal_9174), .A1_f (new_AGEMA_signal_9175), .B0_t (SubBytesIns_Inst_Sbox_15_M23), .B0_f (new_AGEMA_signal_9404), .B1_t (new_AGEMA_signal_9405), .B1_f (new_AGEMA_signal_9406), .Z0_t (SubBytesIns_Inst_Sbox_15_M24), .Z0_f (new_AGEMA_signal_9701), .Z1_t (new_AGEMA_signal_9702), .Z1_f (new_AGEMA_signal_9703) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M22), .A0_f (new_AGEMA_signal_9173), .A1_t (new_AGEMA_signal_9174), .A1_f (new_AGEMA_signal_9175), .B0_t (SubBytesIns_Inst_Sbox_15_M20), .B0_f (new_AGEMA_signal_9167), .B1_t (new_AGEMA_signal_9168), .B1_f (new_AGEMA_signal_9169), .Z0_t (SubBytesIns_Inst_Sbox_15_M25), .Z0_f (new_AGEMA_signal_9407), .Z1_t (new_AGEMA_signal_9408), .Z1_f (new_AGEMA_signal_9409) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M21), .A0_f (new_AGEMA_signal_9170), .A1_t (new_AGEMA_signal_9171), .A1_f (new_AGEMA_signal_9172), .B0_t (SubBytesIns_Inst_Sbox_15_M25), .B0_f (new_AGEMA_signal_9407), .B1_t (new_AGEMA_signal_9408), .B1_f (new_AGEMA_signal_9409), .Z0_t (SubBytesIns_Inst_Sbox_15_M26), .Z0_f (new_AGEMA_signal_9704), .Z1_t (new_AGEMA_signal_9705), .Z1_f (new_AGEMA_signal_9706) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M20), .A0_f (new_AGEMA_signal_9167), .A1_t (new_AGEMA_signal_9168), .A1_f (new_AGEMA_signal_9169), .B0_t (SubBytesIns_Inst_Sbox_15_M21), .B0_f (new_AGEMA_signal_9170), .B1_t (new_AGEMA_signal_9171), .B1_f (new_AGEMA_signal_9172), .Z0_t (SubBytesIns_Inst_Sbox_15_M27), .Z0_f (new_AGEMA_signal_9410), .Z1_t (new_AGEMA_signal_9411), .Z1_f (new_AGEMA_signal_9412) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M23), .A0_f (new_AGEMA_signal_9404), .A1_t (new_AGEMA_signal_9405), .A1_f (new_AGEMA_signal_9406), .B0_t (SubBytesIns_Inst_Sbox_15_M25), .B0_f (new_AGEMA_signal_9407), .B1_t (new_AGEMA_signal_9408), .B1_f (new_AGEMA_signal_9409), .Z0_t (SubBytesIns_Inst_Sbox_15_M28), .Z0_f (new_AGEMA_signal_9707), .Z1_t (new_AGEMA_signal_9708), .Z1_f (new_AGEMA_signal_9709) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M28), .A0_f (new_AGEMA_signal_9707), .A1_t (new_AGEMA_signal_9708), .A1_f (new_AGEMA_signal_9709), .B0_t (SubBytesIns_Inst_Sbox_15_M27), .B0_f (new_AGEMA_signal_9410), .B1_t (new_AGEMA_signal_9411), .B1_f (new_AGEMA_signal_9412), .Z0_t (SubBytesIns_Inst_Sbox_15_M29), .Z0_f (new_AGEMA_signal_10001), .Z1_t (new_AGEMA_signal_10002), .Z1_f (new_AGEMA_signal_10003) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M26), .A0_f (new_AGEMA_signal_9704), .A1_t (new_AGEMA_signal_9705), .A1_f (new_AGEMA_signal_9706), .B0_t (SubBytesIns_Inst_Sbox_15_M24), .B0_f (new_AGEMA_signal_9701), .B1_t (new_AGEMA_signal_9702), .B1_f (new_AGEMA_signal_9703), .Z0_t (SubBytesIns_Inst_Sbox_15_M30), .Z0_f (new_AGEMA_signal_10004), .Z1_t (new_AGEMA_signal_10005), .Z1_f (new_AGEMA_signal_10006) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M20), .A0_f (new_AGEMA_signal_9167), .A1_t (new_AGEMA_signal_9168), .A1_f (new_AGEMA_signal_9169), .B0_t (SubBytesIns_Inst_Sbox_15_M23), .B0_f (new_AGEMA_signal_9404), .B1_t (new_AGEMA_signal_9405), .B1_f (new_AGEMA_signal_9406), .Z0_t (SubBytesIns_Inst_Sbox_15_M31), .Z0_f (new_AGEMA_signal_9710), .Z1_t (new_AGEMA_signal_9711), .Z1_f (new_AGEMA_signal_9712) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M27), .A0_f (new_AGEMA_signal_9410), .A1_t (new_AGEMA_signal_9411), .A1_f (new_AGEMA_signal_9412), .B0_t (SubBytesIns_Inst_Sbox_15_M31), .B0_f (new_AGEMA_signal_9710), .B1_t (new_AGEMA_signal_9711), .B1_f (new_AGEMA_signal_9712), .Z0_t (SubBytesIns_Inst_Sbox_15_M32), .Z0_f (new_AGEMA_signal_10007), .Z1_t (new_AGEMA_signal_10008), .Z1_f (new_AGEMA_signal_10009) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M27), .A0_f (new_AGEMA_signal_9410), .A1_t (new_AGEMA_signal_9411), .A1_f (new_AGEMA_signal_9412), .B0_t (SubBytesIns_Inst_Sbox_15_M25), .B0_f (new_AGEMA_signal_9407), .B1_t (new_AGEMA_signal_9408), .B1_f (new_AGEMA_signal_9409), .Z0_t (SubBytesIns_Inst_Sbox_15_M33), .Z0_f (new_AGEMA_signal_9713), .Z1_t (new_AGEMA_signal_9714), .Z1_f (new_AGEMA_signal_9715) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M21), .A0_f (new_AGEMA_signal_9170), .A1_t (new_AGEMA_signal_9171), .A1_f (new_AGEMA_signal_9172), .B0_t (SubBytesIns_Inst_Sbox_15_M22), .B0_f (new_AGEMA_signal_9173), .B1_t (new_AGEMA_signal_9174), .B1_f (new_AGEMA_signal_9175), .Z0_t (SubBytesIns_Inst_Sbox_15_M34), .Z0_f (new_AGEMA_signal_9413), .Z1_t (new_AGEMA_signal_9414), .Z1_f (new_AGEMA_signal_9415) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M24), .A0_f (new_AGEMA_signal_9701), .A1_t (new_AGEMA_signal_9702), .A1_f (new_AGEMA_signal_9703), .B0_t (SubBytesIns_Inst_Sbox_15_M34), .B0_f (new_AGEMA_signal_9413), .B1_t (new_AGEMA_signal_9414), .B1_f (new_AGEMA_signal_9415), .Z0_t (SubBytesIns_Inst_Sbox_15_M35), .Z0_f (new_AGEMA_signal_10010), .Z1_t (new_AGEMA_signal_10011), .Z1_f (new_AGEMA_signal_10012) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M24), .A0_f (new_AGEMA_signal_9701), .A1_t (new_AGEMA_signal_9702), .A1_f (new_AGEMA_signal_9703), .B0_t (SubBytesIns_Inst_Sbox_15_M25), .B0_f (new_AGEMA_signal_9407), .B1_t (new_AGEMA_signal_9408), .B1_f (new_AGEMA_signal_9409), .Z0_t (SubBytesIns_Inst_Sbox_15_M36), .Z0_f (new_AGEMA_signal_10013), .Z1_t (new_AGEMA_signal_10014), .Z1_f (new_AGEMA_signal_10015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M21), .A0_f (new_AGEMA_signal_9170), .A1_t (new_AGEMA_signal_9171), .A1_f (new_AGEMA_signal_9172), .B0_t (SubBytesIns_Inst_Sbox_15_M29), .B0_f (new_AGEMA_signal_10001), .B1_t (new_AGEMA_signal_10002), .B1_f (new_AGEMA_signal_10003), .Z0_t (SubBytesIns_Inst_Sbox_15_M37), .Z0_f (new_AGEMA_signal_10244), .Z1_t (new_AGEMA_signal_10245), .Z1_f (new_AGEMA_signal_10246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M32), .A0_f (new_AGEMA_signal_10007), .A1_t (new_AGEMA_signal_10008), .A1_f (new_AGEMA_signal_10009), .B0_t (SubBytesIns_Inst_Sbox_15_M33), .B0_f (new_AGEMA_signal_9713), .B1_t (new_AGEMA_signal_9714), .B1_f (new_AGEMA_signal_9715), .Z0_t (SubBytesIns_Inst_Sbox_15_M38), .Z0_f (new_AGEMA_signal_10247), .Z1_t (new_AGEMA_signal_10248), .Z1_f (new_AGEMA_signal_10249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M23), .A0_f (new_AGEMA_signal_9404), .A1_t (new_AGEMA_signal_9405), .A1_f (new_AGEMA_signal_9406), .B0_t (SubBytesIns_Inst_Sbox_15_M30), .B0_f (new_AGEMA_signal_10004), .B1_t (new_AGEMA_signal_10005), .B1_f (new_AGEMA_signal_10006), .Z0_t (SubBytesIns_Inst_Sbox_15_M39), .Z0_f (new_AGEMA_signal_10250), .Z1_t (new_AGEMA_signal_10251), .Z1_f (new_AGEMA_signal_10252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M35), .A0_f (new_AGEMA_signal_10010), .A1_t (new_AGEMA_signal_10011), .A1_f (new_AGEMA_signal_10012), .B0_t (SubBytesIns_Inst_Sbox_15_M36), .B0_f (new_AGEMA_signal_10013), .B1_t (new_AGEMA_signal_10014), .B1_f (new_AGEMA_signal_10015), .Z0_t (SubBytesIns_Inst_Sbox_15_M40), .Z0_f (new_AGEMA_signal_10253), .Z1_t (new_AGEMA_signal_10254), .Z1_f (new_AGEMA_signal_10255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M38), .A0_f (new_AGEMA_signal_10247), .A1_t (new_AGEMA_signal_10248), .A1_f (new_AGEMA_signal_10249), .B0_t (SubBytesIns_Inst_Sbox_15_M40), .B0_f (new_AGEMA_signal_10253), .B1_t (new_AGEMA_signal_10254), .B1_f (new_AGEMA_signal_10255), .Z0_t (SubBytesIns_Inst_Sbox_15_M41), .Z0_f (new_AGEMA_signal_10940), .Z1_t (new_AGEMA_signal_10941), .Z1_f (new_AGEMA_signal_10942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M37), .A0_f (new_AGEMA_signal_10244), .A1_t (new_AGEMA_signal_10245), .A1_f (new_AGEMA_signal_10246), .B0_t (SubBytesIns_Inst_Sbox_15_M39), .B0_f (new_AGEMA_signal_10250), .B1_t (new_AGEMA_signal_10251), .B1_f (new_AGEMA_signal_10252), .Z0_t (SubBytesIns_Inst_Sbox_15_M42), .Z0_f (new_AGEMA_signal_10943), .Z1_t (new_AGEMA_signal_10944), .Z1_f (new_AGEMA_signal_10945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M37), .A0_f (new_AGEMA_signal_10244), .A1_t (new_AGEMA_signal_10245), .A1_f (new_AGEMA_signal_10246), .B0_t (SubBytesIns_Inst_Sbox_15_M38), .B0_f (new_AGEMA_signal_10247), .B1_t (new_AGEMA_signal_10248), .B1_f (new_AGEMA_signal_10249), .Z0_t (SubBytesIns_Inst_Sbox_15_M43), .Z0_f (new_AGEMA_signal_10946), .Z1_t (new_AGEMA_signal_10947), .Z1_f (new_AGEMA_signal_10948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M39), .A0_f (new_AGEMA_signal_10250), .A1_t (new_AGEMA_signal_10251), .A1_f (new_AGEMA_signal_10252), .B0_t (SubBytesIns_Inst_Sbox_15_M40), .B0_f (new_AGEMA_signal_10253), .B1_t (new_AGEMA_signal_10254), .B1_f (new_AGEMA_signal_10255), .Z0_t (SubBytesIns_Inst_Sbox_15_M44), .Z0_f (new_AGEMA_signal_10949), .Z1_t (new_AGEMA_signal_10950), .Z1_f (new_AGEMA_signal_10951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M42), .A0_f (new_AGEMA_signal_10943), .A1_t (new_AGEMA_signal_10944), .A1_f (new_AGEMA_signal_10945), .B0_t (SubBytesIns_Inst_Sbox_15_M41), .B0_f (new_AGEMA_signal_10940), .B1_t (new_AGEMA_signal_10941), .B1_f (new_AGEMA_signal_10942), .Z0_t (SubBytesIns_Inst_Sbox_15_M45), .Z0_f (new_AGEMA_signal_11660), .Z1_t (new_AGEMA_signal_11661), .Z1_f (new_AGEMA_signal_11662) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M44), .A0_f (new_AGEMA_signal_10949), .A1_t (new_AGEMA_signal_10950), .A1_f (new_AGEMA_signal_10951), .B0_t (SubBytesIns_Inst_Sbox_15_T6), .B0_f (new_AGEMA_signal_7288), .B1_t (new_AGEMA_signal_7289), .B1_f (new_AGEMA_signal_7290), .Z0_t (SubBytesIns_Inst_Sbox_15_M46), .Z0_f (new_AGEMA_signal_11663), .Z1_t (new_AGEMA_signal_11664), .Z1_f (new_AGEMA_signal_11665) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M40), .A0_f (new_AGEMA_signal_10253), .A1_t (new_AGEMA_signal_10254), .A1_f (new_AGEMA_signal_10255), .B0_t (SubBytesIns_Inst_Sbox_15_T8), .B0_f (new_AGEMA_signal_8057), .B1_t (new_AGEMA_signal_8058), .B1_f (new_AGEMA_signal_8059), .Z0_t (SubBytesIns_Inst_Sbox_15_M47), .Z0_f (new_AGEMA_signal_10952), .Z1_t (new_AGEMA_signal_10953), .Z1_f (new_AGEMA_signal_10954) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M39), .A0_f (new_AGEMA_signal_10250), .A1_t (new_AGEMA_signal_10251), .A1_f (new_AGEMA_signal_10252), .B0_t (ciphertext_s0_t[120]), .B0_f (ciphertext_s0_f[120]), .B1_t (ciphertext_s1_t[120]), .B1_f (ciphertext_s1_f[120]), .Z0_t (SubBytesIns_Inst_Sbox_15_M48), .Z0_f (new_AGEMA_signal_10955), .Z1_t (new_AGEMA_signal_10956), .Z1_f (new_AGEMA_signal_10957) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M43), .A0_f (new_AGEMA_signal_10946), .A1_t (new_AGEMA_signal_10947), .A1_f (new_AGEMA_signal_10948), .B0_t (SubBytesIns_Inst_Sbox_15_T16), .B0_f (new_AGEMA_signal_7300), .B1_t (new_AGEMA_signal_7301), .B1_f (new_AGEMA_signal_7302), .Z0_t (SubBytesIns_Inst_Sbox_15_M49), .Z0_f (new_AGEMA_signal_11666), .Z1_t (new_AGEMA_signal_11667), .Z1_f (new_AGEMA_signal_11668) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M38), .A0_f (new_AGEMA_signal_10247), .A1_t (new_AGEMA_signal_10248), .A1_f (new_AGEMA_signal_10249), .B0_t (SubBytesIns_Inst_Sbox_15_T9), .B0_f (new_AGEMA_signal_7291), .B1_t (new_AGEMA_signal_7292), .B1_f (new_AGEMA_signal_7293), .Z0_t (SubBytesIns_Inst_Sbox_15_M50), .Z0_f (new_AGEMA_signal_10958), .Z1_t (new_AGEMA_signal_10959), .Z1_f (new_AGEMA_signal_10960) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M37), .A0_f (new_AGEMA_signal_10244), .A1_t (new_AGEMA_signal_10245), .A1_f (new_AGEMA_signal_10246), .B0_t (SubBytesIns_Inst_Sbox_15_T17), .B0_f (new_AGEMA_signal_8066), .B1_t (new_AGEMA_signal_8067), .B1_f (new_AGEMA_signal_8068), .Z0_t (SubBytesIns_Inst_Sbox_15_M51), .Z0_f (new_AGEMA_signal_10961), .Z1_t (new_AGEMA_signal_10962), .Z1_f (new_AGEMA_signal_10963) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M42), .A0_f (new_AGEMA_signal_10943), .A1_t (new_AGEMA_signal_10944), .A1_f (new_AGEMA_signal_10945), .B0_t (SubBytesIns_Inst_Sbox_15_T15), .B0_f (new_AGEMA_signal_7297), .B1_t (new_AGEMA_signal_7298), .B1_f (new_AGEMA_signal_7299), .Z0_t (SubBytesIns_Inst_Sbox_15_M52), .Z0_f (new_AGEMA_signal_11669), .Z1_t (new_AGEMA_signal_11670), .Z1_f (new_AGEMA_signal_11671) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M45), .A0_f (new_AGEMA_signal_11660), .A1_t (new_AGEMA_signal_11661), .A1_f (new_AGEMA_signal_11662), .B0_t (SubBytesIns_Inst_Sbox_15_T27), .B0_f (new_AGEMA_signal_7309), .B1_t (new_AGEMA_signal_7310), .B1_f (new_AGEMA_signal_7311), .Z0_t (SubBytesIns_Inst_Sbox_15_M53), .Z0_f (new_AGEMA_signal_12266), .Z1_t (new_AGEMA_signal_12267), .Z1_f (new_AGEMA_signal_12268) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M41), .A0_f (new_AGEMA_signal_10940), .A1_t (new_AGEMA_signal_10941), .A1_f (new_AGEMA_signal_10942), .B0_t (SubBytesIns_Inst_Sbox_15_T10), .B0_f (new_AGEMA_signal_8060), .B1_t (new_AGEMA_signal_8061), .B1_f (new_AGEMA_signal_8062), .Z0_t (SubBytesIns_Inst_Sbox_15_M54), .Z0_f (new_AGEMA_signal_11672), .Z1_t (new_AGEMA_signal_11673), .Z1_f (new_AGEMA_signal_11674) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M44), .A0_f (new_AGEMA_signal_10949), .A1_t (new_AGEMA_signal_10950), .A1_f (new_AGEMA_signal_10951), .B0_t (SubBytesIns_Inst_Sbox_15_T13), .B0_f (new_AGEMA_signal_7294), .B1_t (new_AGEMA_signal_7295), .B1_f (new_AGEMA_signal_7296), .Z0_t (SubBytesIns_Inst_Sbox_15_M55), .Z0_f (new_AGEMA_signal_11675), .Z1_t (new_AGEMA_signal_11676), .Z1_f (new_AGEMA_signal_11677) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M40), .A0_f (new_AGEMA_signal_10253), .A1_t (new_AGEMA_signal_10254), .A1_f (new_AGEMA_signal_10255), .B0_t (SubBytesIns_Inst_Sbox_15_T23), .B0_f (new_AGEMA_signal_8072), .B1_t (new_AGEMA_signal_8073), .B1_f (new_AGEMA_signal_8074), .Z0_t (SubBytesIns_Inst_Sbox_15_M56), .Z0_f (new_AGEMA_signal_10964), .Z1_t (new_AGEMA_signal_10965), .Z1_f (new_AGEMA_signal_10966) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M39), .A0_f (new_AGEMA_signal_10250), .A1_t (new_AGEMA_signal_10251), .A1_f (new_AGEMA_signal_10252), .B0_t (SubBytesIns_Inst_Sbox_15_T19), .B0_f (new_AGEMA_signal_7303), .B1_t (new_AGEMA_signal_7304), .B1_f (new_AGEMA_signal_7305), .Z0_t (SubBytesIns_Inst_Sbox_15_M57), .Z0_f (new_AGEMA_signal_10967), .Z1_t (new_AGEMA_signal_10968), .Z1_f (new_AGEMA_signal_10969) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M43), .A0_f (new_AGEMA_signal_10946), .A1_t (new_AGEMA_signal_10947), .A1_f (new_AGEMA_signal_10948), .B0_t (SubBytesIns_Inst_Sbox_15_T3), .B0_f (new_AGEMA_signal_6802), .B1_t (new_AGEMA_signal_6803), .B1_f (new_AGEMA_signal_6804), .Z0_t (SubBytesIns_Inst_Sbox_15_M58), .Z0_f (new_AGEMA_signal_11678), .Z1_t (new_AGEMA_signal_11679), .Z1_f (new_AGEMA_signal_11680) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M38), .A0_f (new_AGEMA_signal_10247), .A1_t (new_AGEMA_signal_10248), .A1_f (new_AGEMA_signal_10249), .B0_t (SubBytesIns_Inst_Sbox_15_T22), .B0_f (new_AGEMA_signal_7306), .B1_t (new_AGEMA_signal_7307), .B1_f (new_AGEMA_signal_7308), .Z0_t (SubBytesIns_Inst_Sbox_15_M59), .Z0_f (new_AGEMA_signal_10970), .Z1_t (new_AGEMA_signal_10971), .Z1_f (new_AGEMA_signal_10972) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M37), .A0_f (new_AGEMA_signal_10244), .A1_t (new_AGEMA_signal_10245), .A1_f (new_AGEMA_signal_10246), .B0_t (SubBytesIns_Inst_Sbox_15_T20), .B0_f (new_AGEMA_signal_8069), .B1_t (new_AGEMA_signal_8070), .B1_f (new_AGEMA_signal_8071), .Z0_t (SubBytesIns_Inst_Sbox_15_M60), .Z0_f (new_AGEMA_signal_10973), .Z1_t (new_AGEMA_signal_10974), .Z1_f (new_AGEMA_signal_10975) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M42), .A0_f (new_AGEMA_signal_10943), .A1_t (new_AGEMA_signal_10944), .A1_f (new_AGEMA_signal_10945), .B0_t (SubBytesIns_Inst_Sbox_15_T1), .B0_f (new_AGEMA_signal_6796), .B1_t (new_AGEMA_signal_6797), .B1_f (new_AGEMA_signal_6798), .Z0_t (SubBytesIns_Inst_Sbox_15_M61), .Z0_f (new_AGEMA_signal_11681), .Z1_t (new_AGEMA_signal_11682), .Z1_f (new_AGEMA_signal_11683) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M45), .A0_f (new_AGEMA_signal_11660), .A1_t (new_AGEMA_signal_11661), .A1_f (new_AGEMA_signal_11662), .B0_t (SubBytesIns_Inst_Sbox_15_T4), .B0_f (new_AGEMA_signal_6805), .B1_t (new_AGEMA_signal_6806), .B1_f (new_AGEMA_signal_6807), .Z0_t (SubBytesIns_Inst_Sbox_15_M62), .Z0_f (new_AGEMA_signal_12269), .Z1_t (new_AGEMA_signal_12270), .Z1_f (new_AGEMA_signal_12271) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M41), .A0_f (new_AGEMA_signal_10940), .A1_t (new_AGEMA_signal_10941), .A1_f (new_AGEMA_signal_10942), .B0_t (SubBytesIns_Inst_Sbox_15_T2), .B0_f (new_AGEMA_signal_6799), .B1_t (new_AGEMA_signal_6800), .B1_f (new_AGEMA_signal_6801), .Z0_t (SubBytesIns_Inst_Sbox_15_M63), .Z0_f (new_AGEMA_signal_11684), .Z1_t (new_AGEMA_signal_11685), .Z1_f (new_AGEMA_signal_11686) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M61), .A0_f (new_AGEMA_signal_11681), .A1_t (new_AGEMA_signal_11682), .A1_f (new_AGEMA_signal_11683), .B0_t (SubBytesIns_Inst_Sbox_15_M62), .B0_f (new_AGEMA_signal_12269), .B1_t (new_AGEMA_signal_12270), .B1_f (new_AGEMA_signal_12271), .Z0_t (SubBytesIns_Inst_Sbox_15_L0), .Z0_f (new_AGEMA_signal_12809), .Z1_t (new_AGEMA_signal_12810), .Z1_f (new_AGEMA_signal_12811) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M50), .A0_f (new_AGEMA_signal_10958), .A1_t (new_AGEMA_signal_10959), .A1_f (new_AGEMA_signal_10960), .B0_t (SubBytesIns_Inst_Sbox_15_M56), .B0_f (new_AGEMA_signal_10964), .B1_t (new_AGEMA_signal_10965), .B1_f (new_AGEMA_signal_10966), .Z0_t (SubBytesIns_Inst_Sbox_15_L1), .Z0_f (new_AGEMA_signal_11687), .Z1_t (new_AGEMA_signal_11688), .Z1_f (new_AGEMA_signal_11689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M46), .A0_f (new_AGEMA_signal_11663), .A1_t (new_AGEMA_signal_11664), .A1_f (new_AGEMA_signal_11665), .B0_t (SubBytesIns_Inst_Sbox_15_M48), .B0_f (new_AGEMA_signal_10955), .B1_t (new_AGEMA_signal_10956), .B1_f (new_AGEMA_signal_10957), .Z0_t (SubBytesIns_Inst_Sbox_15_L2), .Z0_f (new_AGEMA_signal_12272), .Z1_t (new_AGEMA_signal_12273), .Z1_f (new_AGEMA_signal_12274) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M47), .A0_f (new_AGEMA_signal_10952), .A1_t (new_AGEMA_signal_10953), .A1_f (new_AGEMA_signal_10954), .B0_t (SubBytesIns_Inst_Sbox_15_M55), .B0_f (new_AGEMA_signal_11675), .B1_t (new_AGEMA_signal_11676), .B1_f (new_AGEMA_signal_11677), .Z0_t (SubBytesIns_Inst_Sbox_15_L3), .Z0_f (new_AGEMA_signal_12275), .Z1_t (new_AGEMA_signal_12276), .Z1_f (new_AGEMA_signal_12277) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M54), .A0_f (new_AGEMA_signal_11672), .A1_t (new_AGEMA_signal_11673), .A1_f (new_AGEMA_signal_11674), .B0_t (SubBytesIns_Inst_Sbox_15_M58), .B0_f (new_AGEMA_signal_11678), .B1_t (new_AGEMA_signal_11679), .B1_f (new_AGEMA_signal_11680), .Z0_t (SubBytesIns_Inst_Sbox_15_L4), .Z0_f (new_AGEMA_signal_12278), .Z1_t (new_AGEMA_signal_12279), .Z1_f (new_AGEMA_signal_12280) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M49), .A0_f (new_AGEMA_signal_11666), .A1_t (new_AGEMA_signal_11667), .A1_f (new_AGEMA_signal_11668), .B0_t (SubBytesIns_Inst_Sbox_15_M61), .B0_f (new_AGEMA_signal_11681), .B1_t (new_AGEMA_signal_11682), .B1_f (new_AGEMA_signal_11683), .Z0_t (SubBytesIns_Inst_Sbox_15_L5), .Z0_f (new_AGEMA_signal_12281), .Z1_t (new_AGEMA_signal_12282), .Z1_f (new_AGEMA_signal_12283) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M62), .A0_f (new_AGEMA_signal_12269), .A1_t (new_AGEMA_signal_12270), .A1_f (new_AGEMA_signal_12271), .B0_t (SubBytesIns_Inst_Sbox_15_L5), .B0_f (new_AGEMA_signal_12281), .B1_t (new_AGEMA_signal_12282), .B1_f (new_AGEMA_signal_12283), .Z0_t (SubBytesIns_Inst_Sbox_15_L6), .Z0_f (new_AGEMA_signal_12812), .Z1_t (new_AGEMA_signal_12813), .Z1_f (new_AGEMA_signal_12814) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M46), .A0_f (new_AGEMA_signal_11663), .A1_t (new_AGEMA_signal_11664), .A1_f (new_AGEMA_signal_11665), .B0_t (SubBytesIns_Inst_Sbox_15_L3), .B0_f (new_AGEMA_signal_12275), .B1_t (new_AGEMA_signal_12276), .B1_f (new_AGEMA_signal_12277), .Z0_t (SubBytesIns_Inst_Sbox_15_L7), .Z0_f (new_AGEMA_signal_12815), .Z1_t (new_AGEMA_signal_12816), .Z1_f (new_AGEMA_signal_12817) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M51), .A0_f (new_AGEMA_signal_10961), .A1_t (new_AGEMA_signal_10962), .A1_f (new_AGEMA_signal_10963), .B0_t (SubBytesIns_Inst_Sbox_15_M59), .B0_f (new_AGEMA_signal_10970), .B1_t (new_AGEMA_signal_10971), .B1_f (new_AGEMA_signal_10972), .Z0_t (SubBytesIns_Inst_Sbox_15_L8), .Z0_f (new_AGEMA_signal_11690), .Z1_t (new_AGEMA_signal_11691), .Z1_f (new_AGEMA_signal_11692) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M52), .A0_f (new_AGEMA_signal_11669), .A1_t (new_AGEMA_signal_11670), .A1_f (new_AGEMA_signal_11671), .B0_t (SubBytesIns_Inst_Sbox_15_M53), .B0_f (new_AGEMA_signal_12266), .B1_t (new_AGEMA_signal_12267), .B1_f (new_AGEMA_signal_12268), .Z0_t (SubBytesIns_Inst_Sbox_15_L9), .Z0_f (new_AGEMA_signal_12818), .Z1_t (new_AGEMA_signal_12819), .Z1_f (new_AGEMA_signal_12820) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M53), .A0_f (new_AGEMA_signal_12266), .A1_t (new_AGEMA_signal_12267), .A1_f (new_AGEMA_signal_12268), .B0_t (SubBytesIns_Inst_Sbox_15_L4), .B0_f (new_AGEMA_signal_12278), .B1_t (new_AGEMA_signal_12279), .B1_f (new_AGEMA_signal_12280), .Z0_t (SubBytesIns_Inst_Sbox_15_L10), .Z0_f (new_AGEMA_signal_12821), .Z1_t (new_AGEMA_signal_12822), .Z1_f (new_AGEMA_signal_12823) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M60), .A0_f (new_AGEMA_signal_10973), .A1_t (new_AGEMA_signal_10974), .A1_f (new_AGEMA_signal_10975), .B0_t (SubBytesIns_Inst_Sbox_15_L2), .B0_f (new_AGEMA_signal_12272), .B1_t (new_AGEMA_signal_12273), .B1_f (new_AGEMA_signal_12274), .Z0_t (SubBytesIns_Inst_Sbox_15_L11), .Z0_f (new_AGEMA_signal_12824), .Z1_t (new_AGEMA_signal_12825), .Z1_f (new_AGEMA_signal_12826) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M48), .A0_f (new_AGEMA_signal_10955), .A1_t (new_AGEMA_signal_10956), .A1_f (new_AGEMA_signal_10957), .B0_t (SubBytesIns_Inst_Sbox_15_M51), .B0_f (new_AGEMA_signal_10961), .B1_t (new_AGEMA_signal_10962), .B1_f (new_AGEMA_signal_10963), .Z0_t (SubBytesIns_Inst_Sbox_15_L12), .Z0_f (new_AGEMA_signal_11693), .Z1_t (new_AGEMA_signal_11694), .Z1_f (new_AGEMA_signal_11695) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M50), .A0_f (new_AGEMA_signal_10958), .A1_t (new_AGEMA_signal_10959), .A1_f (new_AGEMA_signal_10960), .B0_t (SubBytesIns_Inst_Sbox_15_L0), .B0_f (new_AGEMA_signal_12809), .B1_t (new_AGEMA_signal_12810), .B1_f (new_AGEMA_signal_12811), .Z0_t (SubBytesIns_Inst_Sbox_15_L13), .Z0_f (new_AGEMA_signal_13463), .Z1_t (new_AGEMA_signal_13464), .Z1_f (new_AGEMA_signal_13465) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M52), .A0_f (new_AGEMA_signal_11669), .A1_t (new_AGEMA_signal_11670), .A1_f (new_AGEMA_signal_11671), .B0_t (SubBytesIns_Inst_Sbox_15_M61), .B0_f (new_AGEMA_signal_11681), .B1_t (new_AGEMA_signal_11682), .B1_f (new_AGEMA_signal_11683), .Z0_t (SubBytesIns_Inst_Sbox_15_L14), .Z0_f (new_AGEMA_signal_12284), .Z1_t (new_AGEMA_signal_12285), .Z1_f (new_AGEMA_signal_12286) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M55), .A0_f (new_AGEMA_signal_11675), .A1_t (new_AGEMA_signal_11676), .A1_f (new_AGEMA_signal_11677), .B0_t (SubBytesIns_Inst_Sbox_15_L1), .B0_f (new_AGEMA_signal_11687), .B1_t (new_AGEMA_signal_11688), .B1_f (new_AGEMA_signal_11689), .Z0_t (SubBytesIns_Inst_Sbox_15_L15), .Z0_f (new_AGEMA_signal_12287), .Z1_t (new_AGEMA_signal_12288), .Z1_f (new_AGEMA_signal_12289) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M56), .A0_f (new_AGEMA_signal_10964), .A1_t (new_AGEMA_signal_10965), .A1_f (new_AGEMA_signal_10966), .B0_t (SubBytesIns_Inst_Sbox_15_L0), .B0_f (new_AGEMA_signal_12809), .B1_t (new_AGEMA_signal_12810), .B1_f (new_AGEMA_signal_12811), .Z0_t (SubBytesIns_Inst_Sbox_15_L16), .Z0_f (new_AGEMA_signal_13466), .Z1_t (new_AGEMA_signal_13467), .Z1_f (new_AGEMA_signal_13468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M57), .A0_f (new_AGEMA_signal_10967), .A1_t (new_AGEMA_signal_10968), .A1_f (new_AGEMA_signal_10969), .B0_t (SubBytesIns_Inst_Sbox_15_L1), .B0_f (new_AGEMA_signal_11687), .B1_t (new_AGEMA_signal_11688), .B1_f (new_AGEMA_signal_11689), .Z0_t (SubBytesIns_Inst_Sbox_15_L17), .Z0_f (new_AGEMA_signal_12290), .Z1_t (new_AGEMA_signal_12291), .Z1_f (new_AGEMA_signal_12292) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M58), .A0_f (new_AGEMA_signal_11678), .A1_t (new_AGEMA_signal_11679), .A1_f (new_AGEMA_signal_11680), .B0_t (SubBytesIns_Inst_Sbox_15_L8), .B0_f (new_AGEMA_signal_11690), .B1_t (new_AGEMA_signal_11691), .B1_f (new_AGEMA_signal_11692), .Z0_t (SubBytesIns_Inst_Sbox_15_L18), .Z0_f (new_AGEMA_signal_12293), .Z1_t (new_AGEMA_signal_12294), .Z1_f (new_AGEMA_signal_12295) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M63), .A0_f (new_AGEMA_signal_11684), .A1_t (new_AGEMA_signal_11685), .A1_f (new_AGEMA_signal_11686), .B0_t (SubBytesIns_Inst_Sbox_15_L4), .B0_f (new_AGEMA_signal_12278), .B1_t (new_AGEMA_signal_12279), .B1_f (new_AGEMA_signal_12280), .Z0_t (SubBytesIns_Inst_Sbox_15_L19), .Z0_f (new_AGEMA_signal_12827), .Z1_t (new_AGEMA_signal_12828), .Z1_f (new_AGEMA_signal_12829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L0), .A0_f (new_AGEMA_signal_12809), .A1_t (new_AGEMA_signal_12810), .A1_f (new_AGEMA_signal_12811), .B0_t (SubBytesIns_Inst_Sbox_15_L1), .B0_f (new_AGEMA_signal_11687), .B1_t (new_AGEMA_signal_11688), .B1_f (new_AGEMA_signal_11689), .Z0_t (SubBytesIns_Inst_Sbox_15_L20), .Z0_f (new_AGEMA_signal_13469), .Z1_t (new_AGEMA_signal_13470), .Z1_f (new_AGEMA_signal_13471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L1), .A0_f (new_AGEMA_signal_11687), .A1_t (new_AGEMA_signal_11688), .A1_f (new_AGEMA_signal_11689), .B0_t (SubBytesIns_Inst_Sbox_15_L7), .B0_f (new_AGEMA_signal_12815), .B1_t (new_AGEMA_signal_12816), .B1_f (new_AGEMA_signal_12817), .Z0_t (SubBytesIns_Inst_Sbox_15_L21), .Z0_f (new_AGEMA_signal_13472), .Z1_t (new_AGEMA_signal_13473), .Z1_f (new_AGEMA_signal_13474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L3), .A0_f (new_AGEMA_signal_12275), .A1_t (new_AGEMA_signal_12276), .A1_f (new_AGEMA_signal_12277), .B0_t (SubBytesIns_Inst_Sbox_15_L12), .B0_f (new_AGEMA_signal_11693), .B1_t (new_AGEMA_signal_11694), .B1_f (new_AGEMA_signal_11695), .Z0_t (SubBytesIns_Inst_Sbox_15_L22), .Z0_f (new_AGEMA_signal_12830), .Z1_t (new_AGEMA_signal_12831), .Z1_f (new_AGEMA_signal_12832) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L18), .A0_f (new_AGEMA_signal_12293), .A1_t (new_AGEMA_signal_12294), .A1_f (new_AGEMA_signal_12295), .B0_t (SubBytesIns_Inst_Sbox_15_L2), .B0_f (new_AGEMA_signal_12272), .B1_t (new_AGEMA_signal_12273), .B1_f (new_AGEMA_signal_12274), .Z0_t (SubBytesIns_Inst_Sbox_15_L23), .Z0_f (new_AGEMA_signal_12833), .Z1_t (new_AGEMA_signal_12834), .Z1_f (new_AGEMA_signal_12835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L15), .A0_f (new_AGEMA_signal_12287), .A1_t (new_AGEMA_signal_12288), .A1_f (new_AGEMA_signal_12289), .B0_t (SubBytesIns_Inst_Sbox_15_L9), .B0_f (new_AGEMA_signal_12818), .B1_t (new_AGEMA_signal_12819), .B1_f (new_AGEMA_signal_12820), .Z0_t (SubBytesIns_Inst_Sbox_15_L24), .Z0_f (new_AGEMA_signal_13475), .Z1_t (new_AGEMA_signal_13476), .Z1_f (new_AGEMA_signal_13477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L6), .A0_f (new_AGEMA_signal_12812), .A1_t (new_AGEMA_signal_12813), .A1_f (new_AGEMA_signal_12814), .B0_t (SubBytesIns_Inst_Sbox_15_L10), .B0_f (new_AGEMA_signal_12821), .B1_t (new_AGEMA_signal_12822), .B1_f (new_AGEMA_signal_12823), .Z0_t (SubBytesIns_Inst_Sbox_15_L25), .Z0_f (new_AGEMA_signal_13478), .Z1_t (new_AGEMA_signal_13479), .Z1_f (new_AGEMA_signal_13480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L7), .A0_f (new_AGEMA_signal_12815), .A1_t (new_AGEMA_signal_12816), .A1_f (new_AGEMA_signal_12817), .B0_t (SubBytesIns_Inst_Sbox_15_L9), .B0_f (new_AGEMA_signal_12818), .B1_t (new_AGEMA_signal_12819), .B1_f (new_AGEMA_signal_12820), .Z0_t (SubBytesIns_Inst_Sbox_15_L26), .Z0_f (new_AGEMA_signal_13481), .Z1_t (new_AGEMA_signal_13482), .Z1_f (new_AGEMA_signal_13483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L8), .A0_f (new_AGEMA_signal_11690), .A1_t (new_AGEMA_signal_11691), .A1_f (new_AGEMA_signal_11692), .B0_t (SubBytesIns_Inst_Sbox_15_L10), .B0_f (new_AGEMA_signal_12821), .B1_t (new_AGEMA_signal_12822), .B1_f (new_AGEMA_signal_12823), .Z0_t (SubBytesIns_Inst_Sbox_15_L27), .Z0_f (new_AGEMA_signal_13484), .Z1_t (new_AGEMA_signal_13485), .Z1_f (new_AGEMA_signal_13486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L11), .A0_f (new_AGEMA_signal_12824), .A1_t (new_AGEMA_signal_12825), .A1_f (new_AGEMA_signal_12826), .B0_t (SubBytesIns_Inst_Sbox_15_L14), .B0_f (new_AGEMA_signal_12284), .B1_t (new_AGEMA_signal_12285), .B1_f (new_AGEMA_signal_12286), .Z0_t (SubBytesIns_Inst_Sbox_15_L28), .Z0_f (new_AGEMA_signal_13487), .Z1_t (new_AGEMA_signal_13488), .Z1_f (new_AGEMA_signal_13489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L11), .A0_f (new_AGEMA_signal_12824), .A1_t (new_AGEMA_signal_12825), .A1_f (new_AGEMA_signal_12826), .B0_t (SubBytesIns_Inst_Sbox_15_L17), .B0_f (new_AGEMA_signal_12290), .B1_t (new_AGEMA_signal_12291), .B1_f (new_AGEMA_signal_12292), .Z0_t (SubBytesIns_Inst_Sbox_15_L29), .Z0_f (new_AGEMA_signal_13490), .Z1_t (new_AGEMA_signal_13491), .Z1_f (new_AGEMA_signal_13492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L6), .A0_f (new_AGEMA_signal_12812), .A1_t (new_AGEMA_signal_12813), .A1_f (new_AGEMA_signal_12814), .B0_t (SubBytesIns_Inst_Sbox_15_L24), .B0_f (new_AGEMA_signal_13475), .B1_t (new_AGEMA_signal_13476), .B1_f (new_AGEMA_signal_13477), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .Z0_f (new_AGEMA_signal_13955), .Z1_t (new_AGEMA_signal_13956), .Z1_f (new_AGEMA_signal_13957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L16), .A0_f (new_AGEMA_signal_13466), .A1_t (new_AGEMA_signal_13467), .A1_f (new_AGEMA_signal_13468), .B0_t (SubBytesIns_Inst_Sbox_15_L26), .B0_f (new_AGEMA_signal_13481), .B1_t (new_AGEMA_signal_13482), .B1_f (new_AGEMA_signal_13483), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .Z0_f (new_AGEMA_signal_13958), .Z1_t (new_AGEMA_signal_13959), .Z1_f (new_AGEMA_signal_13960) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L19), .A0_f (new_AGEMA_signal_12827), .A1_t (new_AGEMA_signal_12828), .A1_f (new_AGEMA_signal_12829), .B0_t (SubBytesIns_Inst_Sbox_15_L28), .B0_f (new_AGEMA_signal_13487), .B1_t (new_AGEMA_signal_13488), .B1_f (new_AGEMA_signal_13489), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .Z0_f (new_AGEMA_signal_13961), .Z1_t (new_AGEMA_signal_13962), .Z1_f (new_AGEMA_signal_13963) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L6), .A0_f (new_AGEMA_signal_12812), .A1_t (new_AGEMA_signal_12813), .A1_f (new_AGEMA_signal_12814), .B0_t (SubBytesIns_Inst_Sbox_15_L21), .B0_f (new_AGEMA_signal_13472), .B1_t (new_AGEMA_signal_13473), .B1_f (new_AGEMA_signal_13474), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .Z0_f (new_AGEMA_signal_13964), .Z1_t (new_AGEMA_signal_13965), .Z1_f (new_AGEMA_signal_13966) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L20), .A0_f (new_AGEMA_signal_13469), .A1_t (new_AGEMA_signal_13470), .A1_f (new_AGEMA_signal_13471), .B0_t (SubBytesIns_Inst_Sbox_15_L22), .B0_f (new_AGEMA_signal_12830), .B1_t (new_AGEMA_signal_12831), .B1_f (new_AGEMA_signal_12832), .Z0_t (MixColumnsInput[123]), .Z0_f (new_AGEMA_signal_13967), .Z1_t (new_AGEMA_signal_13968), .Z1_f (new_AGEMA_signal_13969) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L25), .A0_f (new_AGEMA_signal_13478), .A1_t (new_AGEMA_signal_13479), .A1_f (new_AGEMA_signal_13480), .B0_t (SubBytesIns_Inst_Sbox_15_L29), .B0_f (new_AGEMA_signal_13490), .B1_t (new_AGEMA_signal_13491), .B1_f (new_AGEMA_signal_13492), .Z0_t (MixColumnsInput[122]), .Z0_f (new_AGEMA_signal_13970), .Z1_t (new_AGEMA_signal_13971), .Z1_f (new_AGEMA_signal_13972) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L13), .A0_f (new_AGEMA_signal_13463), .A1_t (new_AGEMA_signal_13464), .A1_f (new_AGEMA_signal_13465), .B0_t (SubBytesIns_Inst_Sbox_15_L27), .B0_f (new_AGEMA_signal_13484), .B1_t (new_AGEMA_signal_13485), .B1_f (new_AGEMA_signal_13486), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .Z0_f (new_AGEMA_signal_13973), .Z1_t (new_AGEMA_signal_13974), .Z1_f (new_AGEMA_signal_13975) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L6), .A0_f (new_AGEMA_signal_12812), .A1_t (new_AGEMA_signal_12813), .A1_f (new_AGEMA_signal_12814), .B0_t (SubBytesIns_Inst_Sbox_15_L23), .B0_f (new_AGEMA_signal_12833), .B1_t (new_AGEMA_signal_12834), .B1_f (new_AGEMA_signal_12835), .Z0_t (MixColumnsInput[120]), .Z0_f (new_AGEMA_signal_13493), .Z1_t (new_AGEMA_signal_13494), .Z1_f (new_AGEMA_signal_13495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U96 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n192), .A0_f (new_AGEMA_signal_15812), .A1_t (new_AGEMA_signal_15813), .A1_f (new_AGEMA_signal_15814), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13868), .B1_t (new_AGEMA_signal_13869), .B1_f (new_AGEMA_signal_13870), .Z0_t (MixColumnsOutput[105]), .Z0_f (new_AGEMA_signal_16811), .Z1_t (new_AGEMA_signal_16812), .Z1_f (new_AGEMA_signal_16813) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U95 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n191), .A0_f (new_AGEMA_signal_15128), .A1_t (new_AGEMA_signal_15129), .A1_f (new_AGEMA_signal_15130), .B0_t (MixColumnsIns_MixOneColumnInst_0_n190), .B0_f (new_AGEMA_signal_15116), .B1_t (new_AGEMA_signal_15117), .B1_f (new_AGEMA_signal_15118), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n192), .Z0_f (new_AGEMA_signal_15812), .Z1_t (new_AGEMA_signal_15813), .Z1_f (new_AGEMA_signal_15814) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U94 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n189), .A0_f (new_AGEMA_signal_15065), .A1_t (new_AGEMA_signal_15066), .A1_f (new_AGEMA_signal_15067), .B0_t (MixColumnsIns_MixOneColumnInst_0_n188), .B0_f (new_AGEMA_signal_14453), .B1_t (new_AGEMA_signal_14454), .B1_f (new_AGEMA_signal_14455), .Z0_t (MixColumnsOutput[104]), .Z0_f (new_AGEMA_signal_15815), .Z1_t (new_AGEMA_signal_15816), .Z1_f (new_AGEMA_signal_15817) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U93 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n187), .A0_f (new_AGEMA_signal_14483), .A1_t (new_AGEMA_signal_14484), .A1_f (new_AGEMA_signal_14485), .B0_t (MixColumnsInput[112]), .B0_f (new_AGEMA_signal_13328), .B1_t (new_AGEMA_signal_13329), .B1_f (new_AGEMA_signal_13330), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n189), .Z0_f (new_AGEMA_signal_15065), .Z1_t (new_AGEMA_signal_15066), .Z1_f (new_AGEMA_signal_15067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U92 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n186), .A0_f (new_AGEMA_signal_15068), .A1_t (new_AGEMA_signal_15069), .A1_f (new_AGEMA_signal_15070), .B0_t (MixColumnsIns_MixOneColumnInst_0_n185), .B0_f (new_AGEMA_signal_14426), .B1_t (new_AGEMA_signal_14427), .B1_f (new_AGEMA_signal_14428), .Z0_t (MixColumnsOutput[103]), .Z0_f (new_AGEMA_signal_15818), .Z1_t (new_AGEMA_signal_15819), .Z1_f (new_AGEMA_signal_15820) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U91 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n184), .A0_f (new_AGEMA_signal_14459), .A1_t (new_AGEMA_signal_14460), .A1_f (new_AGEMA_signal_14461), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B0_f (new_AGEMA_signal_13745), .B1_t (new_AGEMA_signal_13746), .B1_f (new_AGEMA_signal_13747), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n186), .Z0_f (new_AGEMA_signal_15068), .Z1_t (new_AGEMA_signal_15069), .Z1_f (new_AGEMA_signal_15070) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U90 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n183), .A0_f (new_AGEMA_signal_15071), .A1_t (new_AGEMA_signal_15072), .A1_f (new_AGEMA_signal_15073), .B0_t (MixColumnsIns_MixOneColumnInst_0_n182), .B0_f (new_AGEMA_signal_14429), .B1_t (new_AGEMA_signal_14430), .B1_f (new_AGEMA_signal_14431), .Z0_t (MixColumnsOutput[102]), .Z0_f (new_AGEMA_signal_15821), .Z1_t (new_AGEMA_signal_15822), .Z1_f (new_AGEMA_signal_15823) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U89 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n181), .A0_f (new_AGEMA_signal_14465), .A1_t (new_AGEMA_signal_14466), .A1_f (new_AGEMA_signal_14467), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13748), .B1_t (new_AGEMA_signal_13749), .B1_f (new_AGEMA_signal_13750), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n183), .Z0_f (new_AGEMA_signal_15071), .Z1_t (new_AGEMA_signal_15072), .Z1_f (new_AGEMA_signal_15073) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U88 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n180), .A0_f (new_AGEMA_signal_15074), .A1_t (new_AGEMA_signal_15075), .A1_f (new_AGEMA_signal_15076), .B0_t (MixColumnsIns_MixOneColumnInst_0_n179), .B0_f (new_AGEMA_signal_14432), .B1_t (new_AGEMA_signal_14433), .B1_f (new_AGEMA_signal_14434), .Z0_t (MixColumnsOutput[101]), .Z0_f (new_AGEMA_signal_15824), .Z1_t (new_AGEMA_signal_15825), .Z1_f (new_AGEMA_signal_15826) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U87 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n178), .A0_f (new_AGEMA_signal_14471), .A1_t (new_AGEMA_signal_14472), .A1_f (new_AGEMA_signal_14473), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13751), .B1_t (new_AGEMA_signal_13752), .B1_f (new_AGEMA_signal_13753), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n180), .Z0_f (new_AGEMA_signal_15074), .Z1_t (new_AGEMA_signal_15075), .Z1_f (new_AGEMA_signal_15076) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U86 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n177), .A0_f (new_AGEMA_signal_15827), .A1_t (new_AGEMA_signal_15828), .A1_f (new_AGEMA_signal_15829), .B0_t (MixColumnsIns_MixOneColumnInst_0_n176), .B0_f (new_AGEMA_signal_15089), .B1_t (new_AGEMA_signal_15090), .B1_f (new_AGEMA_signal_15091), .Z0_t (MixColumnsOutput[100]), .Z0_f (new_AGEMA_signal_16814), .Z1_t (new_AGEMA_signal_16815), .Z1_f (new_AGEMA_signal_16816) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U85 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n175), .A0_f (new_AGEMA_signal_15146), .A1_t (new_AGEMA_signal_15147), .A1_f (new_AGEMA_signal_15148), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13754), .B1_t (new_AGEMA_signal_13755), .B1_f (new_AGEMA_signal_13756), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n177), .Z0_f (new_AGEMA_signal_15827), .Z1_t (new_AGEMA_signal_15828), .Z1_f (new_AGEMA_signal_15829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U84 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n174), .A0_f (new_AGEMA_signal_15830), .A1_t (new_AGEMA_signal_15831), .A1_f (new_AGEMA_signal_15832), .B0_t (MixColumnsIns_MixOneColumnInst_0_n173), .B0_f (new_AGEMA_signal_15092), .B1_t (new_AGEMA_signal_15093), .B1_f (new_AGEMA_signal_15094), .Z0_t (MixColumnsOutput[99]), .Z0_f (new_AGEMA_signal_16817), .Z1_t (new_AGEMA_signal_16818), .Z1_f (new_AGEMA_signal_16819) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U83 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n172), .A0_f (new_AGEMA_signal_15152), .A1_t (new_AGEMA_signal_15153), .A1_f (new_AGEMA_signal_15154), .B0_t (MixColumnsInput[107]), .B0_f (new_AGEMA_signal_13757), .B1_t (new_AGEMA_signal_13758), .B1_f (new_AGEMA_signal_13759), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n174), .Z0_f (new_AGEMA_signal_15830), .Z1_t (new_AGEMA_signal_15831), .Z1_f (new_AGEMA_signal_15832) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U82 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n171), .A0_f (new_AGEMA_signal_15077), .A1_t (new_AGEMA_signal_15078), .A1_f (new_AGEMA_signal_15079), .B0_t (MixColumnsIns_MixOneColumnInst_0_n185), .B0_f (new_AGEMA_signal_14426), .B1_t (new_AGEMA_signal_14427), .B1_f (new_AGEMA_signal_14428), .Z0_t (MixColumnsOutput[127]), .Z0_f (new_AGEMA_signal_15833), .Z1_t (new_AGEMA_signal_15834), .Z1_f (new_AGEMA_signal_15835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U81 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13850), .A1_t (new_AGEMA_signal_13851), .A1_f (new_AGEMA_signal_13852), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13958), .B1_t (new_AGEMA_signal_13959), .B1_f (new_AGEMA_signal_13960), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n185), .Z0_f (new_AGEMA_signal_14426), .Z1_t (new_AGEMA_signal_14427), .Z1_f (new_AGEMA_signal_14428) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U80 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13640), .A1_t (new_AGEMA_signal_13641), .A1_f (new_AGEMA_signal_13642), .B0_t (MixColumnsIns_MixOneColumnInst_0_n170), .B0_f (new_AGEMA_signal_14438), .B1_t (new_AGEMA_signal_14439), .B1_f (new_AGEMA_signal_14440), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n171), .Z0_f (new_AGEMA_signal_15077), .Z1_t (new_AGEMA_signal_15078), .Z1_f (new_AGEMA_signal_15079) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U79 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n169), .A0_f (new_AGEMA_signal_15080), .A1_t (new_AGEMA_signal_15081), .A1_f (new_AGEMA_signal_15082), .B0_t (MixColumnsIns_MixOneColumnInst_0_n182), .B0_f (new_AGEMA_signal_14429), .B1_t (new_AGEMA_signal_14430), .B1_f (new_AGEMA_signal_14431), .Z0_t (MixColumnsOutput[126]), .Z0_f (new_AGEMA_signal_15836), .Z1_t (new_AGEMA_signal_15837), .Z1_f (new_AGEMA_signal_15838) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U78 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .A0_f (new_AGEMA_signal_13853), .A1_t (new_AGEMA_signal_13854), .A1_f (new_AGEMA_signal_13855), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13961), .B1_t (new_AGEMA_signal_13962), .B1_f (new_AGEMA_signal_13963), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n182), .Z0_f (new_AGEMA_signal_14429), .Z1_t (new_AGEMA_signal_14430), .Z1_f (new_AGEMA_signal_14431) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U77 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13643), .A1_t (new_AGEMA_signal_13644), .A1_f (new_AGEMA_signal_13645), .B0_t (MixColumnsIns_MixOneColumnInst_0_n168), .B0_f (new_AGEMA_signal_14441), .B1_t (new_AGEMA_signal_14442), .B1_f (new_AGEMA_signal_14443), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n169), .Z0_f (new_AGEMA_signal_15080), .Z1_t (new_AGEMA_signal_15081), .Z1_f (new_AGEMA_signal_15082) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U76 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n167), .A0_f (new_AGEMA_signal_15083), .A1_t (new_AGEMA_signal_15084), .A1_f (new_AGEMA_signal_15085), .B0_t (MixColumnsIns_MixOneColumnInst_0_n166), .B0_f (new_AGEMA_signal_14435), .B1_t (new_AGEMA_signal_14436), .B1_f (new_AGEMA_signal_14437), .Z0_t (MixColumnsOutput[98]), .Z0_f (new_AGEMA_signal_15839), .Z1_t (new_AGEMA_signal_15840), .Z1_f (new_AGEMA_signal_15841) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U75 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n165), .A0_f (new_AGEMA_signal_14477), .A1_t (new_AGEMA_signal_14478), .A1_f (new_AGEMA_signal_14479), .B0_t (MixColumnsInput[106]), .B0_f (new_AGEMA_signal_13760), .B1_t (new_AGEMA_signal_13761), .B1_f (new_AGEMA_signal_13762), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n167), .Z0_f (new_AGEMA_signal_15083), .Z1_t (new_AGEMA_signal_15084), .Z1_f (new_AGEMA_signal_15085) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U74 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n164), .A0_f (new_AGEMA_signal_15086), .A1_t (new_AGEMA_signal_15087), .A1_f (new_AGEMA_signal_15088), .B0_t (MixColumnsIns_MixOneColumnInst_0_n179), .B0_f (new_AGEMA_signal_14432), .B1_t (new_AGEMA_signal_14433), .B1_f (new_AGEMA_signal_14434), .Z0_t (MixColumnsOutput[125]), .Z0_f (new_AGEMA_signal_15842), .Z1_t (new_AGEMA_signal_15843), .Z1_f (new_AGEMA_signal_15844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U73 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .A0_f (new_AGEMA_signal_13856), .A1_t (new_AGEMA_signal_13857), .A1_f (new_AGEMA_signal_13858), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13964), .B1_t (new_AGEMA_signal_13965), .B1_f (new_AGEMA_signal_13966), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n179), .Z0_f (new_AGEMA_signal_14432), .Z1_t (new_AGEMA_signal_14433), .Z1_f (new_AGEMA_signal_14434) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U72 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13646), .A1_t (new_AGEMA_signal_13647), .A1_f (new_AGEMA_signal_13648), .B0_t (MixColumnsIns_MixOneColumnInst_0_n163), .B0_f (new_AGEMA_signal_14444), .B1_t (new_AGEMA_signal_14445), .B1_f (new_AGEMA_signal_14446), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n164), .Z0_f (new_AGEMA_signal_15086), .Z1_t (new_AGEMA_signal_15087), .Z1_f (new_AGEMA_signal_15088) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U71 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n162), .A0_f (new_AGEMA_signal_15845), .A1_t (new_AGEMA_signal_15846), .A1_f (new_AGEMA_signal_15847), .B0_t (MixColumnsIns_MixOneColumnInst_0_n176), .B0_f (new_AGEMA_signal_15089), .B1_t (new_AGEMA_signal_15090), .B1_f (new_AGEMA_signal_15091), .Z0_t (MixColumnsOutput[124]), .Z0_f (new_AGEMA_signal_16820), .Z1_t (new_AGEMA_signal_16821), .Z1_f (new_AGEMA_signal_16822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U70 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .A0_f (new_AGEMA_signal_13859), .A1_t (new_AGEMA_signal_13860), .A1_f (new_AGEMA_signal_13861), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]), .B0_f (new_AGEMA_signal_14486), .B1_t (new_AGEMA_signal_14487), .B1_f (new_AGEMA_signal_14488), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n176), .Z0_f (new_AGEMA_signal_15089), .Z1_t (new_AGEMA_signal_15090), .Z1_f (new_AGEMA_signal_15091) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U69 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13649), .A1_t (new_AGEMA_signal_13650), .A1_f (new_AGEMA_signal_13651), .B0_t (MixColumnsIns_MixOneColumnInst_0_n161), .B0_f (new_AGEMA_signal_15110), .B1_t (new_AGEMA_signal_15111), .B1_f (new_AGEMA_signal_15112), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n162), .Z0_f (new_AGEMA_signal_15845), .Z1_t (new_AGEMA_signal_15846), .Z1_f (new_AGEMA_signal_15847) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U68 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n160), .A0_f (new_AGEMA_signal_15848), .A1_t (new_AGEMA_signal_15849), .A1_f (new_AGEMA_signal_15850), .B0_t (MixColumnsIns_MixOneColumnInst_0_n173), .B0_f (new_AGEMA_signal_15092), .B1_t (new_AGEMA_signal_15093), .B1_f (new_AGEMA_signal_15094), .Z0_t (MixColumnsOutput[123]), .Z0_f (new_AGEMA_signal_16823), .Z1_t (new_AGEMA_signal_16824), .Z1_f (new_AGEMA_signal_16825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U67 ( .A0_t (MixColumnsInput[115]), .A0_f (new_AGEMA_signal_13862), .A1_t (new_AGEMA_signal_13863), .A1_f (new_AGEMA_signal_13864), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]), .B0_f (new_AGEMA_signal_14489), .B1_t (new_AGEMA_signal_14490), .B1_f (new_AGEMA_signal_14491), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n173), .Z0_f (new_AGEMA_signal_15092), .Z1_t (new_AGEMA_signal_15093), .Z1_f (new_AGEMA_signal_15094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U66 ( .A0_t (MixColumnsInput[99]), .A0_f (new_AGEMA_signal_13652), .A1_t (new_AGEMA_signal_13653), .A1_f (new_AGEMA_signal_13654), .B0_t (MixColumnsIns_MixOneColumnInst_0_n159), .B0_f (new_AGEMA_signal_15119), .B1_t (new_AGEMA_signal_15120), .B1_f (new_AGEMA_signal_15121), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n160), .Z0_f (new_AGEMA_signal_15848), .Z1_t (new_AGEMA_signal_15849), .Z1_f (new_AGEMA_signal_15850) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U65 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n158), .A0_f (new_AGEMA_signal_15095), .A1_t (new_AGEMA_signal_15096), .A1_f (new_AGEMA_signal_15097), .B0_t (MixColumnsIns_MixOneColumnInst_0_n166), .B0_f (new_AGEMA_signal_14435), .B1_t (new_AGEMA_signal_14436), .B1_f (new_AGEMA_signal_14437), .Z0_t (MixColumnsOutput[122]), .Z0_f (new_AGEMA_signal_15851), .Z1_t (new_AGEMA_signal_15852), .Z1_f (new_AGEMA_signal_15853) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U64 ( .A0_t (MixColumnsInput[114]), .A0_f (new_AGEMA_signal_13865), .A1_t (new_AGEMA_signal_13866), .A1_f (new_AGEMA_signal_13867), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13973), .B1_t (new_AGEMA_signal_13974), .B1_f (new_AGEMA_signal_13975), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n166), .Z0_f (new_AGEMA_signal_14435), .Z1_t (new_AGEMA_signal_14436), .Z1_f (new_AGEMA_signal_14437) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U63 ( .A0_t (MixColumnsInput[98]), .A0_f (new_AGEMA_signal_13655), .A1_t (new_AGEMA_signal_13656), .A1_f (new_AGEMA_signal_13657), .B0_t (MixColumnsIns_MixOneColumnInst_0_n157), .B0_f (new_AGEMA_signal_14447), .B1_t (new_AGEMA_signal_14448), .B1_f (new_AGEMA_signal_14449), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n158), .Z0_f (new_AGEMA_signal_15095), .Z1_t (new_AGEMA_signal_15096), .Z1_f (new_AGEMA_signal_15097) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U62 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n156), .A0_f (new_AGEMA_signal_15854), .A1_t (new_AGEMA_signal_15855), .A1_f (new_AGEMA_signal_15856), .B0_t (MixColumnsIns_MixOneColumnInst_0_n155), .B0_f (new_AGEMA_signal_15113), .B1_t (new_AGEMA_signal_15114), .B1_f (new_AGEMA_signal_15115), .Z0_t (MixColumnsOutput[121]), .Z0_f (new_AGEMA_signal_16826), .Z1_t (new_AGEMA_signal_16827), .Z1_f (new_AGEMA_signal_16828) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U61 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .A0_f (new_AGEMA_signal_13658), .A1_t (new_AGEMA_signal_13659), .A1_f (new_AGEMA_signal_13660), .B0_t (MixColumnsIns_MixOneColumnInst_0_n154), .B0_f (new_AGEMA_signal_15125), .B1_t (new_AGEMA_signal_15126), .B1_f (new_AGEMA_signal_15127), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n156), .Z0_f (new_AGEMA_signal_15854), .Z1_t (new_AGEMA_signal_15855), .Z1_f (new_AGEMA_signal_15856) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U60 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n153), .A0_f (new_AGEMA_signal_15098), .A1_t (new_AGEMA_signal_15099), .A1_f (new_AGEMA_signal_15100), .B0_t (MixColumnsIns_MixOneColumnInst_0_n152), .B0_f (new_AGEMA_signal_14450), .B1_t (new_AGEMA_signal_14451), .B1_f (new_AGEMA_signal_14452), .Z0_t (MixColumnsOutput[120]), .Z0_f (new_AGEMA_signal_15857), .Z1_t (new_AGEMA_signal_15858), .Z1_f (new_AGEMA_signal_15859) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U59 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n151), .A0_f (new_AGEMA_signal_14480), .A1_t (new_AGEMA_signal_14481), .A1_f (new_AGEMA_signal_14482), .B0_t (MixColumnsInput[96]), .B0_f (new_AGEMA_signal_12998), .B1_t (new_AGEMA_signal_12999), .B1_f (new_AGEMA_signal_13000), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n153), .Z0_f (new_AGEMA_signal_15098), .Z1_t (new_AGEMA_signal_15099), .Z1_f (new_AGEMA_signal_15100) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U58 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n150), .A0_f (new_AGEMA_signal_15101), .A1_t (new_AGEMA_signal_15102), .A1_f (new_AGEMA_signal_15103), .B0_t (MixColumnsIns_MixOneColumnInst_0_n170), .B0_f (new_AGEMA_signal_14438), .B1_t (new_AGEMA_signal_14439), .B1_f (new_AGEMA_signal_14440), .Z0_t (MixColumnsOutput[119]), .Z0_f (new_AGEMA_signal_15860), .Z1_t (new_AGEMA_signal_15861), .Z1_f (new_AGEMA_signal_15862) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U57 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13745), .A1_t (new_AGEMA_signal_13746), .A1_f (new_AGEMA_signal_13747), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13853), .B1_t (new_AGEMA_signal_13854), .B1_f (new_AGEMA_signal_13855), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n170), .Z0_f (new_AGEMA_signal_14438), .Z1_t (new_AGEMA_signal_14439), .Z1_f (new_AGEMA_signal_14440) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U56 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13955), .A1_t (new_AGEMA_signal_13956), .A1_f (new_AGEMA_signal_13957), .B0_t (MixColumnsIns_MixOneColumnInst_0_n149), .B0_f (new_AGEMA_signal_14456), .B1_t (new_AGEMA_signal_14457), .B1_f (new_AGEMA_signal_14458), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n150), .Z0_f (new_AGEMA_signal_15101), .Z1_t (new_AGEMA_signal_15102), .Z1_f (new_AGEMA_signal_15103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U55 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n148), .A0_f (new_AGEMA_signal_15104), .A1_t (new_AGEMA_signal_15105), .A1_f (new_AGEMA_signal_15106), .B0_t (MixColumnsIns_MixOneColumnInst_0_n168), .B0_f (new_AGEMA_signal_14441), .B1_t (new_AGEMA_signal_14442), .B1_f (new_AGEMA_signal_14443), .Z0_t (MixColumnsOutput[118]), .Z0_f (new_AGEMA_signal_15863), .Z1_t (new_AGEMA_signal_15864), .Z1_f (new_AGEMA_signal_15865) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U54 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .A0_f (new_AGEMA_signal_13748), .A1_t (new_AGEMA_signal_13749), .A1_f (new_AGEMA_signal_13750), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13856), .B1_t (new_AGEMA_signal_13857), .B1_f (new_AGEMA_signal_13858), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n168), .Z0_f (new_AGEMA_signal_14441), .Z1_t (new_AGEMA_signal_14442), .Z1_f (new_AGEMA_signal_14443) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U53 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .A0_f (new_AGEMA_signal_13958), .A1_t (new_AGEMA_signal_13959), .A1_f (new_AGEMA_signal_13960), .B0_t (MixColumnsIns_MixOneColumnInst_0_n147), .B0_f (new_AGEMA_signal_14462), .B1_t (new_AGEMA_signal_14463), .B1_f (new_AGEMA_signal_14464), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n148), .Z0_f (new_AGEMA_signal_15104), .Z1_t (new_AGEMA_signal_15105), .Z1_f (new_AGEMA_signal_15106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U52 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n146), .A0_f (new_AGEMA_signal_15107), .A1_t (new_AGEMA_signal_15108), .A1_f (new_AGEMA_signal_15109), .B0_t (MixColumnsIns_MixOneColumnInst_0_n163), .B0_f (new_AGEMA_signal_14444), .B1_t (new_AGEMA_signal_14445), .B1_f (new_AGEMA_signal_14446), .Z0_t (MixColumnsOutput[117]), .Z0_f (new_AGEMA_signal_15866), .Z1_t (new_AGEMA_signal_15867), .Z1_f (new_AGEMA_signal_15868) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U51 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .A0_f (new_AGEMA_signal_13751), .A1_t (new_AGEMA_signal_13752), .A1_f (new_AGEMA_signal_13753), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13859), .B1_t (new_AGEMA_signal_13860), .B1_f (new_AGEMA_signal_13861), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n163), .Z0_f (new_AGEMA_signal_14444), .Z1_t (new_AGEMA_signal_14445), .Z1_f (new_AGEMA_signal_14446) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U50 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .A0_f (new_AGEMA_signal_13961), .A1_t (new_AGEMA_signal_13962), .A1_f (new_AGEMA_signal_13963), .B0_t (MixColumnsIns_MixOneColumnInst_0_n145), .B0_f (new_AGEMA_signal_14468), .B1_t (new_AGEMA_signal_14469), .B1_f (new_AGEMA_signal_14470), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n146), .Z0_f (new_AGEMA_signal_15107), .Z1_t (new_AGEMA_signal_15108), .Z1_f (new_AGEMA_signal_15109) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U49 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n144), .A0_f (new_AGEMA_signal_15869), .A1_t (new_AGEMA_signal_15870), .A1_f (new_AGEMA_signal_15871), .B0_t (MixColumnsIns_MixOneColumnInst_0_n161), .B0_f (new_AGEMA_signal_15110), .B1_t (new_AGEMA_signal_15111), .B1_f (new_AGEMA_signal_15112), .Z0_t (MixColumnsOutput[116]), .Z0_f (new_AGEMA_signal_16829), .Z1_t (new_AGEMA_signal_16830), .Z1_f (new_AGEMA_signal_16831) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U48 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .A0_f (new_AGEMA_signal_13754), .A1_t (new_AGEMA_signal_13755), .A1_f (new_AGEMA_signal_13756), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]), .B0_f (new_AGEMA_signal_14495), .B1_t (new_AGEMA_signal_14496), .B1_f (new_AGEMA_signal_14497), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n161), .Z0_f (new_AGEMA_signal_15110), .Z1_t (new_AGEMA_signal_15111), .Z1_f (new_AGEMA_signal_15112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U47 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .A0_f (new_AGEMA_signal_13964), .A1_t (new_AGEMA_signal_13965), .A1_f (new_AGEMA_signal_13966), .B0_t (MixColumnsIns_MixOneColumnInst_0_n143), .B0_f (new_AGEMA_signal_15143), .B1_t (new_AGEMA_signal_15144), .B1_f (new_AGEMA_signal_15145), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n144), .Z0_f (new_AGEMA_signal_15869), .Z1_t (new_AGEMA_signal_15870), .Z1_f (new_AGEMA_signal_15871) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U46 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n142), .A0_f (new_AGEMA_signal_15872), .A1_t (new_AGEMA_signal_15873), .A1_f (new_AGEMA_signal_15874), .B0_t (MixColumnsIns_MixOneColumnInst_0_n155), .B0_f (new_AGEMA_signal_15113), .B1_t (new_AGEMA_signal_15114), .B1_f (new_AGEMA_signal_15115), .Z0_t (MixColumnsOutput[97]), .Z0_f (new_AGEMA_signal_16832), .Z1_t (new_AGEMA_signal_16833), .Z1_f (new_AGEMA_signal_16834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U45 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .A0_f (new_AGEMA_signal_13868), .A1_t (new_AGEMA_signal_13869), .A1_f (new_AGEMA_signal_13870), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]), .B0_f (new_AGEMA_signal_14492), .B1_t (new_AGEMA_signal_14493), .B1_f (new_AGEMA_signal_14494), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n155), .Z0_f (new_AGEMA_signal_15113), .Z1_t (new_AGEMA_signal_15114), .Z1_f (new_AGEMA_signal_15115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U44 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .A0_f (new_AGEMA_signal_13763), .A1_t (new_AGEMA_signal_13764), .A1_f (new_AGEMA_signal_13765), .B0_t (MixColumnsIns_MixOneColumnInst_0_n190), .B0_f (new_AGEMA_signal_15116), .B1_t (new_AGEMA_signal_15117), .B1_f (new_AGEMA_signal_15118), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n142), .Z0_f (new_AGEMA_signal_15872), .Z1_t (new_AGEMA_signal_15873), .Z1_f (new_AGEMA_signal_15874) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U43 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .A0_f (new_AGEMA_signal_13973), .A1_t (new_AGEMA_signal_13974), .A1_f (new_AGEMA_signal_13975), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]), .B0_f (new_AGEMA_signal_14519), .B1_t (new_AGEMA_signal_14520), .B1_f (new_AGEMA_signal_14521), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n190), .Z0_f (new_AGEMA_signal_15116), .Z1_t (new_AGEMA_signal_15117), .Z1_f (new_AGEMA_signal_15118) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U42 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n141), .A0_f (new_AGEMA_signal_15875), .A1_t (new_AGEMA_signal_15876), .A1_f (new_AGEMA_signal_15877), .B0_t (MixColumnsIns_MixOneColumnInst_0_n159), .B0_f (new_AGEMA_signal_15119), .B1_t (new_AGEMA_signal_15120), .B1_f (new_AGEMA_signal_15121), .Z0_t (MixColumnsOutput[115]), .Z0_f (new_AGEMA_signal_16835), .Z1_t (new_AGEMA_signal_16836), .Z1_f (new_AGEMA_signal_16837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U41 ( .A0_t (MixColumnsInput[107]), .A0_f (new_AGEMA_signal_13757), .A1_t (new_AGEMA_signal_13758), .A1_f (new_AGEMA_signal_13759), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]), .B0_f (new_AGEMA_signal_14498), .B1_t (new_AGEMA_signal_14499), .B1_f (new_AGEMA_signal_14500), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n159), .Z0_f (new_AGEMA_signal_15119), .Z1_t (new_AGEMA_signal_15120), .Z1_f (new_AGEMA_signal_15121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U40 ( .A0_t (MixColumnsInput[123]), .A0_f (new_AGEMA_signal_13967), .A1_t (new_AGEMA_signal_13968), .A1_f (new_AGEMA_signal_13969), .B0_t (MixColumnsIns_MixOneColumnInst_0_n140), .B0_f (new_AGEMA_signal_15149), .B1_t (new_AGEMA_signal_15150), .B1_f (new_AGEMA_signal_15151), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n141), .Z0_f (new_AGEMA_signal_15875), .Z1_t (new_AGEMA_signal_15876), .Z1_f (new_AGEMA_signal_15877) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U39 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n139), .A0_f (new_AGEMA_signal_15122), .A1_t (new_AGEMA_signal_15123), .A1_f (new_AGEMA_signal_15124), .B0_t (MixColumnsIns_MixOneColumnInst_0_n157), .B0_f (new_AGEMA_signal_14447), .B1_t (new_AGEMA_signal_14448), .B1_f (new_AGEMA_signal_14449), .Z0_t (MixColumnsOutput[114]), .Z0_f (new_AGEMA_signal_15878), .Z1_t (new_AGEMA_signal_15879), .Z1_f (new_AGEMA_signal_15880) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U38 ( .A0_t (MixColumnsInput[106]), .A0_f (new_AGEMA_signal_13760), .A1_t (new_AGEMA_signal_13761), .A1_f (new_AGEMA_signal_13762), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13868), .B1_t (new_AGEMA_signal_13869), .B1_f (new_AGEMA_signal_13870), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n157), .Z0_f (new_AGEMA_signal_14447), .Z1_t (new_AGEMA_signal_14448), .Z1_f (new_AGEMA_signal_14449) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U37 ( .A0_t (MixColumnsInput[122]), .A0_f (new_AGEMA_signal_13970), .A1_t (new_AGEMA_signal_13971), .A1_f (new_AGEMA_signal_13972), .B0_t (MixColumnsIns_MixOneColumnInst_0_n138), .B0_f (new_AGEMA_signal_14474), .B1_t (new_AGEMA_signal_14475), .B1_f (new_AGEMA_signal_14476), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n139), .Z0_f (new_AGEMA_signal_15122), .Z1_t (new_AGEMA_signal_15123), .Z1_f (new_AGEMA_signal_15124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U36 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n137), .A0_f (new_AGEMA_signal_15881), .A1_t (new_AGEMA_signal_15882), .A1_f (new_AGEMA_signal_15883), .B0_t (MixColumnsIns_MixOneColumnInst_0_n154), .B0_f (new_AGEMA_signal_15125), .B1_t (new_AGEMA_signal_15126), .B1_f (new_AGEMA_signal_15127), .Z0_t (MixColumnsOutput[113]), .Z0_f (new_AGEMA_signal_16838), .Z1_t (new_AGEMA_signal_16839), .Z1_f (new_AGEMA_signal_16840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U35 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]), .A0_f (new_AGEMA_signal_14501), .A1_t (new_AGEMA_signal_14502), .A1_f (new_AGEMA_signal_14503), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13763), .B1_t (new_AGEMA_signal_13764), .B1_f (new_AGEMA_signal_13765), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n154), .Z0_f (new_AGEMA_signal_15125), .Z1_t (new_AGEMA_signal_15126), .Z1_f (new_AGEMA_signal_15127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U34 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n191), .A0_f (new_AGEMA_signal_15128), .A1_t (new_AGEMA_signal_15129), .A1_f (new_AGEMA_signal_15130), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13973), .B1_t (new_AGEMA_signal_13974), .B1_f (new_AGEMA_signal_13975), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n137), .Z0_f (new_AGEMA_signal_15881), .Z1_t (new_AGEMA_signal_15882), .Z1_f (new_AGEMA_signal_15883) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U33 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]), .A0_f (new_AGEMA_signal_14510), .A1_t (new_AGEMA_signal_14511), .A1_f (new_AGEMA_signal_14512), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .B0_f (new_AGEMA_signal_13658), .B1_t (new_AGEMA_signal_13659), .B1_f (new_AGEMA_signal_13660), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n191), .Z0_f (new_AGEMA_signal_15128), .Z1_t (new_AGEMA_signal_15129), .Z1_f (new_AGEMA_signal_15130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U32 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n136), .A0_f (new_AGEMA_signal_15131), .A1_t (new_AGEMA_signal_15132), .A1_f (new_AGEMA_signal_15133), .B0_t (MixColumnsIns_MixOneColumnInst_0_n152), .B0_f (new_AGEMA_signal_14450), .B1_t (new_AGEMA_signal_14451), .B1_f (new_AGEMA_signal_14452), .Z0_t (MixColumnsOutput[112]), .Z0_f (new_AGEMA_signal_15884), .Z1_t (new_AGEMA_signal_15885), .Z1_f (new_AGEMA_signal_15886) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U31 ( .A0_t (MixColumnsInput[104]), .A0_f (new_AGEMA_signal_13163), .A1_t (new_AGEMA_signal_13164), .A1_f (new_AGEMA_signal_13165), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13850), .B1_t (new_AGEMA_signal_13851), .B1_f (new_AGEMA_signal_13852), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n152), .Z0_f (new_AGEMA_signal_14450), .Z1_t (new_AGEMA_signal_14451), .Z1_f (new_AGEMA_signal_14452) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U30 ( .A0_t (MixColumnsInput[120]), .A0_f (new_AGEMA_signal_13493), .A1_t (new_AGEMA_signal_13494), .A1_f (new_AGEMA_signal_13495), .B0_t (MixColumnsIns_MixOneColumnInst_0_n188), .B0_f (new_AGEMA_signal_14453), .B1_t (new_AGEMA_signal_14454), .B1_f (new_AGEMA_signal_14455), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n136), .Z0_f (new_AGEMA_signal_15131), .Z1_t (new_AGEMA_signal_15132), .Z1_f (new_AGEMA_signal_15133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U29 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13745), .A1_t (new_AGEMA_signal_13746), .A1_f (new_AGEMA_signal_13747), .B0_t (MixColumnsInput[96]), .B0_f (new_AGEMA_signal_12998), .B1_t (new_AGEMA_signal_12999), .B1_f (new_AGEMA_signal_13000), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n188), .Z0_f (new_AGEMA_signal_14453), .Z1_t (new_AGEMA_signal_14454), .Z1_f (new_AGEMA_signal_14455) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U28 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n135), .A0_f (new_AGEMA_signal_15134), .A1_t (new_AGEMA_signal_15135), .A1_f (new_AGEMA_signal_15136), .B0_t (MixColumnsIns_MixOneColumnInst_0_n149), .B0_f (new_AGEMA_signal_14456), .B1_t (new_AGEMA_signal_14457), .B1_f (new_AGEMA_signal_14458), .Z0_t (MixColumnsOutput[111]), .Z0_f (new_AGEMA_signal_15887), .Z1_t (new_AGEMA_signal_15888), .Z1_f (new_AGEMA_signal_15889) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U27 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13640), .A1_t (new_AGEMA_signal_13641), .A1_f (new_AGEMA_signal_13642), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13748), .B1_t (new_AGEMA_signal_13749), .B1_f (new_AGEMA_signal_13750), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n149), .Z0_f (new_AGEMA_signal_14456), .Z1_t (new_AGEMA_signal_14457), .Z1_f (new_AGEMA_signal_14458) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U26 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n184), .A0_f (new_AGEMA_signal_14459), .A1_t (new_AGEMA_signal_14460), .A1_f (new_AGEMA_signal_14461), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13850), .B1_t (new_AGEMA_signal_13851), .B1_f (new_AGEMA_signal_13852), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n135), .Z0_f (new_AGEMA_signal_15134), .Z1_t (new_AGEMA_signal_15135), .Z1_f (new_AGEMA_signal_15136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U25 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13643), .A1_t (new_AGEMA_signal_13644), .A1_f (new_AGEMA_signal_13645), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13955), .B1_t (new_AGEMA_signal_13956), .B1_f (new_AGEMA_signal_13957), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n184), .Z0_f (new_AGEMA_signal_14459), .Z1_t (new_AGEMA_signal_14460), .Z1_f (new_AGEMA_signal_14461) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U24 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n134), .A0_f (new_AGEMA_signal_15137), .A1_t (new_AGEMA_signal_15138), .A1_f (new_AGEMA_signal_15139), .B0_t (MixColumnsIns_MixOneColumnInst_0_n147), .B0_f (new_AGEMA_signal_14462), .B1_t (new_AGEMA_signal_14463), .B1_f (new_AGEMA_signal_14464), .Z0_t (MixColumnsOutput[110]), .Z0_f (new_AGEMA_signal_15890), .Z1_t (new_AGEMA_signal_15891), .Z1_f (new_AGEMA_signal_15892) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U23 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13643), .A1_t (new_AGEMA_signal_13644), .A1_f (new_AGEMA_signal_13645), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13751), .B1_t (new_AGEMA_signal_13752), .B1_f (new_AGEMA_signal_13753), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n147), .Z0_f (new_AGEMA_signal_14462), .Z1_t (new_AGEMA_signal_14463), .Z1_f (new_AGEMA_signal_14464) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U22 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n181), .A0_f (new_AGEMA_signal_14465), .A1_t (new_AGEMA_signal_14466), .A1_f (new_AGEMA_signal_14467), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13853), .B1_t (new_AGEMA_signal_13854), .B1_f (new_AGEMA_signal_13855), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n134), .Z0_f (new_AGEMA_signal_15137), .Z1_t (new_AGEMA_signal_15138), .Z1_f (new_AGEMA_signal_15139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U21 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13646), .A1_t (new_AGEMA_signal_13647), .A1_f (new_AGEMA_signal_13648), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13958), .B1_t (new_AGEMA_signal_13959), .B1_f (new_AGEMA_signal_13960), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n181), .Z0_f (new_AGEMA_signal_14465), .Z1_t (new_AGEMA_signal_14466), .Z1_f (new_AGEMA_signal_14467) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U20 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n133), .A0_f (new_AGEMA_signal_15140), .A1_t (new_AGEMA_signal_15141), .A1_f (new_AGEMA_signal_15142), .B0_t (MixColumnsIns_MixOneColumnInst_0_n145), .B0_f (new_AGEMA_signal_14468), .B1_t (new_AGEMA_signal_14469), .B1_f (new_AGEMA_signal_14470), .Z0_t (MixColumnsOutput[109]), .Z0_f (new_AGEMA_signal_15893), .Z1_t (new_AGEMA_signal_15894), .Z1_f (new_AGEMA_signal_15895) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U19 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13646), .A1_t (new_AGEMA_signal_13647), .A1_f (new_AGEMA_signal_13648), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13754), .B1_t (new_AGEMA_signal_13755), .B1_f (new_AGEMA_signal_13756), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n145), .Z0_f (new_AGEMA_signal_14468), .Z1_t (new_AGEMA_signal_14469), .Z1_f (new_AGEMA_signal_14470) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U18 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n178), .A0_f (new_AGEMA_signal_14471), .A1_t (new_AGEMA_signal_14472), .A1_f (new_AGEMA_signal_14473), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13856), .B1_t (new_AGEMA_signal_13857), .B1_f (new_AGEMA_signal_13858), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n133), .Z0_f (new_AGEMA_signal_15140), .Z1_t (new_AGEMA_signal_15141), .Z1_f (new_AGEMA_signal_15142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U17 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13649), .A1_t (new_AGEMA_signal_13650), .A1_f (new_AGEMA_signal_13651), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13961), .B1_t (new_AGEMA_signal_13962), .B1_f (new_AGEMA_signal_13963), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n178), .Z0_f (new_AGEMA_signal_14471), .Z1_t (new_AGEMA_signal_14472), .Z1_f (new_AGEMA_signal_14473) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U16 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n132), .A0_f (new_AGEMA_signal_15896), .A1_t (new_AGEMA_signal_15897), .A1_f (new_AGEMA_signal_15898), .B0_t (MixColumnsIns_MixOneColumnInst_0_n143), .B0_f (new_AGEMA_signal_15143), .B1_t (new_AGEMA_signal_15144), .B1_f (new_AGEMA_signal_15145), .Z0_t (MixColumnsOutput[108]), .Z0_f (new_AGEMA_signal_16841), .Z1_t (new_AGEMA_signal_16842), .Z1_f (new_AGEMA_signal_16843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U15 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13649), .A1_t (new_AGEMA_signal_13650), .A1_f (new_AGEMA_signal_13651), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]), .B0_f (new_AGEMA_signal_14504), .B1_t (new_AGEMA_signal_14505), .B1_f (new_AGEMA_signal_14506), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n143), .Z0_f (new_AGEMA_signal_15143), .Z1_t (new_AGEMA_signal_15144), .Z1_f (new_AGEMA_signal_15145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U14 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n175), .A0_f (new_AGEMA_signal_15146), .A1_t (new_AGEMA_signal_15147), .A1_f (new_AGEMA_signal_15148), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13859), .B1_t (new_AGEMA_signal_13860), .B1_f (new_AGEMA_signal_13861), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n132), .Z0_f (new_AGEMA_signal_15896), .Z1_t (new_AGEMA_signal_15897), .Z1_f (new_AGEMA_signal_15898) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U13 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]), .A0_f (new_AGEMA_signal_14513), .A1_t (new_AGEMA_signal_14514), .A1_f (new_AGEMA_signal_14515), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13964), .B1_t (new_AGEMA_signal_13965), .B1_f (new_AGEMA_signal_13966), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n175), .Z0_f (new_AGEMA_signal_15146), .Z1_t (new_AGEMA_signal_15147), .Z1_f (new_AGEMA_signal_15148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U12 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n131), .A0_f (new_AGEMA_signal_15899), .A1_t (new_AGEMA_signal_15900), .A1_f (new_AGEMA_signal_15901), .B0_t (MixColumnsIns_MixOneColumnInst_0_n140), .B0_f (new_AGEMA_signal_15149), .B1_t (new_AGEMA_signal_15150), .B1_f (new_AGEMA_signal_15151), .Z0_t (MixColumnsOutput[107]), .Z0_f (new_AGEMA_signal_16844), .Z1_t (new_AGEMA_signal_16845), .Z1_f (new_AGEMA_signal_16846) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U11 ( .A0_t (MixColumnsInput[99]), .A0_f (new_AGEMA_signal_13652), .A1_t (new_AGEMA_signal_13653), .A1_f (new_AGEMA_signal_13654), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]), .B0_f (new_AGEMA_signal_14507), .B1_t (new_AGEMA_signal_14508), .B1_f (new_AGEMA_signal_14509), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n140), .Z0_f (new_AGEMA_signal_15149), .Z1_t (new_AGEMA_signal_15150), .Z1_f (new_AGEMA_signal_15151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U10 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n172), .A0_f (new_AGEMA_signal_15152), .A1_t (new_AGEMA_signal_15153), .A1_f (new_AGEMA_signal_15154), .B0_t (MixColumnsInput[115]), .B0_f (new_AGEMA_signal_13862), .B1_t (new_AGEMA_signal_13863), .B1_f (new_AGEMA_signal_13864), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n131), .Z0_f (new_AGEMA_signal_15899), .Z1_t (new_AGEMA_signal_15900), .Z1_f (new_AGEMA_signal_15901) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U9 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]), .A0_f (new_AGEMA_signal_14516), .A1_t (new_AGEMA_signal_14517), .A1_f (new_AGEMA_signal_14518), .B0_t (MixColumnsInput[123]), .B0_f (new_AGEMA_signal_13967), .B1_t (new_AGEMA_signal_13968), .B1_f (new_AGEMA_signal_13969), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n172), .Z0_f (new_AGEMA_signal_15152), .Z1_t (new_AGEMA_signal_15153), .Z1_f (new_AGEMA_signal_15154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U8 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n130), .A0_f (new_AGEMA_signal_15155), .A1_t (new_AGEMA_signal_15156), .A1_f (new_AGEMA_signal_15157), .B0_t (MixColumnsIns_MixOneColumnInst_0_n138), .B0_f (new_AGEMA_signal_14474), .B1_t (new_AGEMA_signal_14475), .B1_f (new_AGEMA_signal_14476), .Z0_t (MixColumnsOutput[106]), .Z0_f (new_AGEMA_signal_15902), .Z1_t (new_AGEMA_signal_15903), .Z1_f (new_AGEMA_signal_15904) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U7 ( .A0_t (MixColumnsInput[98]), .A0_f (new_AGEMA_signal_13655), .A1_t (new_AGEMA_signal_13656), .A1_f (new_AGEMA_signal_13657), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13763), .B1_t (new_AGEMA_signal_13764), .B1_f (new_AGEMA_signal_13765), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n138), .Z0_f (new_AGEMA_signal_14474), .Z1_t (new_AGEMA_signal_14475), .Z1_f (new_AGEMA_signal_14476) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U6 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n165), .A0_f (new_AGEMA_signal_14477), .A1_t (new_AGEMA_signal_14478), .A1_f (new_AGEMA_signal_14479), .B0_t (MixColumnsInput[114]), .B0_f (new_AGEMA_signal_13865), .B1_t (new_AGEMA_signal_13866), .B1_f (new_AGEMA_signal_13867), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n130), .Z0_f (new_AGEMA_signal_15155), .Z1_t (new_AGEMA_signal_15156), .Z1_f (new_AGEMA_signal_15157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U5 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .A0_f (new_AGEMA_signal_13658), .A1_t (new_AGEMA_signal_13659), .A1_f (new_AGEMA_signal_13660), .B0_t (MixColumnsInput[122]), .B0_f (new_AGEMA_signal_13970), .B1_t (new_AGEMA_signal_13971), .B1_f (new_AGEMA_signal_13972), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n165), .Z0_f (new_AGEMA_signal_14477), .Z1_t (new_AGEMA_signal_14478), .Z1_f (new_AGEMA_signal_14479) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n129), .A0_f (new_AGEMA_signal_15158), .A1_t (new_AGEMA_signal_15159), .A1_f (new_AGEMA_signal_15160), .B0_t (MixColumnsInput[104]), .B0_f (new_AGEMA_signal_13163), .B1_t (new_AGEMA_signal_13164), .B1_f (new_AGEMA_signal_13165), .Z0_t (MixColumnsOutput[96]), .Z0_f (new_AGEMA_signal_15905), .Z1_t (new_AGEMA_signal_15906), .Z1_f (new_AGEMA_signal_15907) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n187), .A0_f (new_AGEMA_signal_14483), .A1_t (new_AGEMA_signal_14484), .A1_f (new_AGEMA_signal_14485), .B0_t (MixColumnsIns_MixOneColumnInst_0_n151), .B0_f (new_AGEMA_signal_14480), .B1_t (new_AGEMA_signal_14481), .B1_f (new_AGEMA_signal_14482), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n129), .Z0_f (new_AGEMA_signal_15158), .Z1_t (new_AGEMA_signal_15159), .Z1_f (new_AGEMA_signal_15160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U2 ( .A0_t (MixColumnsInput[112]), .A0_f (new_AGEMA_signal_13328), .A1_t (new_AGEMA_signal_13329), .A1_f (new_AGEMA_signal_13330), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13955), .B1_t (new_AGEMA_signal_13956), .B1_f (new_AGEMA_signal_13957), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n151), .Z0_f (new_AGEMA_signal_14480), .Z1_t (new_AGEMA_signal_14481), .Z1_f (new_AGEMA_signal_14482) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U1 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13640), .A1_t (new_AGEMA_signal_13641), .A1_f (new_AGEMA_signal_13642), .B0_t (MixColumnsInput[120]), .B0_f (new_AGEMA_signal_13493), .B1_t (new_AGEMA_signal_13494), .B1_f (new_AGEMA_signal_13495), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n187), .Z0_f (new_AGEMA_signal_14483), .Z1_t (new_AGEMA_signal_14484), .Z1_f (new_AGEMA_signal_14485) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13955), .A1_t (new_AGEMA_signal_13956), .A1_f (new_AGEMA_signal_13957), .B0_t (MixColumnsInput[123]), .B0_f (new_AGEMA_signal_13967), .B1_t (new_AGEMA_signal_13968), .B1_f (new_AGEMA_signal_13969), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]), .Z0_f (new_AGEMA_signal_14486), .Z1_t (new_AGEMA_signal_14487), .Z1_f (new_AGEMA_signal_14488) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13955), .A1_t (new_AGEMA_signal_13956), .A1_f (new_AGEMA_signal_13957), .B0_t (MixColumnsInput[122]), .B0_f (new_AGEMA_signal_13970), .B1_t (new_AGEMA_signal_13971), .B1_f (new_AGEMA_signal_13972), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]), .Z0_f (new_AGEMA_signal_14489), .Z1_t (new_AGEMA_signal_14490), .Z1_f (new_AGEMA_signal_14491) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13955), .A1_t (new_AGEMA_signal_13956), .A1_f (new_AGEMA_signal_13957), .B0_t (MixColumnsInput[120]), .B0_f (new_AGEMA_signal_13493), .B1_t (new_AGEMA_signal_13494), .B1_f (new_AGEMA_signal_13495), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]), .Z0_f (new_AGEMA_signal_14492), .Z1_t (new_AGEMA_signal_14493), .Z1_f (new_AGEMA_signal_14494) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13850), .A1_t (new_AGEMA_signal_13851), .A1_f (new_AGEMA_signal_13852), .B0_t (MixColumnsInput[115]), .B0_f (new_AGEMA_signal_13862), .B1_t (new_AGEMA_signal_13863), .B1_f (new_AGEMA_signal_13864), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]), .Z0_f (new_AGEMA_signal_14495), .Z1_t (new_AGEMA_signal_14496), .Z1_f (new_AGEMA_signal_14497) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13850), .A1_t (new_AGEMA_signal_13851), .A1_f (new_AGEMA_signal_13852), .B0_t (MixColumnsInput[114]), .B0_f (new_AGEMA_signal_13865), .B1_t (new_AGEMA_signal_13866), .B1_f (new_AGEMA_signal_13867), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]), .Z0_f (new_AGEMA_signal_14498), .Z1_t (new_AGEMA_signal_14499), .Z1_f (new_AGEMA_signal_14500) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13850), .A1_t (new_AGEMA_signal_13851), .A1_f (new_AGEMA_signal_13852), .B0_t (MixColumnsInput[112]), .B0_f (new_AGEMA_signal_13328), .B1_t (new_AGEMA_signal_13329), .B1_f (new_AGEMA_signal_13330), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]), .Z0_f (new_AGEMA_signal_14501), .Z1_t (new_AGEMA_signal_14502), .Z1_f (new_AGEMA_signal_14503) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13745), .A1_t (new_AGEMA_signal_13746), .A1_f (new_AGEMA_signal_13747), .B0_t (MixColumnsInput[107]), .B0_f (new_AGEMA_signal_13757), .B1_t (new_AGEMA_signal_13758), .B1_f (new_AGEMA_signal_13759), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]), .Z0_f (new_AGEMA_signal_14504), .Z1_t (new_AGEMA_signal_14505), .Z1_f (new_AGEMA_signal_14506) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13745), .A1_t (new_AGEMA_signal_13746), .A1_f (new_AGEMA_signal_13747), .B0_t (MixColumnsInput[106]), .B0_f (new_AGEMA_signal_13760), .B1_t (new_AGEMA_signal_13761), .B1_f (new_AGEMA_signal_13762), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]), .Z0_f (new_AGEMA_signal_14507), .Z1_t (new_AGEMA_signal_14508), .Z1_f (new_AGEMA_signal_14509) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13745), .A1_t (new_AGEMA_signal_13746), .A1_f (new_AGEMA_signal_13747), .B0_t (MixColumnsInput[104]), .B0_f (new_AGEMA_signal_13163), .B1_t (new_AGEMA_signal_13164), .B1_f (new_AGEMA_signal_13165), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]), .Z0_f (new_AGEMA_signal_14510), .Z1_t (new_AGEMA_signal_14511), .Z1_f (new_AGEMA_signal_14512) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13640), .A1_t (new_AGEMA_signal_13641), .A1_f (new_AGEMA_signal_13642), .B0_t (MixColumnsInput[99]), .B0_f (new_AGEMA_signal_13652), .B1_t (new_AGEMA_signal_13653), .B1_f (new_AGEMA_signal_13654), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]), .Z0_f (new_AGEMA_signal_14513), .Z1_t (new_AGEMA_signal_14514), .Z1_f (new_AGEMA_signal_14515) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13640), .A1_t (new_AGEMA_signal_13641), .A1_f (new_AGEMA_signal_13642), .B0_t (MixColumnsInput[98]), .B0_f (new_AGEMA_signal_13655), .B1_t (new_AGEMA_signal_13656), .B1_f (new_AGEMA_signal_13657), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]), .Z0_f (new_AGEMA_signal_14516), .Z1_t (new_AGEMA_signal_14517), .Z1_f (new_AGEMA_signal_14518) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13640), .A1_t (new_AGEMA_signal_13641), .A1_f (new_AGEMA_signal_13642), .B0_t (MixColumnsInput[96]), .B0_f (new_AGEMA_signal_12998), .B1_t (new_AGEMA_signal_12999), .B1_f (new_AGEMA_signal_13000), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]), .Z0_f (new_AGEMA_signal_14519), .Z1_t (new_AGEMA_signal_14520), .Z1_f (new_AGEMA_signal_14521) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U96 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n192), .A0_f (new_AGEMA_signal_15908), .A1_t (new_AGEMA_signal_15909), .A1_f (new_AGEMA_signal_15910), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13784), .B1_t (new_AGEMA_signal_13785), .B1_f (new_AGEMA_signal_13786), .Z0_t (MixColumnsOutput[73]), .Z0_f (new_AGEMA_signal_16847), .Z1_t (new_AGEMA_signal_16848), .Z1_f (new_AGEMA_signal_16849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U95 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n191), .A0_f (new_AGEMA_signal_15224), .A1_t (new_AGEMA_signal_15225), .A1_f (new_AGEMA_signal_15226), .B0_t (MixColumnsIns_MixOneColumnInst_1_n190), .B0_f (new_AGEMA_signal_15212), .B1_t (new_AGEMA_signal_15213), .B1_f (new_AGEMA_signal_15214), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n192), .Z0_f (new_AGEMA_signal_15908), .Z1_t (new_AGEMA_signal_15909), .Z1_f (new_AGEMA_signal_15910) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U94 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n189), .A0_f (new_AGEMA_signal_15161), .A1_t (new_AGEMA_signal_15162), .A1_f (new_AGEMA_signal_15163), .B0_t (MixColumnsIns_MixOneColumnInst_1_n188), .B0_f (new_AGEMA_signal_14549), .B1_t (new_AGEMA_signal_14550), .B1_f (new_AGEMA_signal_14551), .Z0_t (MixColumnsOutput[72]), .Z0_f (new_AGEMA_signal_15911), .Z1_t (new_AGEMA_signal_15912), .Z1_f (new_AGEMA_signal_15913) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U93 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n187), .A0_f (new_AGEMA_signal_14579), .A1_t (new_AGEMA_signal_14580), .A1_f (new_AGEMA_signal_14581), .B0_t (MixColumnsInput[80]), .B0_f (new_AGEMA_signal_13196), .B1_t (new_AGEMA_signal_13197), .B1_f (new_AGEMA_signal_13198), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n189), .Z0_f (new_AGEMA_signal_15161), .Z1_t (new_AGEMA_signal_15162), .Z1_f (new_AGEMA_signal_15163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U92 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n186), .A0_f (new_AGEMA_signal_15164), .A1_t (new_AGEMA_signal_15165), .A1_f (new_AGEMA_signal_15166), .B0_t (MixColumnsIns_MixOneColumnInst_1_n185), .B0_f (new_AGEMA_signal_14522), .B1_t (new_AGEMA_signal_14523), .B1_f (new_AGEMA_signal_14524), .Z0_t (MixColumnsOutput[71]), .Z0_f (new_AGEMA_signal_15914), .Z1_t (new_AGEMA_signal_15915), .Z1_f (new_AGEMA_signal_15916) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U91 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n184), .A0_f (new_AGEMA_signal_14555), .A1_t (new_AGEMA_signal_14556), .A1_f (new_AGEMA_signal_14557), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B0_f (new_AGEMA_signal_13661), .B1_t (new_AGEMA_signal_13662), .B1_f (new_AGEMA_signal_13663), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n186), .Z0_f (new_AGEMA_signal_15164), .Z1_t (new_AGEMA_signal_15165), .Z1_f (new_AGEMA_signal_15166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U90 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n183), .A0_f (new_AGEMA_signal_15167), .A1_t (new_AGEMA_signal_15168), .A1_f (new_AGEMA_signal_15169), .B0_t (MixColumnsIns_MixOneColumnInst_1_n182), .B0_f (new_AGEMA_signal_14525), .B1_t (new_AGEMA_signal_14526), .B1_f (new_AGEMA_signal_14527), .Z0_t (MixColumnsOutput[70]), .Z0_f (new_AGEMA_signal_15917), .Z1_t (new_AGEMA_signal_15918), .Z1_f (new_AGEMA_signal_15919) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U89 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n181), .A0_f (new_AGEMA_signal_14561), .A1_t (new_AGEMA_signal_14562), .A1_f (new_AGEMA_signal_14563), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13664), .B1_t (new_AGEMA_signal_13665), .B1_f (new_AGEMA_signal_13666), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n183), .Z0_f (new_AGEMA_signal_15167), .Z1_t (new_AGEMA_signal_15168), .Z1_f (new_AGEMA_signal_15169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U88 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n180), .A0_f (new_AGEMA_signal_15170), .A1_t (new_AGEMA_signal_15171), .A1_f (new_AGEMA_signal_15172), .B0_t (MixColumnsIns_MixOneColumnInst_1_n179), .B0_f (new_AGEMA_signal_14528), .B1_t (new_AGEMA_signal_14529), .B1_f (new_AGEMA_signal_14530), .Z0_t (MixColumnsOutput[69]), .Z0_f (new_AGEMA_signal_15920), .Z1_t (new_AGEMA_signal_15921), .Z1_f (new_AGEMA_signal_15922) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U87 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n178), .A0_f (new_AGEMA_signal_14567), .A1_t (new_AGEMA_signal_14568), .A1_f (new_AGEMA_signal_14569), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13667), .B1_t (new_AGEMA_signal_13668), .B1_f (new_AGEMA_signal_13669), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n180), .Z0_f (new_AGEMA_signal_15170), .Z1_t (new_AGEMA_signal_15171), .Z1_f (new_AGEMA_signal_15172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U86 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n177), .A0_f (new_AGEMA_signal_15923), .A1_t (new_AGEMA_signal_15924), .A1_f (new_AGEMA_signal_15925), .B0_t (MixColumnsIns_MixOneColumnInst_1_n176), .B0_f (new_AGEMA_signal_15185), .B1_t (new_AGEMA_signal_15186), .B1_f (new_AGEMA_signal_15187), .Z0_t (MixColumnsOutput[68]), .Z0_f (new_AGEMA_signal_16850), .Z1_t (new_AGEMA_signal_16851), .Z1_f (new_AGEMA_signal_16852) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U85 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n175), .A0_f (new_AGEMA_signal_15242), .A1_t (new_AGEMA_signal_15243), .A1_f (new_AGEMA_signal_15244), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13670), .B1_t (new_AGEMA_signal_13671), .B1_f (new_AGEMA_signal_13672), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n177), .Z0_f (new_AGEMA_signal_15923), .Z1_t (new_AGEMA_signal_15924), .Z1_f (new_AGEMA_signal_15925) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U84 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n174), .A0_f (new_AGEMA_signal_15926), .A1_t (new_AGEMA_signal_15927), .A1_f (new_AGEMA_signal_15928), .B0_t (MixColumnsIns_MixOneColumnInst_1_n173), .B0_f (new_AGEMA_signal_15188), .B1_t (new_AGEMA_signal_15189), .B1_f (new_AGEMA_signal_15190), .Z0_t (MixColumnsOutput[67]), .Z0_f (new_AGEMA_signal_16853), .Z1_t (new_AGEMA_signal_16854), .Z1_f (new_AGEMA_signal_16855) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U83 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n172), .A0_f (new_AGEMA_signal_15248), .A1_t (new_AGEMA_signal_15249), .A1_f (new_AGEMA_signal_15250), .B0_t (MixColumnsInput[75]), .B0_f (new_AGEMA_signal_13673), .B1_t (new_AGEMA_signal_13674), .B1_f (new_AGEMA_signal_13675), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n174), .Z0_f (new_AGEMA_signal_15926), .Z1_t (new_AGEMA_signal_15927), .Z1_f (new_AGEMA_signal_15928) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U82 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n171), .A0_f (new_AGEMA_signal_15173), .A1_t (new_AGEMA_signal_15174), .A1_f (new_AGEMA_signal_15175), .B0_t (MixColumnsIns_MixOneColumnInst_1_n185), .B0_f (new_AGEMA_signal_14522), .B1_t (new_AGEMA_signal_14523), .B1_f (new_AGEMA_signal_14524), .Z0_t (MixColumnsOutput[95]), .Z0_f (new_AGEMA_signal_15929), .Z1_t (new_AGEMA_signal_15930), .Z1_f (new_AGEMA_signal_15931) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U81 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13766), .A1_t (new_AGEMA_signal_13767), .A1_f (new_AGEMA_signal_13768), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13874), .B1_t (new_AGEMA_signal_13875), .B1_f (new_AGEMA_signal_13876), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n185), .Z0_f (new_AGEMA_signal_14522), .Z1_t (new_AGEMA_signal_14523), .Z1_f (new_AGEMA_signal_14524) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U80 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13892), .A1_t (new_AGEMA_signal_13893), .A1_f (new_AGEMA_signal_13894), .B0_t (MixColumnsIns_MixOneColumnInst_1_n170), .B0_f (new_AGEMA_signal_14534), .B1_t (new_AGEMA_signal_14535), .B1_f (new_AGEMA_signal_14536), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n171), .Z0_f (new_AGEMA_signal_15173), .Z1_t (new_AGEMA_signal_15174), .Z1_f (new_AGEMA_signal_15175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U79 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n169), .A0_f (new_AGEMA_signal_15176), .A1_t (new_AGEMA_signal_15177), .A1_f (new_AGEMA_signal_15178), .B0_t (MixColumnsIns_MixOneColumnInst_1_n182), .B0_f (new_AGEMA_signal_14525), .B1_t (new_AGEMA_signal_14526), .B1_f (new_AGEMA_signal_14527), .Z0_t (MixColumnsOutput[94]), .Z0_f (new_AGEMA_signal_15932), .Z1_t (new_AGEMA_signal_15933), .Z1_f (new_AGEMA_signal_15934) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U78 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .A0_f (new_AGEMA_signal_13769), .A1_t (new_AGEMA_signal_13770), .A1_f (new_AGEMA_signal_13771), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13877), .B1_t (new_AGEMA_signal_13878), .B1_f (new_AGEMA_signal_13879), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n182), .Z0_f (new_AGEMA_signal_14525), .Z1_t (new_AGEMA_signal_14526), .Z1_f (new_AGEMA_signal_14527) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U77 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13895), .A1_t (new_AGEMA_signal_13896), .A1_f (new_AGEMA_signal_13897), .B0_t (MixColumnsIns_MixOneColumnInst_1_n168), .B0_f (new_AGEMA_signal_14537), .B1_t (new_AGEMA_signal_14538), .B1_f (new_AGEMA_signal_14539), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n169), .Z0_f (new_AGEMA_signal_15176), .Z1_t (new_AGEMA_signal_15177), .Z1_f (new_AGEMA_signal_15178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U76 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n167), .A0_f (new_AGEMA_signal_15179), .A1_t (new_AGEMA_signal_15180), .A1_f (new_AGEMA_signal_15181), .B0_t (MixColumnsIns_MixOneColumnInst_1_n166), .B0_f (new_AGEMA_signal_14531), .B1_t (new_AGEMA_signal_14532), .B1_f (new_AGEMA_signal_14533), .Z0_t (MixColumnsOutput[66]), .Z0_f (new_AGEMA_signal_15935), .Z1_t (new_AGEMA_signal_15936), .Z1_f (new_AGEMA_signal_15937) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U75 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n165), .A0_f (new_AGEMA_signal_14573), .A1_t (new_AGEMA_signal_14574), .A1_f (new_AGEMA_signal_14575), .B0_t (MixColumnsInput[74]), .B0_f (new_AGEMA_signal_13676), .B1_t (new_AGEMA_signal_13677), .B1_f (new_AGEMA_signal_13678), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n167), .Z0_f (new_AGEMA_signal_15179), .Z1_t (new_AGEMA_signal_15180), .Z1_f (new_AGEMA_signal_15181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U74 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n164), .A0_f (new_AGEMA_signal_15182), .A1_t (new_AGEMA_signal_15183), .A1_f (new_AGEMA_signal_15184), .B0_t (MixColumnsIns_MixOneColumnInst_1_n179), .B0_f (new_AGEMA_signal_14528), .B1_t (new_AGEMA_signal_14529), .B1_f (new_AGEMA_signal_14530), .Z0_t (MixColumnsOutput[93]), .Z0_f (new_AGEMA_signal_15938), .Z1_t (new_AGEMA_signal_15939), .Z1_f (new_AGEMA_signal_15940) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U73 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .A0_f (new_AGEMA_signal_13772), .A1_t (new_AGEMA_signal_13773), .A1_f (new_AGEMA_signal_13774), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13880), .B1_t (new_AGEMA_signal_13881), .B1_f (new_AGEMA_signal_13882), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n179), .Z0_f (new_AGEMA_signal_14528), .Z1_t (new_AGEMA_signal_14529), .Z1_f (new_AGEMA_signal_14530) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U72 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13898), .A1_t (new_AGEMA_signal_13899), .A1_f (new_AGEMA_signal_13900), .B0_t (MixColumnsIns_MixOneColumnInst_1_n163), .B0_f (new_AGEMA_signal_14540), .B1_t (new_AGEMA_signal_14541), .B1_f (new_AGEMA_signal_14542), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n164), .Z0_f (new_AGEMA_signal_15182), .Z1_t (new_AGEMA_signal_15183), .Z1_f (new_AGEMA_signal_15184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U71 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n162), .A0_f (new_AGEMA_signal_15941), .A1_t (new_AGEMA_signal_15942), .A1_f (new_AGEMA_signal_15943), .B0_t (MixColumnsIns_MixOneColumnInst_1_n176), .B0_f (new_AGEMA_signal_15185), .B1_t (new_AGEMA_signal_15186), .B1_f (new_AGEMA_signal_15187), .Z0_t (MixColumnsOutput[92]), .Z0_f (new_AGEMA_signal_16856), .Z1_t (new_AGEMA_signal_16857), .Z1_f (new_AGEMA_signal_16858) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U70 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .A0_f (new_AGEMA_signal_13775), .A1_t (new_AGEMA_signal_13776), .A1_f (new_AGEMA_signal_13777), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]), .B0_f (new_AGEMA_signal_14582), .B1_t (new_AGEMA_signal_14583), .B1_f (new_AGEMA_signal_14584), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n176), .Z0_f (new_AGEMA_signal_15185), .Z1_t (new_AGEMA_signal_15186), .Z1_f (new_AGEMA_signal_15187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U69 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13901), .A1_t (new_AGEMA_signal_13902), .A1_f (new_AGEMA_signal_13903), .B0_t (MixColumnsIns_MixOneColumnInst_1_n161), .B0_f (new_AGEMA_signal_15206), .B1_t (new_AGEMA_signal_15207), .B1_f (new_AGEMA_signal_15208), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n162), .Z0_f (new_AGEMA_signal_15941), .Z1_t (new_AGEMA_signal_15942), .Z1_f (new_AGEMA_signal_15943) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U68 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n160), .A0_f (new_AGEMA_signal_15944), .A1_t (new_AGEMA_signal_15945), .A1_f (new_AGEMA_signal_15946), .B0_t (MixColumnsIns_MixOneColumnInst_1_n173), .B0_f (new_AGEMA_signal_15188), .B1_t (new_AGEMA_signal_15189), .B1_f (new_AGEMA_signal_15190), .Z0_t (MixColumnsOutput[91]), .Z0_f (new_AGEMA_signal_16859), .Z1_t (new_AGEMA_signal_16860), .Z1_f (new_AGEMA_signal_16861) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U67 ( .A0_t (MixColumnsInput[83]), .A0_f (new_AGEMA_signal_13778), .A1_t (new_AGEMA_signal_13779), .A1_f (new_AGEMA_signal_13780), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]), .B0_f (new_AGEMA_signal_14585), .B1_t (new_AGEMA_signal_14586), .B1_f (new_AGEMA_signal_14587), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n173), .Z0_f (new_AGEMA_signal_15188), .Z1_t (new_AGEMA_signal_15189), .Z1_f (new_AGEMA_signal_15190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U66 ( .A0_t (MixColumnsInput[67]), .A0_f (new_AGEMA_signal_13904), .A1_t (new_AGEMA_signal_13905), .A1_f (new_AGEMA_signal_13906), .B0_t (MixColumnsIns_MixOneColumnInst_1_n159), .B0_f (new_AGEMA_signal_15215), .B1_t (new_AGEMA_signal_15216), .B1_f (new_AGEMA_signal_15217), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n160), .Z0_f (new_AGEMA_signal_15944), .Z1_t (new_AGEMA_signal_15945), .Z1_f (new_AGEMA_signal_15946) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U65 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n158), .A0_f (new_AGEMA_signal_15191), .A1_t (new_AGEMA_signal_15192), .A1_f (new_AGEMA_signal_15193), .B0_t (MixColumnsIns_MixOneColumnInst_1_n166), .B0_f (new_AGEMA_signal_14531), .B1_t (new_AGEMA_signal_14532), .B1_f (new_AGEMA_signal_14533), .Z0_t (MixColumnsOutput[90]), .Z0_f (new_AGEMA_signal_15947), .Z1_t (new_AGEMA_signal_15948), .Z1_f (new_AGEMA_signal_15949) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U64 ( .A0_t (MixColumnsInput[82]), .A0_f (new_AGEMA_signal_13781), .A1_t (new_AGEMA_signal_13782), .A1_f (new_AGEMA_signal_13783), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13889), .B1_t (new_AGEMA_signal_13890), .B1_f (new_AGEMA_signal_13891), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n166), .Z0_f (new_AGEMA_signal_14531), .Z1_t (new_AGEMA_signal_14532), .Z1_f (new_AGEMA_signal_14533) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U63 ( .A0_t (MixColumnsInput[66]), .A0_f (new_AGEMA_signal_13907), .A1_t (new_AGEMA_signal_13908), .A1_f (new_AGEMA_signal_13909), .B0_t (MixColumnsIns_MixOneColumnInst_1_n157), .B0_f (new_AGEMA_signal_14543), .B1_t (new_AGEMA_signal_14544), .B1_f (new_AGEMA_signal_14545), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n158), .Z0_f (new_AGEMA_signal_15191), .Z1_t (new_AGEMA_signal_15192), .Z1_f (new_AGEMA_signal_15193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U62 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n156), .A0_f (new_AGEMA_signal_15950), .A1_t (new_AGEMA_signal_15951), .A1_f (new_AGEMA_signal_15952), .B0_t (MixColumnsIns_MixOneColumnInst_1_n155), .B0_f (new_AGEMA_signal_15209), .B1_t (new_AGEMA_signal_15210), .B1_f (new_AGEMA_signal_15211), .Z0_t (MixColumnsOutput[89]), .Z0_f (new_AGEMA_signal_16862), .Z1_t (new_AGEMA_signal_16863), .Z1_f (new_AGEMA_signal_16864) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U61 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .A0_f (new_AGEMA_signal_13910), .A1_t (new_AGEMA_signal_13911), .A1_f (new_AGEMA_signal_13912), .B0_t (MixColumnsIns_MixOneColumnInst_1_n154), .B0_f (new_AGEMA_signal_15221), .B1_t (new_AGEMA_signal_15222), .B1_f (new_AGEMA_signal_15223), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n156), .Z0_f (new_AGEMA_signal_15950), .Z1_t (new_AGEMA_signal_15951), .Z1_f (new_AGEMA_signal_15952) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U60 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n153), .A0_f (new_AGEMA_signal_15194), .A1_t (new_AGEMA_signal_15195), .A1_f (new_AGEMA_signal_15196), .B0_t (MixColumnsIns_MixOneColumnInst_1_n152), .B0_f (new_AGEMA_signal_14546), .B1_t (new_AGEMA_signal_14547), .B1_f (new_AGEMA_signal_14548), .Z0_t (MixColumnsOutput[88]), .Z0_f (new_AGEMA_signal_15953), .Z1_t (new_AGEMA_signal_15954), .Z1_f (new_AGEMA_signal_15955) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U59 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n151), .A0_f (new_AGEMA_signal_14576), .A1_t (new_AGEMA_signal_14577), .A1_f (new_AGEMA_signal_14578), .B0_t (MixColumnsInput[64]), .B0_f (new_AGEMA_signal_13394), .B1_t (new_AGEMA_signal_13395), .B1_f (new_AGEMA_signal_13396), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n153), .Z0_f (new_AGEMA_signal_15194), .Z1_t (new_AGEMA_signal_15195), .Z1_f (new_AGEMA_signal_15196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U58 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n150), .A0_f (new_AGEMA_signal_15197), .A1_t (new_AGEMA_signal_15198), .A1_f (new_AGEMA_signal_15199), .B0_t (MixColumnsIns_MixOneColumnInst_1_n170), .B0_f (new_AGEMA_signal_14534), .B1_t (new_AGEMA_signal_14535), .B1_f (new_AGEMA_signal_14536), .Z0_t (MixColumnsOutput[87]), .Z0_f (new_AGEMA_signal_15956), .Z1_t (new_AGEMA_signal_15957), .Z1_f (new_AGEMA_signal_15958) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U57 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13661), .A1_t (new_AGEMA_signal_13662), .A1_f (new_AGEMA_signal_13663), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13769), .B1_t (new_AGEMA_signal_13770), .B1_f (new_AGEMA_signal_13771), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n170), .Z0_f (new_AGEMA_signal_14534), .Z1_t (new_AGEMA_signal_14535), .Z1_f (new_AGEMA_signal_14536) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U56 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13871), .A1_t (new_AGEMA_signal_13872), .A1_f (new_AGEMA_signal_13873), .B0_t (MixColumnsIns_MixOneColumnInst_1_n149), .B0_f (new_AGEMA_signal_14552), .B1_t (new_AGEMA_signal_14553), .B1_f (new_AGEMA_signal_14554), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n150), .Z0_f (new_AGEMA_signal_15197), .Z1_t (new_AGEMA_signal_15198), .Z1_f (new_AGEMA_signal_15199) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U55 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n148), .A0_f (new_AGEMA_signal_15200), .A1_t (new_AGEMA_signal_15201), .A1_f (new_AGEMA_signal_15202), .B0_t (MixColumnsIns_MixOneColumnInst_1_n168), .B0_f (new_AGEMA_signal_14537), .B1_t (new_AGEMA_signal_14538), .B1_f (new_AGEMA_signal_14539), .Z0_t (MixColumnsOutput[86]), .Z0_f (new_AGEMA_signal_15959), .Z1_t (new_AGEMA_signal_15960), .Z1_f (new_AGEMA_signal_15961) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U54 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .A0_f (new_AGEMA_signal_13664), .A1_t (new_AGEMA_signal_13665), .A1_f (new_AGEMA_signal_13666), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13772), .B1_t (new_AGEMA_signal_13773), .B1_f (new_AGEMA_signal_13774), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n168), .Z0_f (new_AGEMA_signal_14537), .Z1_t (new_AGEMA_signal_14538), .Z1_f (new_AGEMA_signal_14539) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U53 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .A0_f (new_AGEMA_signal_13874), .A1_t (new_AGEMA_signal_13875), .A1_f (new_AGEMA_signal_13876), .B0_t (MixColumnsIns_MixOneColumnInst_1_n147), .B0_f (new_AGEMA_signal_14558), .B1_t (new_AGEMA_signal_14559), .B1_f (new_AGEMA_signal_14560), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n148), .Z0_f (new_AGEMA_signal_15200), .Z1_t (new_AGEMA_signal_15201), .Z1_f (new_AGEMA_signal_15202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U52 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n146), .A0_f (new_AGEMA_signal_15203), .A1_t (new_AGEMA_signal_15204), .A1_f (new_AGEMA_signal_15205), .B0_t (MixColumnsIns_MixOneColumnInst_1_n163), .B0_f (new_AGEMA_signal_14540), .B1_t (new_AGEMA_signal_14541), .B1_f (new_AGEMA_signal_14542), .Z0_t (MixColumnsOutput[85]), .Z0_f (new_AGEMA_signal_15962), .Z1_t (new_AGEMA_signal_15963), .Z1_f (new_AGEMA_signal_15964) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U51 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .A0_f (new_AGEMA_signal_13667), .A1_t (new_AGEMA_signal_13668), .A1_f (new_AGEMA_signal_13669), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13775), .B1_t (new_AGEMA_signal_13776), .B1_f (new_AGEMA_signal_13777), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n163), .Z0_f (new_AGEMA_signal_14540), .Z1_t (new_AGEMA_signal_14541), .Z1_f (new_AGEMA_signal_14542) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U50 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .A0_f (new_AGEMA_signal_13877), .A1_t (new_AGEMA_signal_13878), .A1_f (new_AGEMA_signal_13879), .B0_t (MixColumnsIns_MixOneColumnInst_1_n145), .B0_f (new_AGEMA_signal_14564), .B1_t (new_AGEMA_signal_14565), .B1_f (new_AGEMA_signal_14566), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n146), .Z0_f (new_AGEMA_signal_15203), .Z1_t (new_AGEMA_signal_15204), .Z1_f (new_AGEMA_signal_15205) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U49 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n144), .A0_f (new_AGEMA_signal_15965), .A1_t (new_AGEMA_signal_15966), .A1_f (new_AGEMA_signal_15967), .B0_t (MixColumnsIns_MixOneColumnInst_1_n161), .B0_f (new_AGEMA_signal_15206), .B1_t (new_AGEMA_signal_15207), .B1_f (new_AGEMA_signal_15208), .Z0_t (MixColumnsOutput[84]), .Z0_f (new_AGEMA_signal_16865), .Z1_t (new_AGEMA_signal_16866), .Z1_f (new_AGEMA_signal_16867) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U48 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .A0_f (new_AGEMA_signal_13670), .A1_t (new_AGEMA_signal_13671), .A1_f (new_AGEMA_signal_13672), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]), .B0_f (new_AGEMA_signal_14591), .B1_t (new_AGEMA_signal_14592), .B1_f (new_AGEMA_signal_14593), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n161), .Z0_f (new_AGEMA_signal_15206), .Z1_t (new_AGEMA_signal_15207), .Z1_f (new_AGEMA_signal_15208) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U47 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .A0_f (new_AGEMA_signal_13880), .A1_t (new_AGEMA_signal_13881), .A1_f (new_AGEMA_signal_13882), .B0_t (MixColumnsIns_MixOneColumnInst_1_n143), .B0_f (new_AGEMA_signal_15239), .B1_t (new_AGEMA_signal_15240), .B1_f (new_AGEMA_signal_15241), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n144), .Z0_f (new_AGEMA_signal_15965), .Z1_t (new_AGEMA_signal_15966), .Z1_f (new_AGEMA_signal_15967) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U46 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n142), .A0_f (new_AGEMA_signal_15968), .A1_t (new_AGEMA_signal_15969), .A1_f (new_AGEMA_signal_15970), .B0_t (MixColumnsIns_MixOneColumnInst_1_n155), .B0_f (new_AGEMA_signal_15209), .B1_t (new_AGEMA_signal_15210), .B1_f (new_AGEMA_signal_15211), .Z0_t (MixColumnsOutput[65]), .Z0_f (new_AGEMA_signal_16868), .Z1_t (new_AGEMA_signal_16869), .Z1_f (new_AGEMA_signal_16870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U45 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .A0_f (new_AGEMA_signal_13784), .A1_t (new_AGEMA_signal_13785), .A1_f (new_AGEMA_signal_13786), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]), .B0_f (new_AGEMA_signal_14588), .B1_t (new_AGEMA_signal_14589), .B1_f (new_AGEMA_signal_14590), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n155), .Z0_f (new_AGEMA_signal_15209), .Z1_t (new_AGEMA_signal_15210), .Z1_f (new_AGEMA_signal_15211) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U44 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .A0_f (new_AGEMA_signal_13679), .A1_t (new_AGEMA_signal_13680), .A1_f (new_AGEMA_signal_13681), .B0_t (MixColumnsIns_MixOneColumnInst_1_n190), .B0_f (new_AGEMA_signal_15212), .B1_t (new_AGEMA_signal_15213), .B1_f (new_AGEMA_signal_15214), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n142), .Z0_f (new_AGEMA_signal_15968), .Z1_t (new_AGEMA_signal_15969), .Z1_f (new_AGEMA_signal_15970) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U43 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .A0_f (new_AGEMA_signal_13889), .A1_t (new_AGEMA_signal_13890), .A1_f (new_AGEMA_signal_13891), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]), .B0_f (new_AGEMA_signal_14615), .B1_t (new_AGEMA_signal_14616), .B1_f (new_AGEMA_signal_14617), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n190), .Z0_f (new_AGEMA_signal_15212), .Z1_t (new_AGEMA_signal_15213), .Z1_f (new_AGEMA_signal_15214) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U42 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n141), .A0_f (new_AGEMA_signal_15971), .A1_t (new_AGEMA_signal_15972), .A1_f (new_AGEMA_signal_15973), .B0_t (MixColumnsIns_MixOneColumnInst_1_n159), .B0_f (new_AGEMA_signal_15215), .B1_t (new_AGEMA_signal_15216), .B1_f (new_AGEMA_signal_15217), .Z0_t (MixColumnsOutput[83]), .Z0_f (new_AGEMA_signal_16871), .Z1_t (new_AGEMA_signal_16872), .Z1_f (new_AGEMA_signal_16873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U41 ( .A0_t (MixColumnsInput[75]), .A0_f (new_AGEMA_signal_13673), .A1_t (new_AGEMA_signal_13674), .A1_f (new_AGEMA_signal_13675), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]), .B0_f (new_AGEMA_signal_14594), .B1_t (new_AGEMA_signal_14595), .B1_f (new_AGEMA_signal_14596), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n159), .Z0_f (new_AGEMA_signal_15215), .Z1_t (new_AGEMA_signal_15216), .Z1_f (new_AGEMA_signal_15217) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U40 ( .A0_t (MixColumnsInput[91]), .A0_f (new_AGEMA_signal_13883), .A1_t (new_AGEMA_signal_13884), .A1_f (new_AGEMA_signal_13885), .B0_t (MixColumnsIns_MixOneColumnInst_1_n140), .B0_f (new_AGEMA_signal_15245), .B1_t (new_AGEMA_signal_15246), .B1_f (new_AGEMA_signal_15247), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n141), .Z0_f (new_AGEMA_signal_15971), .Z1_t (new_AGEMA_signal_15972), .Z1_f (new_AGEMA_signal_15973) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U39 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n139), .A0_f (new_AGEMA_signal_15218), .A1_t (new_AGEMA_signal_15219), .A1_f (new_AGEMA_signal_15220), .B0_t (MixColumnsIns_MixOneColumnInst_1_n157), .B0_f (new_AGEMA_signal_14543), .B1_t (new_AGEMA_signal_14544), .B1_f (new_AGEMA_signal_14545), .Z0_t (MixColumnsOutput[82]), .Z0_f (new_AGEMA_signal_15974), .Z1_t (new_AGEMA_signal_15975), .Z1_f (new_AGEMA_signal_15976) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U38 ( .A0_t (MixColumnsInput[74]), .A0_f (new_AGEMA_signal_13676), .A1_t (new_AGEMA_signal_13677), .A1_f (new_AGEMA_signal_13678), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13784), .B1_t (new_AGEMA_signal_13785), .B1_f (new_AGEMA_signal_13786), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n157), .Z0_f (new_AGEMA_signal_14543), .Z1_t (new_AGEMA_signal_14544), .Z1_f (new_AGEMA_signal_14545) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U37 ( .A0_t (MixColumnsInput[90]), .A0_f (new_AGEMA_signal_13886), .A1_t (new_AGEMA_signal_13887), .A1_f (new_AGEMA_signal_13888), .B0_t (MixColumnsIns_MixOneColumnInst_1_n138), .B0_f (new_AGEMA_signal_14570), .B1_t (new_AGEMA_signal_14571), .B1_f (new_AGEMA_signal_14572), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n139), .Z0_f (new_AGEMA_signal_15218), .Z1_t (new_AGEMA_signal_15219), .Z1_f (new_AGEMA_signal_15220) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U36 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n137), .A0_f (new_AGEMA_signal_15977), .A1_t (new_AGEMA_signal_15978), .A1_f (new_AGEMA_signal_15979), .B0_t (MixColumnsIns_MixOneColumnInst_1_n154), .B0_f (new_AGEMA_signal_15221), .B1_t (new_AGEMA_signal_15222), .B1_f (new_AGEMA_signal_15223), .Z0_t (MixColumnsOutput[81]), .Z0_f (new_AGEMA_signal_16874), .Z1_t (new_AGEMA_signal_16875), .Z1_f (new_AGEMA_signal_16876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U35 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]), .A0_f (new_AGEMA_signal_14597), .A1_t (new_AGEMA_signal_14598), .A1_f (new_AGEMA_signal_14599), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13679), .B1_t (new_AGEMA_signal_13680), .B1_f (new_AGEMA_signal_13681), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n154), .Z0_f (new_AGEMA_signal_15221), .Z1_t (new_AGEMA_signal_15222), .Z1_f (new_AGEMA_signal_15223) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U34 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n191), .A0_f (new_AGEMA_signal_15224), .A1_t (new_AGEMA_signal_15225), .A1_f (new_AGEMA_signal_15226), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13889), .B1_t (new_AGEMA_signal_13890), .B1_f (new_AGEMA_signal_13891), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n137), .Z0_f (new_AGEMA_signal_15977), .Z1_t (new_AGEMA_signal_15978), .Z1_f (new_AGEMA_signal_15979) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U33 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]), .A0_f (new_AGEMA_signal_14606), .A1_t (new_AGEMA_signal_14607), .A1_f (new_AGEMA_signal_14608), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .B0_f (new_AGEMA_signal_13910), .B1_t (new_AGEMA_signal_13911), .B1_f (new_AGEMA_signal_13912), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n191), .Z0_f (new_AGEMA_signal_15224), .Z1_t (new_AGEMA_signal_15225), .Z1_f (new_AGEMA_signal_15226) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U32 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n136), .A0_f (new_AGEMA_signal_15227), .A1_t (new_AGEMA_signal_15228), .A1_f (new_AGEMA_signal_15229), .B0_t (MixColumnsIns_MixOneColumnInst_1_n152), .B0_f (new_AGEMA_signal_14546), .B1_t (new_AGEMA_signal_14547), .B1_f (new_AGEMA_signal_14548), .Z0_t (MixColumnsOutput[80]), .Z0_f (new_AGEMA_signal_15980), .Z1_t (new_AGEMA_signal_15981), .Z1_f (new_AGEMA_signal_15982) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U31 ( .A0_t (MixColumnsInput[72]), .A0_f (new_AGEMA_signal_13031), .A1_t (new_AGEMA_signal_13032), .A1_f (new_AGEMA_signal_13033), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13766), .B1_t (new_AGEMA_signal_13767), .B1_f (new_AGEMA_signal_13768), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n152), .Z0_f (new_AGEMA_signal_14546), .Z1_t (new_AGEMA_signal_14547), .Z1_f (new_AGEMA_signal_14548) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U30 ( .A0_t (MixColumnsInput[88]), .A0_f (new_AGEMA_signal_13361), .A1_t (new_AGEMA_signal_13362), .A1_f (new_AGEMA_signal_13363), .B0_t (MixColumnsIns_MixOneColumnInst_1_n188), .B0_f (new_AGEMA_signal_14549), .B1_t (new_AGEMA_signal_14550), .B1_f (new_AGEMA_signal_14551), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n136), .Z0_f (new_AGEMA_signal_15227), .Z1_t (new_AGEMA_signal_15228), .Z1_f (new_AGEMA_signal_15229) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U29 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13661), .A1_t (new_AGEMA_signal_13662), .A1_f (new_AGEMA_signal_13663), .B0_t (MixColumnsInput[64]), .B0_f (new_AGEMA_signal_13394), .B1_t (new_AGEMA_signal_13395), .B1_f (new_AGEMA_signal_13396), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n188), .Z0_f (new_AGEMA_signal_14549), .Z1_t (new_AGEMA_signal_14550), .Z1_f (new_AGEMA_signal_14551) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U28 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n135), .A0_f (new_AGEMA_signal_15230), .A1_t (new_AGEMA_signal_15231), .A1_f (new_AGEMA_signal_15232), .B0_t (MixColumnsIns_MixOneColumnInst_1_n149), .B0_f (new_AGEMA_signal_14552), .B1_t (new_AGEMA_signal_14553), .B1_f (new_AGEMA_signal_14554), .Z0_t (MixColumnsOutput[79]), .Z0_f (new_AGEMA_signal_15983), .Z1_t (new_AGEMA_signal_15984), .Z1_f (new_AGEMA_signal_15985) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U27 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13892), .A1_t (new_AGEMA_signal_13893), .A1_f (new_AGEMA_signal_13894), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13664), .B1_t (new_AGEMA_signal_13665), .B1_f (new_AGEMA_signal_13666), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n149), .Z0_f (new_AGEMA_signal_14552), .Z1_t (new_AGEMA_signal_14553), .Z1_f (new_AGEMA_signal_14554) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U26 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n184), .A0_f (new_AGEMA_signal_14555), .A1_t (new_AGEMA_signal_14556), .A1_f (new_AGEMA_signal_14557), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13766), .B1_t (new_AGEMA_signal_13767), .B1_f (new_AGEMA_signal_13768), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n135), .Z0_f (new_AGEMA_signal_15230), .Z1_t (new_AGEMA_signal_15231), .Z1_f (new_AGEMA_signal_15232) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U25 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13895), .A1_t (new_AGEMA_signal_13896), .A1_f (new_AGEMA_signal_13897), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13871), .B1_t (new_AGEMA_signal_13872), .B1_f (new_AGEMA_signal_13873), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n184), .Z0_f (new_AGEMA_signal_14555), .Z1_t (new_AGEMA_signal_14556), .Z1_f (new_AGEMA_signal_14557) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U24 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n134), .A0_f (new_AGEMA_signal_15233), .A1_t (new_AGEMA_signal_15234), .A1_f (new_AGEMA_signal_15235), .B0_t (MixColumnsIns_MixOneColumnInst_1_n147), .B0_f (new_AGEMA_signal_14558), .B1_t (new_AGEMA_signal_14559), .B1_f (new_AGEMA_signal_14560), .Z0_t (MixColumnsOutput[78]), .Z0_f (new_AGEMA_signal_15986), .Z1_t (new_AGEMA_signal_15987), .Z1_f (new_AGEMA_signal_15988) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U23 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13895), .A1_t (new_AGEMA_signal_13896), .A1_f (new_AGEMA_signal_13897), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13667), .B1_t (new_AGEMA_signal_13668), .B1_f (new_AGEMA_signal_13669), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n147), .Z0_f (new_AGEMA_signal_14558), .Z1_t (new_AGEMA_signal_14559), .Z1_f (new_AGEMA_signal_14560) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U22 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n181), .A0_f (new_AGEMA_signal_14561), .A1_t (new_AGEMA_signal_14562), .A1_f (new_AGEMA_signal_14563), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13769), .B1_t (new_AGEMA_signal_13770), .B1_f (new_AGEMA_signal_13771), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n134), .Z0_f (new_AGEMA_signal_15233), .Z1_t (new_AGEMA_signal_15234), .Z1_f (new_AGEMA_signal_15235) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U21 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13898), .A1_t (new_AGEMA_signal_13899), .A1_f (new_AGEMA_signal_13900), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13874), .B1_t (new_AGEMA_signal_13875), .B1_f (new_AGEMA_signal_13876), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n181), .Z0_f (new_AGEMA_signal_14561), .Z1_t (new_AGEMA_signal_14562), .Z1_f (new_AGEMA_signal_14563) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U20 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n133), .A0_f (new_AGEMA_signal_15236), .A1_t (new_AGEMA_signal_15237), .A1_f (new_AGEMA_signal_15238), .B0_t (MixColumnsIns_MixOneColumnInst_1_n145), .B0_f (new_AGEMA_signal_14564), .B1_t (new_AGEMA_signal_14565), .B1_f (new_AGEMA_signal_14566), .Z0_t (MixColumnsOutput[77]), .Z0_f (new_AGEMA_signal_15989), .Z1_t (new_AGEMA_signal_15990), .Z1_f (new_AGEMA_signal_15991) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U19 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13898), .A1_t (new_AGEMA_signal_13899), .A1_f (new_AGEMA_signal_13900), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13670), .B1_t (new_AGEMA_signal_13671), .B1_f (new_AGEMA_signal_13672), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n145), .Z0_f (new_AGEMA_signal_14564), .Z1_t (new_AGEMA_signal_14565), .Z1_f (new_AGEMA_signal_14566) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U18 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n178), .A0_f (new_AGEMA_signal_14567), .A1_t (new_AGEMA_signal_14568), .A1_f (new_AGEMA_signal_14569), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13772), .B1_t (new_AGEMA_signal_13773), .B1_f (new_AGEMA_signal_13774), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n133), .Z0_f (new_AGEMA_signal_15236), .Z1_t (new_AGEMA_signal_15237), .Z1_f (new_AGEMA_signal_15238) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U17 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13901), .A1_t (new_AGEMA_signal_13902), .A1_f (new_AGEMA_signal_13903), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13877), .B1_t (new_AGEMA_signal_13878), .B1_f (new_AGEMA_signal_13879), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n178), .Z0_f (new_AGEMA_signal_14567), .Z1_t (new_AGEMA_signal_14568), .Z1_f (new_AGEMA_signal_14569) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U16 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n132), .A0_f (new_AGEMA_signal_15992), .A1_t (new_AGEMA_signal_15993), .A1_f (new_AGEMA_signal_15994), .B0_t (MixColumnsIns_MixOneColumnInst_1_n143), .B0_f (new_AGEMA_signal_15239), .B1_t (new_AGEMA_signal_15240), .B1_f (new_AGEMA_signal_15241), .Z0_t (MixColumnsOutput[76]), .Z0_f (new_AGEMA_signal_16877), .Z1_t (new_AGEMA_signal_16878), .Z1_f (new_AGEMA_signal_16879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U15 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13901), .A1_t (new_AGEMA_signal_13902), .A1_f (new_AGEMA_signal_13903), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]), .B0_f (new_AGEMA_signal_14600), .B1_t (new_AGEMA_signal_14601), .B1_f (new_AGEMA_signal_14602), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n143), .Z0_f (new_AGEMA_signal_15239), .Z1_t (new_AGEMA_signal_15240), .Z1_f (new_AGEMA_signal_15241) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U14 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n175), .A0_f (new_AGEMA_signal_15242), .A1_t (new_AGEMA_signal_15243), .A1_f (new_AGEMA_signal_15244), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13775), .B1_t (new_AGEMA_signal_13776), .B1_f (new_AGEMA_signal_13777), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n132), .Z0_f (new_AGEMA_signal_15992), .Z1_t (new_AGEMA_signal_15993), .Z1_f (new_AGEMA_signal_15994) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U13 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]), .A0_f (new_AGEMA_signal_14609), .A1_t (new_AGEMA_signal_14610), .A1_f (new_AGEMA_signal_14611), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13880), .B1_t (new_AGEMA_signal_13881), .B1_f (new_AGEMA_signal_13882), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n175), .Z0_f (new_AGEMA_signal_15242), .Z1_t (new_AGEMA_signal_15243), .Z1_f (new_AGEMA_signal_15244) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U12 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n131), .A0_f (new_AGEMA_signal_15995), .A1_t (new_AGEMA_signal_15996), .A1_f (new_AGEMA_signal_15997), .B0_t (MixColumnsIns_MixOneColumnInst_1_n140), .B0_f (new_AGEMA_signal_15245), .B1_t (new_AGEMA_signal_15246), .B1_f (new_AGEMA_signal_15247), .Z0_t (MixColumnsOutput[75]), .Z0_f (new_AGEMA_signal_16880), .Z1_t (new_AGEMA_signal_16881), .Z1_f (new_AGEMA_signal_16882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U11 ( .A0_t (MixColumnsInput[67]), .A0_f (new_AGEMA_signal_13904), .A1_t (new_AGEMA_signal_13905), .A1_f (new_AGEMA_signal_13906), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]), .B0_f (new_AGEMA_signal_14603), .B1_t (new_AGEMA_signal_14604), .B1_f (new_AGEMA_signal_14605), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n140), .Z0_f (new_AGEMA_signal_15245), .Z1_t (new_AGEMA_signal_15246), .Z1_f (new_AGEMA_signal_15247) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U10 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n172), .A0_f (new_AGEMA_signal_15248), .A1_t (new_AGEMA_signal_15249), .A1_f (new_AGEMA_signal_15250), .B0_t (MixColumnsInput[83]), .B0_f (new_AGEMA_signal_13778), .B1_t (new_AGEMA_signal_13779), .B1_f (new_AGEMA_signal_13780), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n131), .Z0_f (new_AGEMA_signal_15995), .Z1_t (new_AGEMA_signal_15996), .Z1_f (new_AGEMA_signal_15997) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U9 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]), .A0_f (new_AGEMA_signal_14612), .A1_t (new_AGEMA_signal_14613), .A1_f (new_AGEMA_signal_14614), .B0_t (MixColumnsInput[91]), .B0_f (new_AGEMA_signal_13883), .B1_t (new_AGEMA_signal_13884), .B1_f (new_AGEMA_signal_13885), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n172), .Z0_f (new_AGEMA_signal_15248), .Z1_t (new_AGEMA_signal_15249), .Z1_f (new_AGEMA_signal_15250) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U8 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n130), .A0_f (new_AGEMA_signal_15251), .A1_t (new_AGEMA_signal_15252), .A1_f (new_AGEMA_signal_15253), .B0_t (MixColumnsIns_MixOneColumnInst_1_n138), .B0_f (new_AGEMA_signal_14570), .B1_t (new_AGEMA_signal_14571), .B1_f (new_AGEMA_signal_14572), .Z0_t (MixColumnsOutput[74]), .Z0_f (new_AGEMA_signal_15998), .Z1_t (new_AGEMA_signal_15999), .Z1_f (new_AGEMA_signal_16000) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U7 ( .A0_t (MixColumnsInput[66]), .A0_f (new_AGEMA_signal_13907), .A1_t (new_AGEMA_signal_13908), .A1_f (new_AGEMA_signal_13909), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13679), .B1_t (new_AGEMA_signal_13680), .B1_f (new_AGEMA_signal_13681), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n138), .Z0_f (new_AGEMA_signal_14570), .Z1_t (new_AGEMA_signal_14571), .Z1_f (new_AGEMA_signal_14572) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U6 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n165), .A0_f (new_AGEMA_signal_14573), .A1_t (new_AGEMA_signal_14574), .A1_f (new_AGEMA_signal_14575), .B0_t (MixColumnsInput[82]), .B0_f (new_AGEMA_signal_13781), .B1_t (new_AGEMA_signal_13782), .B1_f (new_AGEMA_signal_13783), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n130), .Z0_f (new_AGEMA_signal_15251), .Z1_t (new_AGEMA_signal_15252), .Z1_f (new_AGEMA_signal_15253) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U5 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .A0_f (new_AGEMA_signal_13910), .A1_t (new_AGEMA_signal_13911), .A1_f (new_AGEMA_signal_13912), .B0_t (MixColumnsInput[90]), .B0_f (new_AGEMA_signal_13886), .B1_t (new_AGEMA_signal_13887), .B1_f (new_AGEMA_signal_13888), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n165), .Z0_f (new_AGEMA_signal_14573), .Z1_t (new_AGEMA_signal_14574), .Z1_f (new_AGEMA_signal_14575) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n129), .A0_f (new_AGEMA_signal_15254), .A1_t (new_AGEMA_signal_15255), .A1_f (new_AGEMA_signal_15256), .B0_t (MixColumnsInput[72]), .B0_f (new_AGEMA_signal_13031), .B1_t (new_AGEMA_signal_13032), .B1_f (new_AGEMA_signal_13033), .Z0_t (MixColumnsOutput[64]), .Z0_f (new_AGEMA_signal_16001), .Z1_t (new_AGEMA_signal_16002), .Z1_f (new_AGEMA_signal_16003) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n187), .A0_f (new_AGEMA_signal_14579), .A1_t (new_AGEMA_signal_14580), .A1_f (new_AGEMA_signal_14581), .B0_t (MixColumnsIns_MixOneColumnInst_1_n151), .B0_f (new_AGEMA_signal_14576), .B1_t (new_AGEMA_signal_14577), .B1_f (new_AGEMA_signal_14578), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n129), .Z0_f (new_AGEMA_signal_15254), .Z1_t (new_AGEMA_signal_15255), .Z1_f (new_AGEMA_signal_15256) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U2 ( .A0_t (MixColumnsInput[80]), .A0_f (new_AGEMA_signal_13196), .A1_t (new_AGEMA_signal_13197), .A1_f (new_AGEMA_signal_13198), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13871), .B1_t (new_AGEMA_signal_13872), .B1_f (new_AGEMA_signal_13873), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n151), .Z0_f (new_AGEMA_signal_14576), .Z1_t (new_AGEMA_signal_14577), .Z1_f (new_AGEMA_signal_14578) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U1 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13892), .A1_t (new_AGEMA_signal_13893), .A1_f (new_AGEMA_signal_13894), .B0_t (MixColumnsInput[88]), .B0_f (new_AGEMA_signal_13361), .B1_t (new_AGEMA_signal_13362), .B1_f (new_AGEMA_signal_13363), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n187), .Z0_f (new_AGEMA_signal_14579), .Z1_t (new_AGEMA_signal_14580), .Z1_f (new_AGEMA_signal_14581) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13871), .A1_t (new_AGEMA_signal_13872), .A1_f (new_AGEMA_signal_13873), .B0_t (MixColumnsInput[91]), .B0_f (new_AGEMA_signal_13883), .B1_t (new_AGEMA_signal_13884), .B1_f (new_AGEMA_signal_13885), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]), .Z0_f (new_AGEMA_signal_14582), .Z1_t (new_AGEMA_signal_14583), .Z1_f (new_AGEMA_signal_14584) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13871), .A1_t (new_AGEMA_signal_13872), .A1_f (new_AGEMA_signal_13873), .B0_t (MixColumnsInput[90]), .B0_f (new_AGEMA_signal_13886), .B1_t (new_AGEMA_signal_13887), .B1_f (new_AGEMA_signal_13888), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]), .Z0_f (new_AGEMA_signal_14585), .Z1_t (new_AGEMA_signal_14586), .Z1_f (new_AGEMA_signal_14587) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13871), .A1_t (new_AGEMA_signal_13872), .A1_f (new_AGEMA_signal_13873), .B0_t (MixColumnsInput[88]), .B0_f (new_AGEMA_signal_13361), .B1_t (new_AGEMA_signal_13362), .B1_f (new_AGEMA_signal_13363), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]), .Z0_f (new_AGEMA_signal_14588), .Z1_t (new_AGEMA_signal_14589), .Z1_f (new_AGEMA_signal_14590) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13766), .A1_t (new_AGEMA_signal_13767), .A1_f (new_AGEMA_signal_13768), .B0_t (MixColumnsInput[83]), .B0_f (new_AGEMA_signal_13778), .B1_t (new_AGEMA_signal_13779), .B1_f (new_AGEMA_signal_13780), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]), .Z0_f (new_AGEMA_signal_14591), .Z1_t (new_AGEMA_signal_14592), .Z1_f (new_AGEMA_signal_14593) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13766), .A1_t (new_AGEMA_signal_13767), .A1_f (new_AGEMA_signal_13768), .B0_t (MixColumnsInput[82]), .B0_f (new_AGEMA_signal_13781), .B1_t (new_AGEMA_signal_13782), .B1_f (new_AGEMA_signal_13783), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]), .Z0_f (new_AGEMA_signal_14594), .Z1_t (new_AGEMA_signal_14595), .Z1_f (new_AGEMA_signal_14596) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13766), .A1_t (new_AGEMA_signal_13767), .A1_f (new_AGEMA_signal_13768), .B0_t (MixColumnsInput[80]), .B0_f (new_AGEMA_signal_13196), .B1_t (new_AGEMA_signal_13197), .B1_f (new_AGEMA_signal_13198), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]), .Z0_f (new_AGEMA_signal_14597), .Z1_t (new_AGEMA_signal_14598), .Z1_f (new_AGEMA_signal_14599) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13661), .A1_t (new_AGEMA_signal_13662), .A1_f (new_AGEMA_signal_13663), .B0_t (MixColumnsInput[75]), .B0_f (new_AGEMA_signal_13673), .B1_t (new_AGEMA_signal_13674), .B1_f (new_AGEMA_signal_13675), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]), .Z0_f (new_AGEMA_signal_14600), .Z1_t (new_AGEMA_signal_14601), .Z1_f (new_AGEMA_signal_14602) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13661), .A1_t (new_AGEMA_signal_13662), .A1_f (new_AGEMA_signal_13663), .B0_t (MixColumnsInput[74]), .B0_f (new_AGEMA_signal_13676), .B1_t (new_AGEMA_signal_13677), .B1_f (new_AGEMA_signal_13678), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]), .Z0_f (new_AGEMA_signal_14603), .Z1_t (new_AGEMA_signal_14604), .Z1_f (new_AGEMA_signal_14605) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13661), .A1_t (new_AGEMA_signal_13662), .A1_f (new_AGEMA_signal_13663), .B0_t (MixColumnsInput[72]), .B0_f (new_AGEMA_signal_13031), .B1_t (new_AGEMA_signal_13032), .B1_f (new_AGEMA_signal_13033), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]), .Z0_f (new_AGEMA_signal_14606), .Z1_t (new_AGEMA_signal_14607), .Z1_f (new_AGEMA_signal_14608) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13892), .A1_t (new_AGEMA_signal_13893), .A1_f (new_AGEMA_signal_13894), .B0_t (MixColumnsInput[67]), .B0_f (new_AGEMA_signal_13904), .B1_t (new_AGEMA_signal_13905), .B1_f (new_AGEMA_signal_13906), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]), .Z0_f (new_AGEMA_signal_14609), .Z1_t (new_AGEMA_signal_14610), .Z1_f (new_AGEMA_signal_14611) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13892), .A1_t (new_AGEMA_signal_13893), .A1_f (new_AGEMA_signal_13894), .B0_t (MixColumnsInput[66]), .B0_f (new_AGEMA_signal_13907), .B1_t (new_AGEMA_signal_13908), .B1_f (new_AGEMA_signal_13909), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]), .Z0_f (new_AGEMA_signal_14612), .Z1_t (new_AGEMA_signal_14613), .Z1_f (new_AGEMA_signal_14614) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13892), .A1_t (new_AGEMA_signal_13893), .A1_f (new_AGEMA_signal_13894), .B0_t (MixColumnsInput[64]), .B0_f (new_AGEMA_signal_13394), .B1_t (new_AGEMA_signal_13395), .B1_f (new_AGEMA_signal_13396), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]), .Z0_f (new_AGEMA_signal_14615), .Z1_t (new_AGEMA_signal_14616), .Z1_f (new_AGEMA_signal_14617) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U96 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n192), .A0_f (new_AGEMA_signal_16004), .A1_t (new_AGEMA_signal_16005), .A1_f (new_AGEMA_signal_16006), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13700), .B1_t (new_AGEMA_signal_13701), .B1_f (new_AGEMA_signal_13702), .Z0_t (MixColumnsOutput[41]), .Z0_f (new_AGEMA_signal_16883), .Z1_t (new_AGEMA_signal_16884), .Z1_f (new_AGEMA_signal_16885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U95 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n191), .A0_f (new_AGEMA_signal_15320), .A1_t (new_AGEMA_signal_15321), .A1_f (new_AGEMA_signal_15322), .B0_t (MixColumnsIns_MixOneColumnInst_2_n190), .B0_f (new_AGEMA_signal_15308), .B1_t (new_AGEMA_signal_15309), .B1_f (new_AGEMA_signal_15310), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n192), .Z0_f (new_AGEMA_signal_16004), .Z1_t (new_AGEMA_signal_16005), .Z1_f (new_AGEMA_signal_16006) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U94 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n189), .A0_f (new_AGEMA_signal_15257), .A1_t (new_AGEMA_signal_15258), .A1_f (new_AGEMA_signal_15259), .B0_t (MixColumnsIns_MixOneColumnInst_2_n188), .B0_f (new_AGEMA_signal_14645), .B1_t (new_AGEMA_signal_14646), .B1_f (new_AGEMA_signal_14647), .Z0_t (MixColumnsOutput[40]), .Z0_f (new_AGEMA_signal_16007), .Z1_t (new_AGEMA_signal_16008), .Z1_f (new_AGEMA_signal_16009) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U93 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n187), .A0_f (new_AGEMA_signal_14675), .A1_t (new_AGEMA_signal_14676), .A1_f (new_AGEMA_signal_14677), .B0_t (MixColumnsInput[48]), .B0_f (new_AGEMA_signal_13064), .B1_t (new_AGEMA_signal_13065), .B1_f (new_AGEMA_signal_13066), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n189), .Z0_f (new_AGEMA_signal_15257), .Z1_t (new_AGEMA_signal_15258), .Z1_f (new_AGEMA_signal_15259) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U92 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n186), .A0_f (new_AGEMA_signal_15260), .A1_t (new_AGEMA_signal_15261), .A1_f (new_AGEMA_signal_15262), .B0_t (MixColumnsIns_MixOneColumnInst_2_n185), .B0_f (new_AGEMA_signal_14618), .B1_t (new_AGEMA_signal_14619), .B1_f (new_AGEMA_signal_14620), .Z0_t (MixColumnsOutput[39]), .Z0_f (new_AGEMA_signal_16010), .Z1_t (new_AGEMA_signal_16011), .Z1_f (new_AGEMA_signal_16012) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U91 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n184), .A0_f (new_AGEMA_signal_14651), .A1_t (new_AGEMA_signal_14652), .A1_f (new_AGEMA_signal_14653), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B0_f (new_AGEMA_signal_13913), .B1_t (new_AGEMA_signal_13914), .B1_f (new_AGEMA_signal_13915), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n186), .Z0_f (new_AGEMA_signal_15260), .Z1_t (new_AGEMA_signal_15261), .Z1_f (new_AGEMA_signal_15262) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U90 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n183), .A0_f (new_AGEMA_signal_15263), .A1_t (new_AGEMA_signal_15264), .A1_f (new_AGEMA_signal_15265), .B0_t (MixColumnsIns_MixOneColumnInst_2_n182), .B0_f (new_AGEMA_signal_14621), .B1_t (new_AGEMA_signal_14622), .B1_f (new_AGEMA_signal_14623), .Z0_t (MixColumnsOutput[38]), .Z0_f (new_AGEMA_signal_16013), .Z1_t (new_AGEMA_signal_16014), .Z1_f (new_AGEMA_signal_16015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U89 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n181), .A0_f (new_AGEMA_signal_14657), .A1_t (new_AGEMA_signal_14658), .A1_f (new_AGEMA_signal_14659), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13916), .B1_t (new_AGEMA_signal_13917), .B1_f (new_AGEMA_signal_13918), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n183), .Z0_f (new_AGEMA_signal_15263), .Z1_t (new_AGEMA_signal_15264), .Z1_f (new_AGEMA_signal_15265) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U88 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n180), .A0_f (new_AGEMA_signal_15266), .A1_t (new_AGEMA_signal_15267), .A1_f (new_AGEMA_signal_15268), .B0_t (MixColumnsIns_MixOneColumnInst_2_n179), .B0_f (new_AGEMA_signal_14624), .B1_t (new_AGEMA_signal_14625), .B1_f (new_AGEMA_signal_14626), .Z0_t (MixColumnsOutput[37]), .Z0_f (new_AGEMA_signal_16016), .Z1_t (new_AGEMA_signal_16017), .Z1_f (new_AGEMA_signal_16018) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U87 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n178), .A0_f (new_AGEMA_signal_14663), .A1_t (new_AGEMA_signal_14664), .A1_f (new_AGEMA_signal_14665), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13919), .B1_t (new_AGEMA_signal_13920), .B1_f (new_AGEMA_signal_13921), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n180), .Z0_f (new_AGEMA_signal_15266), .Z1_t (new_AGEMA_signal_15267), .Z1_f (new_AGEMA_signal_15268) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U86 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n177), .A0_f (new_AGEMA_signal_16019), .A1_t (new_AGEMA_signal_16020), .A1_f (new_AGEMA_signal_16021), .B0_t (MixColumnsIns_MixOneColumnInst_2_n176), .B0_f (new_AGEMA_signal_15281), .B1_t (new_AGEMA_signal_15282), .B1_f (new_AGEMA_signal_15283), .Z0_t (MixColumnsOutput[36]), .Z0_f (new_AGEMA_signal_16886), .Z1_t (new_AGEMA_signal_16887), .Z1_f (new_AGEMA_signal_16888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U85 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n175), .A0_f (new_AGEMA_signal_15338), .A1_t (new_AGEMA_signal_15339), .A1_f (new_AGEMA_signal_15340), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13922), .B1_t (new_AGEMA_signal_13923), .B1_f (new_AGEMA_signal_13924), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n177), .Z0_f (new_AGEMA_signal_16019), .Z1_t (new_AGEMA_signal_16020), .Z1_f (new_AGEMA_signal_16021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U84 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n174), .A0_f (new_AGEMA_signal_16022), .A1_t (new_AGEMA_signal_16023), .A1_f (new_AGEMA_signal_16024), .B0_t (MixColumnsIns_MixOneColumnInst_2_n173), .B0_f (new_AGEMA_signal_15284), .B1_t (new_AGEMA_signal_15285), .B1_f (new_AGEMA_signal_15286), .Z0_t (MixColumnsOutput[35]), .Z0_f (new_AGEMA_signal_16889), .Z1_t (new_AGEMA_signal_16890), .Z1_f (new_AGEMA_signal_16891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U83 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n172), .A0_f (new_AGEMA_signal_15344), .A1_t (new_AGEMA_signal_15345), .A1_f (new_AGEMA_signal_15346), .B0_t (MixColumnsInput[43]), .B0_f (new_AGEMA_signal_13925), .B1_t (new_AGEMA_signal_13926), .B1_f (new_AGEMA_signal_13927), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n174), .Z0_f (new_AGEMA_signal_16022), .Z1_t (new_AGEMA_signal_16023), .Z1_f (new_AGEMA_signal_16024) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U82 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n171), .A0_f (new_AGEMA_signal_15269), .A1_t (new_AGEMA_signal_15270), .A1_f (new_AGEMA_signal_15271), .B0_t (MixColumnsIns_MixOneColumnInst_2_n185), .B0_f (new_AGEMA_signal_14618), .B1_t (new_AGEMA_signal_14619), .B1_f (new_AGEMA_signal_14620), .Z0_t (MixColumnsOutput[63]), .Z0_f (new_AGEMA_signal_16025), .Z1_t (new_AGEMA_signal_16026), .Z1_f (new_AGEMA_signal_16027) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U81 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13682), .A1_t (new_AGEMA_signal_13683), .A1_f (new_AGEMA_signal_13684), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13790), .B1_t (new_AGEMA_signal_13791), .B1_f (new_AGEMA_signal_13792), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n185), .Z0_f (new_AGEMA_signal_14618), .Z1_t (new_AGEMA_signal_14619), .Z1_f (new_AGEMA_signal_14620) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U80 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13808), .A1_t (new_AGEMA_signal_13809), .A1_f (new_AGEMA_signal_13810), .B0_t (MixColumnsIns_MixOneColumnInst_2_n170), .B0_f (new_AGEMA_signal_14630), .B1_t (new_AGEMA_signal_14631), .B1_f (new_AGEMA_signal_14632), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n171), .Z0_f (new_AGEMA_signal_15269), .Z1_t (new_AGEMA_signal_15270), .Z1_f (new_AGEMA_signal_15271) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U79 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n169), .A0_f (new_AGEMA_signal_15272), .A1_t (new_AGEMA_signal_15273), .A1_f (new_AGEMA_signal_15274), .B0_t (MixColumnsIns_MixOneColumnInst_2_n182), .B0_f (new_AGEMA_signal_14621), .B1_t (new_AGEMA_signal_14622), .B1_f (new_AGEMA_signal_14623), .Z0_t (MixColumnsOutput[62]), .Z0_f (new_AGEMA_signal_16028), .Z1_t (new_AGEMA_signal_16029), .Z1_f (new_AGEMA_signal_16030) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U78 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .A0_f (new_AGEMA_signal_13685), .A1_t (new_AGEMA_signal_13686), .A1_f (new_AGEMA_signal_13687), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13793), .B1_t (new_AGEMA_signal_13794), .B1_f (new_AGEMA_signal_13795), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n182), .Z0_f (new_AGEMA_signal_14621), .Z1_t (new_AGEMA_signal_14622), .Z1_f (new_AGEMA_signal_14623) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U77 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13811), .A1_t (new_AGEMA_signal_13812), .A1_f (new_AGEMA_signal_13813), .B0_t (MixColumnsIns_MixOneColumnInst_2_n168), .B0_f (new_AGEMA_signal_14633), .B1_t (new_AGEMA_signal_14634), .B1_f (new_AGEMA_signal_14635), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n169), .Z0_f (new_AGEMA_signal_15272), .Z1_t (new_AGEMA_signal_15273), .Z1_f (new_AGEMA_signal_15274) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U76 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n167), .A0_f (new_AGEMA_signal_15275), .A1_t (new_AGEMA_signal_15276), .A1_f (new_AGEMA_signal_15277), .B0_t (MixColumnsIns_MixOneColumnInst_2_n166), .B0_f (new_AGEMA_signal_14627), .B1_t (new_AGEMA_signal_14628), .B1_f (new_AGEMA_signal_14629), .Z0_t (MixColumnsOutput[34]), .Z0_f (new_AGEMA_signal_16031), .Z1_t (new_AGEMA_signal_16032), .Z1_f (new_AGEMA_signal_16033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U75 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n165), .A0_f (new_AGEMA_signal_14669), .A1_t (new_AGEMA_signal_14670), .A1_f (new_AGEMA_signal_14671), .B0_t (MixColumnsInput[42]), .B0_f (new_AGEMA_signal_13928), .B1_t (new_AGEMA_signal_13929), .B1_f (new_AGEMA_signal_13930), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n167), .Z0_f (new_AGEMA_signal_15275), .Z1_t (new_AGEMA_signal_15276), .Z1_f (new_AGEMA_signal_15277) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U74 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n164), .A0_f (new_AGEMA_signal_15278), .A1_t (new_AGEMA_signal_15279), .A1_f (new_AGEMA_signal_15280), .B0_t (MixColumnsIns_MixOneColumnInst_2_n179), .B0_f (new_AGEMA_signal_14624), .B1_t (new_AGEMA_signal_14625), .B1_f (new_AGEMA_signal_14626), .Z0_t (MixColumnsOutput[61]), .Z0_f (new_AGEMA_signal_16034), .Z1_t (new_AGEMA_signal_16035), .Z1_f (new_AGEMA_signal_16036) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U73 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .A0_f (new_AGEMA_signal_13688), .A1_t (new_AGEMA_signal_13689), .A1_f (new_AGEMA_signal_13690), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13796), .B1_t (new_AGEMA_signal_13797), .B1_f (new_AGEMA_signal_13798), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n179), .Z0_f (new_AGEMA_signal_14624), .Z1_t (new_AGEMA_signal_14625), .Z1_f (new_AGEMA_signal_14626) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U72 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13814), .A1_t (new_AGEMA_signal_13815), .A1_f (new_AGEMA_signal_13816), .B0_t (MixColumnsIns_MixOneColumnInst_2_n163), .B0_f (new_AGEMA_signal_14636), .B1_t (new_AGEMA_signal_14637), .B1_f (new_AGEMA_signal_14638), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n164), .Z0_f (new_AGEMA_signal_15278), .Z1_t (new_AGEMA_signal_15279), .Z1_f (new_AGEMA_signal_15280) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U71 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n162), .A0_f (new_AGEMA_signal_16037), .A1_t (new_AGEMA_signal_16038), .A1_f (new_AGEMA_signal_16039), .B0_t (MixColumnsIns_MixOneColumnInst_2_n176), .B0_f (new_AGEMA_signal_15281), .B1_t (new_AGEMA_signal_15282), .B1_f (new_AGEMA_signal_15283), .Z0_t (MixColumnsOutput[60]), .Z0_f (new_AGEMA_signal_16892), .Z1_t (new_AGEMA_signal_16893), .Z1_f (new_AGEMA_signal_16894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U70 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .A0_f (new_AGEMA_signal_13691), .A1_t (new_AGEMA_signal_13692), .A1_f (new_AGEMA_signal_13693), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]), .B0_f (new_AGEMA_signal_14678), .B1_t (new_AGEMA_signal_14679), .B1_f (new_AGEMA_signal_14680), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n176), .Z0_f (new_AGEMA_signal_15281), .Z1_t (new_AGEMA_signal_15282), .Z1_f (new_AGEMA_signal_15283) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U69 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13817), .A1_t (new_AGEMA_signal_13818), .A1_f (new_AGEMA_signal_13819), .B0_t (MixColumnsIns_MixOneColumnInst_2_n161), .B0_f (new_AGEMA_signal_15302), .B1_t (new_AGEMA_signal_15303), .B1_f (new_AGEMA_signal_15304), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n162), .Z0_f (new_AGEMA_signal_16037), .Z1_t (new_AGEMA_signal_16038), .Z1_f (new_AGEMA_signal_16039) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U68 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n160), .A0_f (new_AGEMA_signal_16040), .A1_t (new_AGEMA_signal_16041), .A1_f (new_AGEMA_signal_16042), .B0_t (MixColumnsIns_MixOneColumnInst_2_n173), .B0_f (new_AGEMA_signal_15284), .B1_t (new_AGEMA_signal_15285), .B1_f (new_AGEMA_signal_15286), .Z0_t (MixColumnsOutput[59]), .Z0_f (new_AGEMA_signal_16895), .Z1_t (new_AGEMA_signal_16896), .Z1_f (new_AGEMA_signal_16897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U67 ( .A0_t (MixColumnsInput[51]), .A0_f (new_AGEMA_signal_13694), .A1_t (new_AGEMA_signal_13695), .A1_f (new_AGEMA_signal_13696), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]), .B0_f (new_AGEMA_signal_14681), .B1_t (new_AGEMA_signal_14682), .B1_f (new_AGEMA_signal_14683), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n173), .Z0_f (new_AGEMA_signal_15284), .Z1_t (new_AGEMA_signal_15285), .Z1_f (new_AGEMA_signal_15286) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U66 ( .A0_t (MixColumnsInput[35]), .A0_f (new_AGEMA_signal_13820), .A1_t (new_AGEMA_signal_13821), .A1_f (new_AGEMA_signal_13822), .B0_t (MixColumnsIns_MixOneColumnInst_2_n159), .B0_f (new_AGEMA_signal_15311), .B1_t (new_AGEMA_signal_15312), .B1_f (new_AGEMA_signal_15313), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n160), .Z0_f (new_AGEMA_signal_16040), .Z1_t (new_AGEMA_signal_16041), .Z1_f (new_AGEMA_signal_16042) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U65 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n158), .A0_f (new_AGEMA_signal_15287), .A1_t (new_AGEMA_signal_15288), .A1_f (new_AGEMA_signal_15289), .B0_t (MixColumnsIns_MixOneColumnInst_2_n166), .B0_f (new_AGEMA_signal_14627), .B1_t (new_AGEMA_signal_14628), .B1_f (new_AGEMA_signal_14629), .Z0_t (MixColumnsOutput[58]), .Z0_f (new_AGEMA_signal_16043), .Z1_t (new_AGEMA_signal_16044), .Z1_f (new_AGEMA_signal_16045) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U64 ( .A0_t (MixColumnsInput[50]), .A0_f (new_AGEMA_signal_13697), .A1_t (new_AGEMA_signal_13698), .A1_f (new_AGEMA_signal_13699), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13805), .B1_t (new_AGEMA_signal_13806), .B1_f (new_AGEMA_signal_13807), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n166), .Z0_f (new_AGEMA_signal_14627), .Z1_t (new_AGEMA_signal_14628), .Z1_f (new_AGEMA_signal_14629) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U63 ( .A0_t (MixColumnsInput[34]), .A0_f (new_AGEMA_signal_13823), .A1_t (new_AGEMA_signal_13824), .A1_f (new_AGEMA_signal_13825), .B0_t (MixColumnsIns_MixOneColumnInst_2_n157), .B0_f (new_AGEMA_signal_14639), .B1_t (new_AGEMA_signal_14640), .B1_f (new_AGEMA_signal_14641), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n158), .Z0_f (new_AGEMA_signal_15287), .Z1_t (new_AGEMA_signal_15288), .Z1_f (new_AGEMA_signal_15289) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U62 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n156), .A0_f (new_AGEMA_signal_16046), .A1_t (new_AGEMA_signal_16047), .A1_f (new_AGEMA_signal_16048), .B0_t (MixColumnsIns_MixOneColumnInst_2_n155), .B0_f (new_AGEMA_signal_15305), .B1_t (new_AGEMA_signal_15306), .B1_f (new_AGEMA_signal_15307), .Z0_t (MixColumnsOutput[57]), .Z0_f (new_AGEMA_signal_16898), .Z1_t (new_AGEMA_signal_16899), .Z1_f (new_AGEMA_signal_16900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U61 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .A0_f (new_AGEMA_signal_13826), .A1_t (new_AGEMA_signal_13827), .A1_f (new_AGEMA_signal_13828), .B0_t (MixColumnsIns_MixOneColumnInst_2_n154), .B0_f (new_AGEMA_signal_15317), .B1_t (new_AGEMA_signal_15318), .B1_f (new_AGEMA_signal_15319), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n156), .Z0_f (new_AGEMA_signal_16046), .Z1_t (new_AGEMA_signal_16047), .Z1_f (new_AGEMA_signal_16048) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U60 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n153), .A0_f (new_AGEMA_signal_15290), .A1_t (new_AGEMA_signal_15291), .A1_f (new_AGEMA_signal_15292), .B0_t (MixColumnsIns_MixOneColumnInst_2_n152), .B0_f (new_AGEMA_signal_14642), .B1_t (new_AGEMA_signal_14643), .B1_f (new_AGEMA_signal_14644), .Z0_t (MixColumnsOutput[56]), .Z0_f (new_AGEMA_signal_16049), .Z1_t (new_AGEMA_signal_16050), .Z1_f (new_AGEMA_signal_16051) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U59 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n151), .A0_f (new_AGEMA_signal_14672), .A1_t (new_AGEMA_signal_14673), .A1_f (new_AGEMA_signal_14674), .B0_t (MixColumnsInput[32]), .B0_f (new_AGEMA_signal_13262), .B1_t (new_AGEMA_signal_13263), .B1_f (new_AGEMA_signal_13264), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n153), .Z0_f (new_AGEMA_signal_15290), .Z1_t (new_AGEMA_signal_15291), .Z1_f (new_AGEMA_signal_15292) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U58 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n150), .A0_f (new_AGEMA_signal_15293), .A1_t (new_AGEMA_signal_15294), .A1_f (new_AGEMA_signal_15295), .B0_t (MixColumnsIns_MixOneColumnInst_2_n170), .B0_f (new_AGEMA_signal_14630), .B1_t (new_AGEMA_signal_14631), .B1_f (new_AGEMA_signal_14632), .Z0_t (MixColumnsOutput[55]), .Z0_f (new_AGEMA_signal_16052), .Z1_t (new_AGEMA_signal_16053), .Z1_f (new_AGEMA_signal_16054) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U57 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13913), .A1_t (new_AGEMA_signal_13914), .A1_f (new_AGEMA_signal_13915), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13685), .B1_t (new_AGEMA_signal_13686), .B1_f (new_AGEMA_signal_13687), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n170), .Z0_f (new_AGEMA_signal_14630), .Z1_t (new_AGEMA_signal_14631), .Z1_f (new_AGEMA_signal_14632) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U56 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13787), .A1_t (new_AGEMA_signal_13788), .A1_f (new_AGEMA_signal_13789), .B0_t (MixColumnsIns_MixOneColumnInst_2_n149), .B0_f (new_AGEMA_signal_14648), .B1_t (new_AGEMA_signal_14649), .B1_f (new_AGEMA_signal_14650), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n150), .Z0_f (new_AGEMA_signal_15293), .Z1_t (new_AGEMA_signal_15294), .Z1_f (new_AGEMA_signal_15295) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U55 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n148), .A0_f (new_AGEMA_signal_15296), .A1_t (new_AGEMA_signal_15297), .A1_f (new_AGEMA_signal_15298), .B0_t (MixColumnsIns_MixOneColumnInst_2_n168), .B0_f (new_AGEMA_signal_14633), .B1_t (new_AGEMA_signal_14634), .B1_f (new_AGEMA_signal_14635), .Z0_t (MixColumnsOutput[54]), .Z0_f (new_AGEMA_signal_16055), .Z1_t (new_AGEMA_signal_16056), .Z1_f (new_AGEMA_signal_16057) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U54 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .A0_f (new_AGEMA_signal_13916), .A1_t (new_AGEMA_signal_13917), .A1_f (new_AGEMA_signal_13918), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13688), .B1_t (new_AGEMA_signal_13689), .B1_f (new_AGEMA_signal_13690), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n168), .Z0_f (new_AGEMA_signal_14633), .Z1_t (new_AGEMA_signal_14634), .Z1_f (new_AGEMA_signal_14635) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U53 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .A0_f (new_AGEMA_signal_13790), .A1_t (new_AGEMA_signal_13791), .A1_f (new_AGEMA_signal_13792), .B0_t (MixColumnsIns_MixOneColumnInst_2_n147), .B0_f (new_AGEMA_signal_14654), .B1_t (new_AGEMA_signal_14655), .B1_f (new_AGEMA_signal_14656), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n148), .Z0_f (new_AGEMA_signal_15296), .Z1_t (new_AGEMA_signal_15297), .Z1_f (new_AGEMA_signal_15298) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U52 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n146), .A0_f (new_AGEMA_signal_15299), .A1_t (new_AGEMA_signal_15300), .A1_f (new_AGEMA_signal_15301), .B0_t (MixColumnsIns_MixOneColumnInst_2_n163), .B0_f (new_AGEMA_signal_14636), .B1_t (new_AGEMA_signal_14637), .B1_f (new_AGEMA_signal_14638), .Z0_t (MixColumnsOutput[53]), .Z0_f (new_AGEMA_signal_16058), .Z1_t (new_AGEMA_signal_16059), .Z1_f (new_AGEMA_signal_16060) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U51 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .A0_f (new_AGEMA_signal_13919), .A1_t (new_AGEMA_signal_13920), .A1_f (new_AGEMA_signal_13921), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13691), .B1_t (new_AGEMA_signal_13692), .B1_f (new_AGEMA_signal_13693), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n163), .Z0_f (new_AGEMA_signal_14636), .Z1_t (new_AGEMA_signal_14637), .Z1_f (new_AGEMA_signal_14638) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U50 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .A0_f (new_AGEMA_signal_13793), .A1_t (new_AGEMA_signal_13794), .A1_f (new_AGEMA_signal_13795), .B0_t (MixColumnsIns_MixOneColumnInst_2_n145), .B0_f (new_AGEMA_signal_14660), .B1_t (new_AGEMA_signal_14661), .B1_f (new_AGEMA_signal_14662), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n146), .Z0_f (new_AGEMA_signal_15299), .Z1_t (new_AGEMA_signal_15300), .Z1_f (new_AGEMA_signal_15301) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U49 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n144), .A0_f (new_AGEMA_signal_16061), .A1_t (new_AGEMA_signal_16062), .A1_f (new_AGEMA_signal_16063), .B0_t (MixColumnsIns_MixOneColumnInst_2_n161), .B0_f (new_AGEMA_signal_15302), .B1_t (new_AGEMA_signal_15303), .B1_f (new_AGEMA_signal_15304), .Z0_t (MixColumnsOutput[52]), .Z0_f (new_AGEMA_signal_16901), .Z1_t (new_AGEMA_signal_16902), .Z1_f (new_AGEMA_signal_16903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U48 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .A0_f (new_AGEMA_signal_13922), .A1_t (new_AGEMA_signal_13923), .A1_f (new_AGEMA_signal_13924), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]), .B0_f (new_AGEMA_signal_14687), .B1_t (new_AGEMA_signal_14688), .B1_f (new_AGEMA_signal_14689), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n161), .Z0_f (new_AGEMA_signal_15302), .Z1_t (new_AGEMA_signal_15303), .Z1_f (new_AGEMA_signal_15304) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U47 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .A0_f (new_AGEMA_signal_13796), .A1_t (new_AGEMA_signal_13797), .A1_f (new_AGEMA_signal_13798), .B0_t (MixColumnsIns_MixOneColumnInst_2_n143), .B0_f (new_AGEMA_signal_15335), .B1_t (new_AGEMA_signal_15336), .B1_f (new_AGEMA_signal_15337), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n144), .Z0_f (new_AGEMA_signal_16061), .Z1_t (new_AGEMA_signal_16062), .Z1_f (new_AGEMA_signal_16063) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U46 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n142), .A0_f (new_AGEMA_signal_16064), .A1_t (new_AGEMA_signal_16065), .A1_f (new_AGEMA_signal_16066), .B0_t (MixColumnsIns_MixOneColumnInst_2_n155), .B0_f (new_AGEMA_signal_15305), .B1_t (new_AGEMA_signal_15306), .B1_f (new_AGEMA_signal_15307), .Z0_t (MixColumnsOutput[33]), .Z0_f (new_AGEMA_signal_16904), .Z1_t (new_AGEMA_signal_16905), .Z1_f (new_AGEMA_signal_16906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U45 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .A0_f (new_AGEMA_signal_13700), .A1_t (new_AGEMA_signal_13701), .A1_f (new_AGEMA_signal_13702), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]), .B0_f (new_AGEMA_signal_14684), .B1_t (new_AGEMA_signal_14685), .B1_f (new_AGEMA_signal_14686), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n155), .Z0_f (new_AGEMA_signal_15305), .Z1_t (new_AGEMA_signal_15306), .Z1_f (new_AGEMA_signal_15307) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U44 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .A0_f (new_AGEMA_signal_13931), .A1_t (new_AGEMA_signal_13932), .A1_f (new_AGEMA_signal_13933), .B0_t (MixColumnsIns_MixOneColumnInst_2_n190), .B0_f (new_AGEMA_signal_15308), .B1_t (new_AGEMA_signal_15309), .B1_f (new_AGEMA_signal_15310), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n142), .Z0_f (new_AGEMA_signal_16064), .Z1_t (new_AGEMA_signal_16065), .Z1_f (new_AGEMA_signal_16066) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U43 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .A0_f (new_AGEMA_signal_13805), .A1_t (new_AGEMA_signal_13806), .A1_f (new_AGEMA_signal_13807), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]), .B0_f (new_AGEMA_signal_14711), .B1_t (new_AGEMA_signal_14712), .B1_f (new_AGEMA_signal_14713), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n190), .Z0_f (new_AGEMA_signal_15308), .Z1_t (new_AGEMA_signal_15309), .Z1_f (new_AGEMA_signal_15310) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U42 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n141), .A0_f (new_AGEMA_signal_16067), .A1_t (new_AGEMA_signal_16068), .A1_f (new_AGEMA_signal_16069), .B0_t (MixColumnsIns_MixOneColumnInst_2_n159), .B0_f (new_AGEMA_signal_15311), .B1_t (new_AGEMA_signal_15312), .B1_f (new_AGEMA_signal_15313), .Z0_t (MixColumnsOutput[51]), .Z0_f (new_AGEMA_signal_16907), .Z1_t (new_AGEMA_signal_16908), .Z1_f (new_AGEMA_signal_16909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U41 ( .A0_t (MixColumnsInput[43]), .A0_f (new_AGEMA_signal_13925), .A1_t (new_AGEMA_signal_13926), .A1_f (new_AGEMA_signal_13927), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]), .B0_f (new_AGEMA_signal_14690), .B1_t (new_AGEMA_signal_14691), .B1_f (new_AGEMA_signal_14692), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n159), .Z0_f (new_AGEMA_signal_15311), .Z1_t (new_AGEMA_signal_15312), .Z1_f (new_AGEMA_signal_15313) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U40 ( .A0_t (MixColumnsInput[59]), .A0_f (new_AGEMA_signal_13799), .A1_t (new_AGEMA_signal_13800), .A1_f (new_AGEMA_signal_13801), .B0_t (MixColumnsIns_MixOneColumnInst_2_n140), .B0_f (new_AGEMA_signal_15341), .B1_t (new_AGEMA_signal_15342), .B1_f (new_AGEMA_signal_15343), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n141), .Z0_f (new_AGEMA_signal_16067), .Z1_t (new_AGEMA_signal_16068), .Z1_f (new_AGEMA_signal_16069) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U39 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n139), .A0_f (new_AGEMA_signal_15314), .A1_t (new_AGEMA_signal_15315), .A1_f (new_AGEMA_signal_15316), .B0_t (MixColumnsIns_MixOneColumnInst_2_n157), .B0_f (new_AGEMA_signal_14639), .B1_t (new_AGEMA_signal_14640), .B1_f (new_AGEMA_signal_14641), .Z0_t (MixColumnsOutput[50]), .Z0_f (new_AGEMA_signal_16070), .Z1_t (new_AGEMA_signal_16071), .Z1_f (new_AGEMA_signal_16072) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U38 ( .A0_t (MixColumnsInput[42]), .A0_f (new_AGEMA_signal_13928), .A1_t (new_AGEMA_signal_13929), .A1_f (new_AGEMA_signal_13930), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13700), .B1_t (new_AGEMA_signal_13701), .B1_f (new_AGEMA_signal_13702), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n157), .Z0_f (new_AGEMA_signal_14639), .Z1_t (new_AGEMA_signal_14640), .Z1_f (new_AGEMA_signal_14641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U37 ( .A0_t (MixColumnsInput[58]), .A0_f (new_AGEMA_signal_13802), .A1_t (new_AGEMA_signal_13803), .A1_f (new_AGEMA_signal_13804), .B0_t (MixColumnsIns_MixOneColumnInst_2_n138), .B0_f (new_AGEMA_signal_14666), .B1_t (new_AGEMA_signal_14667), .B1_f (new_AGEMA_signal_14668), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n139), .Z0_f (new_AGEMA_signal_15314), .Z1_t (new_AGEMA_signal_15315), .Z1_f (new_AGEMA_signal_15316) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U36 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n137), .A0_f (new_AGEMA_signal_16073), .A1_t (new_AGEMA_signal_16074), .A1_f (new_AGEMA_signal_16075), .B0_t (MixColumnsIns_MixOneColumnInst_2_n154), .B0_f (new_AGEMA_signal_15317), .B1_t (new_AGEMA_signal_15318), .B1_f (new_AGEMA_signal_15319), .Z0_t (MixColumnsOutput[49]), .Z0_f (new_AGEMA_signal_16910), .Z1_t (new_AGEMA_signal_16911), .Z1_f (new_AGEMA_signal_16912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U35 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]), .A0_f (new_AGEMA_signal_14693), .A1_t (new_AGEMA_signal_14694), .A1_f (new_AGEMA_signal_14695), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13931), .B1_t (new_AGEMA_signal_13932), .B1_f (new_AGEMA_signal_13933), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n154), .Z0_f (new_AGEMA_signal_15317), .Z1_t (new_AGEMA_signal_15318), .Z1_f (new_AGEMA_signal_15319) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U34 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n191), .A0_f (new_AGEMA_signal_15320), .A1_t (new_AGEMA_signal_15321), .A1_f (new_AGEMA_signal_15322), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13805), .B1_t (new_AGEMA_signal_13806), .B1_f (new_AGEMA_signal_13807), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n137), .Z0_f (new_AGEMA_signal_16073), .Z1_t (new_AGEMA_signal_16074), .Z1_f (new_AGEMA_signal_16075) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U33 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]), .A0_f (new_AGEMA_signal_14702), .A1_t (new_AGEMA_signal_14703), .A1_f (new_AGEMA_signal_14704), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .B0_f (new_AGEMA_signal_13826), .B1_t (new_AGEMA_signal_13827), .B1_f (new_AGEMA_signal_13828), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n191), .Z0_f (new_AGEMA_signal_15320), .Z1_t (new_AGEMA_signal_15321), .Z1_f (new_AGEMA_signal_15322) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U32 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n136), .A0_f (new_AGEMA_signal_15323), .A1_t (new_AGEMA_signal_15324), .A1_f (new_AGEMA_signal_15325), .B0_t (MixColumnsIns_MixOneColumnInst_2_n152), .B0_f (new_AGEMA_signal_14642), .B1_t (new_AGEMA_signal_14643), .B1_f (new_AGEMA_signal_14644), .Z0_t (MixColumnsOutput[48]), .Z0_f (new_AGEMA_signal_16076), .Z1_t (new_AGEMA_signal_16077), .Z1_f (new_AGEMA_signal_16078) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U31 ( .A0_t (MixColumnsInput[40]), .A0_f (new_AGEMA_signal_13427), .A1_t (new_AGEMA_signal_13428), .A1_f (new_AGEMA_signal_13429), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13682), .B1_t (new_AGEMA_signal_13683), .B1_f (new_AGEMA_signal_13684), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n152), .Z0_f (new_AGEMA_signal_14642), .Z1_t (new_AGEMA_signal_14643), .Z1_f (new_AGEMA_signal_14644) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U30 ( .A0_t (MixColumnsInput[56]), .A0_f (new_AGEMA_signal_13229), .A1_t (new_AGEMA_signal_13230), .A1_f (new_AGEMA_signal_13231), .B0_t (MixColumnsIns_MixOneColumnInst_2_n188), .B0_f (new_AGEMA_signal_14645), .B1_t (new_AGEMA_signal_14646), .B1_f (new_AGEMA_signal_14647), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n136), .Z0_f (new_AGEMA_signal_15323), .Z1_t (new_AGEMA_signal_15324), .Z1_f (new_AGEMA_signal_15325) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U29 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13913), .A1_t (new_AGEMA_signal_13914), .A1_f (new_AGEMA_signal_13915), .B0_t (MixColumnsInput[32]), .B0_f (new_AGEMA_signal_13262), .B1_t (new_AGEMA_signal_13263), .B1_f (new_AGEMA_signal_13264), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n188), .Z0_f (new_AGEMA_signal_14645), .Z1_t (new_AGEMA_signal_14646), .Z1_f (new_AGEMA_signal_14647) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U28 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n135), .A0_f (new_AGEMA_signal_15326), .A1_t (new_AGEMA_signal_15327), .A1_f (new_AGEMA_signal_15328), .B0_t (MixColumnsIns_MixOneColumnInst_2_n149), .B0_f (new_AGEMA_signal_14648), .B1_t (new_AGEMA_signal_14649), .B1_f (new_AGEMA_signal_14650), .Z0_t (MixColumnsOutput[47]), .Z0_f (new_AGEMA_signal_16079), .Z1_t (new_AGEMA_signal_16080), .Z1_f (new_AGEMA_signal_16081) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U27 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13808), .A1_t (new_AGEMA_signal_13809), .A1_f (new_AGEMA_signal_13810), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13916), .B1_t (new_AGEMA_signal_13917), .B1_f (new_AGEMA_signal_13918), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n149), .Z0_f (new_AGEMA_signal_14648), .Z1_t (new_AGEMA_signal_14649), .Z1_f (new_AGEMA_signal_14650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U26 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n184), .A0_f (new_AGEMA_signal_14651), .A1_t (new_AGEMA_signal_14652), .A1_f (new_AGEMA_signal_14653), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13682), .B1_t (new_AGEMA_signal_13683), .B1_f (new_AGEMA_signal_13684), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n135), .Z0_f (new_AGEMA_signal_15326), .Z1_t (new_AGEMA_signal_15327), .Z1_f (new_AGEMA_signal_15328) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U25 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13811), .A1_t (new_AGEMA_signal_13812), .A1_f (new_AGEMA_signal_13813), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13787), .B1_t (new_AGEMA_signal_13788), .B1_f (new_AGEMA_signal_13789), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n184), .Z0_f (new_AGEMA_signal_14651), .Z1_t (new_AGEMA_signal_14652), .Z1_f (new_AGEMA_signal_14653) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U24 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n134), .A0_f (new_AGEMA_signal_15329), .A1_t (new_AGEMA_signal_15330), .A1_f (new_AGEMA_signal_15331), .B0_t (MixColumnsIns_MixOneColumnInst_2_n147), .B0_f (new_AGEMA_signal_14654), .B1_t (new_AGEMA_signal_14655), .B1_f (new_AGEMA_signal_14656), .Z0_t (MixColumnsOutput[46]), .Z0_f (new_AGEMA_signal_16082), .Z1_t (new_AGEMA_signal_16083), .Z1_f (new_AGEMA_signal_16084) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U23 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13811), .A1_t (new_AGEMA_signal_13812), .A1_f (new_AGEMA_signal_13813), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13919), .B1_t (new_AGEMA_signal_13920), .B1_f (new_AGEMA_signal_13921), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n147), .Z0_f (new_AGEMA_signal_14654), .Z1_t (new_AGEMA_signal_14655), .Z1_f (new_AGEMA_signal_14656) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U22 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n181), .A0_f (new_AGEMA_signal_14657), .A1_t (new_AGEMA_signal_14658), .A1_f (new_AGEMA_signal_14659), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13685), .B1_t (new_AGEMA_signal_13686), .B1_f (new_AGEMA_signal_13687), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n134), .Z0_f (new_AGEMA_signal_15329), .Z1_t (new_AGEMA_signal_15330), .Z1_f (new_AGEMA_signal_15331) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U21 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13814), .A1_t (new_AGEMA_signal_13815), .A1_f (new_AGEMA_signal_13816), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13790), .B1_t (new_AGEMA_signal_13791), .B1_f (new_AGEMA_signal_13792), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n181), .Z0_f (new_AGEMA_signal_14657), .Z1_t (new_AGEMA_signal_14658), .Z1_f (new_AGEMA_signal_14659) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U20 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n133), .A0_f (new_AGEMA_signal_15332), .A1_t (new_AGEMA_signal_15333), .A1_f (new_AGEMA_signal_15334), .B0_t (MixColumnsIns_MixOneColumnInst_2_n145), .B0_f (new_AGEMA_signal_14660), .B1_t (new_AGEMA_signal_14661), .B1_f (new_AGEMA_signal_14662), .Z0_t (MixColumnsOutput[45]), .Z0_f (new_AGEMA_signal_16085), .Z1_t (new_AGEMA_signal_16086), .Z1_f (new_AGEMA_signal_16087) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U19 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13814), .A1_t (new_AGEMA_signal_13815), .A1_f (new_AGEMA_signal_13816), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13922), .B1_t (new_AGEMA_signal_13923), .B1_f (new_AGEMA_signal_13924), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n145), .Z0_f (new_AGEMA_signal_14660), .Z1_t (new_AGEMA_signal_14661), .Z1_f (new_AGEMA_signal_14662) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U18 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n178), .A0_f (new_AGEMA_signal_14663), .A1_t (new_AGEMA_signal_14664), .A1_f (new_AGEMA_signal_14665), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13688), .B1_t (new_AGEMA_signal_13689), .B1_f (new_AGEMA_signal_13690), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n133), .Z0_f (new_AGEMA_signal_15332), .Z1_t (new_AGEMA_signal_15333), .Z1_f (new_AGEMA_signal_15334) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U17 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13817), .A1_t (new_AGEMA_signal_13818), .A1_f (new_AGEMA_signal_13819), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13793), .B1_t (new_AGEMA_signal_13794), .B1_f (new_AGEMA_signal_13795), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n178), .Z0_f (new_AGEMA_signal_14663), .Z1_t (new_AGEMA_signal_14664), .Z1_f (new_AGEMA_signal_14665) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U16 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n132), .A0_f (new_AGEMA_signal_16088), .A1_t (new_AGEMA_signal_16089), .A1_f (new_AGEMA_signal_16090), .B0_t (MixColumnsIns_MixOneColumnInst_2_n143), .B0_f (new_AGEMA_signal_15335), .B1_t (new_AGEMA_signal_15336), .B1_f (new_AGEMA_signal_15337), .Z0_t (MixColumnsOutput[44]), .Z0_f (new_AGEMA_signal_16913), .Z1_t (new_AGEMA_signal_16914), .Z1_f (new_AGEMA_signal_16915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U15 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13817), .A1_t (new_AGEMA_signal_13818), .A1_f (new_AGEMA_signal_13819), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]), .B0_f (new_AGEMA_signal_14696), .B1_t (new_AGEMA_signal_14697), .B1_f (new_AGEMA_signal_14698), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n143), .Z0_f (new_AGEMA_signal_15335), .Z1_t (new_AGEMA_signal_15336), .Z1_f (new_AGEMA_signal_15337) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U14 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n175), .A0_f (new_AGEMA_signal_15338), .A1_t (new_AGEMA_signal_15339), .A1_f (new_AGEMA_signal_15340), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13691), .B1_t (new_AGEMA_signal_13692), .B1_f (new_AGEMA_signal_13693), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n132), .Z0_f (new_AGEMA_signal_16088), .Z1_t (new_AGEMA_signal_16089), .Z1_f (new_AGEMA_signal_16090) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U13 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]), .A0_f (new_AGEMA_signal_14705), .A1_t (new_AGEMA_signal_14706), .A1_f (new_AGEMA_signal_14707), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13796), .B1_t (new_AGEMA_signal_13797), .B1_f (new_AGEMA_signal_13798), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n175), .Z0_f (new_AGEMA_signal_15338), .Z1_t (new_AGEMA_signal_15339), .Z1_f (new_AGEMA_signal_15340) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U12 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n131), .A0_f (new_AGEMA_signal_16091), .A1_t (new_AGEMA_signal_16092), .A1_f (new_AGEMA_signal_16093), .B0_t (MixColumnsIns_MixOneColumnInst_2_n140), .B0_f (new_AGEMA_signal_15341), .B1_t (new_AGEMA_signal_15342), .B1_f (new_AGEMA_signal_15343), .Z0_t (MixColumnsOutput[43]), .Z0_f (new_AGEMA_signal_16916), .Z1_t (new_AGEMA_signal_16917), .Z1_f (new_AGEMA_signal_16918) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U11 ( .A0_t (MixColumnsInput[35]), .A0_f (new_AGEMA_signal_13820), .A1_t (new_AGEMA_signal_13821), .A1_f (new_AGEMA_signal_13822), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]), .B0_f (new_AGEMA_signal_14699), .B1_t (new_AGEMA_signal_14700), .B1_f (new_AGEMA_signal_14701), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n140), .Z0_f (new_AGEMA_signal_15341), .Z1_t (new_AGEMA_signal_15342), .Z1_f (new_AGEMA_signal_15343) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U10 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n172), .A0_f (new_AGEMA_signal_15344), .A1_t (new_AGEMA_signal_15345), .A1_f (new_AGEMA_signal_15346), .B0_t (MixColumnsInput[51]), .B0_f (new_AGEMA_signal_13694), .B1_t (new_AGEMA_signal_13695), .B1_f (new_AGEMA_signal_13696), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n131), .Z0_f (new_AGEMA_signal_16091), .Z1_t (new_AGEMA_signal_16092), .Z1_f (new_AGEMA_signal_16093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U9 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]), .A0_f (new_AGEMA_signal_14708), .A1_t (new_AGEMA_signal_14709), .A1_f (new_AGEMA_signal_14710), .B0_t (MixColumnsInput[59]), .B0_f (new_AGEMA_signal_13799), .B1_t (new_AGEMA_signal_13800), .B1_f (new_AGEMA_signal_13801), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n172), .Z0_f (new_AGEMA_signal_15344), .Z1_t (new_AGEMA_signal_15345), .Z1_f (new_AGEMA_signal_15346) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U8 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n130), .A0_f (new_AGEMA_signal_15347), .A1_t (new_AGEMA_signal_15348), .A1_f (new_AGEMA_signal_15349), .B0_t (MixColumnsIns_MixOneColumnInst_2_n138), .B0_f (new_AGEMA_signal_14666), .B1_t (new_AGEMA_signal_14667), .B1_f (new_AGEMA_signal_14668), .Z0_t (MixColumnsOutput[42]), .Z0_f (new_AGEMA_signal_16094), .Z1_t (new_AGEMA_signal_16095), .Z1_f (new_AGEMA_signal_16096) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U7 ( .A0_t (MixColumnsInput[34]), .A0_f (new_AGEMA_signal_13823), .A1_t (new_AGEMA_signal_13824), .A1_f (new_AGEMA_signal_13825), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13931), .B1_t (new_AGEMA_signal_13932), .B1_f (new_AGEMA_signal_13933), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n138), .Z0_f (new_AGEMA_signal_14666), .Z1_t (new_AGEMA_signal_14667), .Z1_f (new_AGEMA_signal_14668) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U6 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n165), .A0_f (new_AGEMA_signal_14669), .A1_t (new_AGEMA_signal_14670), .A1_f (new_AGEMA_signal_14671), .B0_t (MixColumnsInput[50]), .B0_f (new_AGEMA_signal_13697), .B1_t (new_AGEMA_signal_13698), .B1_f (new_AGEMA_signal_13699), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n130), .Z0_f (new_AGEMA_signal_15347), .Z1_t (new_AGEMA_signal_15348), .Z1_f (new_AGEMA_signal_15349) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U5 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .A0_f (new_AGEMA_signal_13826), .A1_t (new_AGEMA_signal_13827), .A1_f (new_AGEMA_signal_13828), .B0_t (MixColumnsInput[58]), .B0_f (new_AGEMA_signal_13802), .B1_t (new_AGEMA_signal_13803), .B1_f (new_AGEMA_signal_13804), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n165), .Z0_f (new_AGEMA_signal_14669), .Z1_t (new_AGEMA_signal_14670), .Z1_f (new_AGEMA_signal_14671) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n129), .A0_f (new_AGEMA_signal_15350), .A1_t (new_AGEMA_signal_15351), .A1_f (new_AGEMA_signal_15352), .B0_t (MixColumnsInput[40]), .B0_f (new_AGEMA_signal_13427), .B1_t (new_AGEMA_signal_13428), .B1_f (new_AGEMA_signal_13429), .Z0_t (MixColumnsOutput[32]), .Z0_f (new_AGEMA_signal_16097), .Z1_t (new_AGEMA_signal_16098), .Z1_f (new_AGEMA_signal_16099) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n187), .A0_f (new_AGEMA_signal_14675), .A1_t (new_AGEMA_signal_14676), .A1_f (new_AGEMA_signal_14677), .B0_t (MixColumnsIns_MixOneColumnInst_2_n151), .B0_f (new_AGEMA_signal_14672), .B1_t (new_AGEMA_signal_14673), .B1_f (new_AGEMA_signal_14674), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n129), .Z0_f (new_AGEMA_signal_15350), .Z1_t (new_AGEMA_signal_15351), .Z1_f (new_AGEMA_signal_15352) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U2 ( .A0_t (MixColumnsInput[48]), .A0_f (new_AGEMA_signal_13064), .A1_t (new_AGEMA_signal_13065), .A1_f (new_AGEMA_signal_13066), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13787), .B1_t (new_AGEMA_signal_13788), .B1_f (new_AGEMA_signal_13789), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n151), .Z0_f (new_AGEMA_signal_14672), .Z1_t (new_AGEMA_signal_14673), .Z1_f (new_AGEMA_signal_14674) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U1 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13808), .A1_t (new_AGEMA_signal_13809), .A1_f (new_AGEMA_signal_13810), .B0_t (MixColumnsInput[56]), .B0_f (new_AGEMA_signal_13229), .B1_t (new_AGEMA_signal_13230), .B1_f (new_AGEMA_signal_13231), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n187), .Z0_f (new_AGEMA_signal_14675), .Z1_t (new_AGEMA_signal_14676), .Z1_f (new_AGEMA_signal_14677) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13787), .A1_t (new_AGEMA_signal_13788), .A1_f (new_AGEMA_signal_13789), .B0_t (MixColumnsInput[59]), .B0_f (new_AGEMA_signal_13799), .B1_t (new_AGEMA_signal_13800), .B1_f (new_AGEMA_signal_13801), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]), .Z0_f (new_AGEMA_signal_14678), .Z1_t (new_AGEMA_signal_14679), .Z1_f (new_AGEMA_signal_14680) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13787), .A1_t (new_AGEMA_signal_13788), .A1_f (new_AGEMA_signal_13789), .B0_t (MixColumnsInput[58]), .B0_f (new_AGEMA_signal_13802), .B1_t (new_AGEMA_signal_13803), .B1_f (new_AGEMA_signal_13804), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]), .Z0_f (new_AGEMA_signal_14681), .Z1_t (new_AGEMA_signal_14682), .Z1_f (new_AGEMA_signal_14683) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13787), .A1_t (new_AGEMA_signal_13788), .A1_f (new_AGEMA_signal_13789), .B0_t (MixColumnsInput[56]), .B0_f (new_AGEMA_signal_13229), .B1_t (new_AGEMA_signal_13230), .B1_f (new_AGEMA_signal_13231), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]), .Z0_f (new_AGEMA_signal_14684), .Z1_t (new_AGEMA_signal_14685), .Z1_f (new_AGEMA_signal_14686) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13682), .A1_t (new_AGEMA_signal_13683), .A1_f (new_AGEMA_signal_13684), .B0_t (MixColumnsInput[51]), .B0_f (new_AGEMA_signal_13694), .B1_t (new_AGEMA_signal_13695), .B1_f (new_AGEMA_signal_13696), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]), .Z0_f (new_AGEMA_signal_14687), .Z1_t (new_AGEMA_signal_14688), .Z1_f (new_AGEMA_signal_14689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13682), .A1_t (new_AGEMA_signal_13683), .A1_f (new_AGEMA_signal_13684), .B0_t (MixColumnsInput[50]), .B0_f (new_AGEMA_signal_13697), .B1_t (new_AGEMA_signal_13698), .B1_f (new_AGEMA_signal_13699), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]), .Z0_f (new_AGEMA_signal_14690), .Z1_t (new_AGEMA_signal_14691), .Z1_f (new_AGEMA_signal_14692) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13682), .A1_t (new_AGEMA_signal_13683), .A1_f (new_AGEMA_signal_13684), .B0_t (MixColumnsInput[48]), .B0_f (new_AGEMA_signal_13064), .B1_t (new_AGEMA_signal_13065), .B1_f (new_AGEMA_signal_13066), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]), .Z0_f (new_AGEMA_signal_14693), .Z1_t (new_AGEMA_signal_14694), .Z1_f (new_AGEMA_signal_14695) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13913), .A1_t (new_AGEMA_signal_13914), .A1_f (new_AGEMA_signal_13915), .B0_t (MixColumnsInput[43]), .B0_f (new_AGEMA_signal_13925), .B1_t (new_AGEMA_signal_13926), .B1_f (new_AGEMA_signal_13927), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]), .Z0_f (new_AGEMA_signal_14696), .Z1_t (new_AGEMA_signal_14697), .Z1_f (new_AGEMA_signal_14698) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13913), .A1_t (new_AGEMA_signal_13914), .A1_f (new_AGEMA_signal_13915), .B0_t (MixColumnsInput[42]), .B0_f (new_AGEMA_signal_13928), .B1_t (new_AGEMA_signal_13929), .B1_f (new_AGEMA_signal_13930), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]), .Z0_f (new_AGEMA_signal_14699), .Z1_t (new_AGEMA_signal_14700), .Z1_f (new_AGEMA_signal_14701) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13913), .A1_t (new_AGEMA_signal_13914), .A1_f (new_AGEMA_signal_13915), .B0_t (MixColumnsInput[40]), .B0_f (new_AGEMA_signal_13427), .B1_t (new_AGEMA_signal_13428), .B1_f (new_AGEMA_signal_13429), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]), .Z0_f (new_AGEMA_signal_14702), .Z1_t (new_AGEMA_signal_14703), .Z1_f (new_AGEMA_signal_14704) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13808), .A1_t (new_AGEMA_signal_13809), .A1_f (new_AGEMA_signal_13810), .B0_t (MixColumnsInput[35]), .B0_f (new_AGEMA_signal_13820), .B1_t (new_AGEMA_signal_13821), .B1_f (new_AGEMA_signal_13822), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]), .Z0_f (new_AGEMA_signal_14705), .Z1_t (new_AGEMA_signal_14706), .Z1_f (new_AGEMA_signal_14707) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13808), .A1_t (new_AGEMA_signal_13809), .A1_f (new_AGEMA_signal_13810), .B0_t (MixColumnsInput[34]), .B0_f (new_AGEMA_signal_13823), .B1_t (new_AGEMA_signal_13824), .B1_f (new_AGEMA_signal_13825), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]), .Z0_f (new_AGEMA_signal_14708), .Z1_t (new_AGEMA_signal_14709), .Z1_f (new_AGEMA_signal_14710) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13808), .A1_t (new_AGEMA_signal_13809), .A1_f (new_AGEMA_signal_13810), .B0_t (MixColumnsInput[32]), .B0_f (new_AGEMA_signal_13262), .B1_t (new_AGEMA_signal_13263), .B1_f (new_AGEMA_signal_13264), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]), .Z0_f (new_AGEMA_signal_14711), .Z1_t (new_AGEMA_signal_14712), .Z1_f (new_AGEMA_signal_14713) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U96 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n192), .A0_f (new_AGEMA_signal_16100), .A1_t (new_AGEMA_signal_16101), .A1_f (new_AGEMA_signal_16102), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13952), .B1_t (new_AGEMA_signal_13953), .B1_f (new_AGEMA_signal_13954), .Z0_t (MixColumnsOutput[9]), .Z0_f (new_AGEMA_signal_16919), .Z1_t (new_AGEMA_signal_16920), .Z1_f (new_AGEMA_signal_16921) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U95 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n191), .A0_f (new_AGEMA_signal_15416), .A1_t (new_AGEMA_signal_15417), .A1_f (new_AGEMA_signal_15418), .B0_t (MixColumnsIns_MixOneColumnInst_3_n190), .B0_f (new_AGEMA_signal_15404), .B1_t (new_AGEMA_signal_15405), .B1_f (new_AGEMA_signal_15406), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n192), .Z0_f (new_AGEMA_signal_16100), .Z1_t (new_AGEMA_signal_16101), .Z1_f (new_AGEMA_signal_16102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U94 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n189), .A0_f (new_AGEMA_signal_15353), .A1_t (new_AGEMA_signal_15354), .A1_f (new_AGEMA_signal_15355), .B0_t (MixColumnsIns_MixOneColumnInst_3_n188), .B0_f (new_AGEMA_signal_14741), .B1_t (new_AGEMA_signal_14742), .B1_f (new_AGEMA_signal_14743), .Z0_t (MixColumnsOutput[8]), .Z0_f (new_AGEMA_signal_16103), .Z1_t (new_AGEMA_signal_16104), .Z1_f (new_AGEMA_signal_16105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U93 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n187), .A0_f (new_AGEMA_signal_14771), .A1_t (new_AGEMA_signal_14772), .A1_f (new_AGEMA_signal_14773), .B0_t (MixColumnsInput[16]), .B0_f (new_AGEMA_signal_13460), .B1_t (new_AGEMA_signal_13461), .B1_f (new_AGEMA_signal_13462), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n189), .Z0_f (new_AGEMA_signal_15353), .Z1_t (new_AGEMA_signal_15354), .Z1_f (new_AGEMA_signal_15355) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U92 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n186), .A0_f (new_AGEMA_signal_15356), .A1_t (new_AGEMA_signal_15357), .A1_f (new_AGEMA_signal_15358), .B0_t (MixColumnsIns_MixOneColumnInst_3_n185), .B0_f (new_AGEMA_signal_14714), .B1_t (new_AGEMA_signal_14715), .B1_f (new_AGEMA_signal_14716), .Z0_t (MixColumnsOutput[7]), .Z0_f (new_AGEMA_signal_16106), .Z1_t (new_AGEMA_signal_16107), .Z1_f (new_AGEMA_signal_16108) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U91 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n184), .A0_f (new_AGEMA_signal_14747), .A1_t (new_AGEMA_signal_14748), .A1_f (new_AGEMA_signal_14749), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B0_f (new_AGEMA_signal_13829), .B1_t (new_AGEMA_signal_13830), .B1_f (new_AGEMA_signal_13831), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n186), .Z0_f (new_AGEMA_signal_15356), .Z1_t (new_AGEMA_signal_15357), .Z1_f (new_AGEMA_signal_15358) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U90 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n183), .A0_f (new_AGEMA_signal_15359), .A1_t (new_AGEMA_signal_15360), .A1_f (new_AGEMA_signal_15361), .B0_t (MixColumnsIns_MixOneColumnInst_3_n182), .B0_f (new_AGEMA_signal_14717), .B1_t (new_AGEMA_signal_14718), .B1_f (new_AGEMA_signal_14719), .Z0_t (MixColumnsOutput[6]), .Z0_f (new_AGEMA_signal_16109), .Z1_t (new_AGEMA_signal_16110), .Z1_f (new_AGEMA_signal_16111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U89 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n181), .A0_f (new_AGEMA_signal_14753), .A1_t (new_AGEMA_signal_14754), .A1_f (new_AGEMA_signal_14755), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13832), .B1_t (new_AGEMA_signal_13833), .B1_f (new_AGEMA_signal_13834), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n183), .Z0_f (new_AGEMA_signal_15359), .Z1_t (new_AGEMA_signal_15360), .Z1_f (new_AGEMA_signal_15361) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U88 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n180), .A0_f (new_AGEMA_signal_15362), .A1_t (new_AGEMA_signal_15363), .A1_f (new_AGEMA_signal_15364), .B0_t (MixColumnsIns_MixOneColumnInst_3_n179), .B0_f (new_AGEMA_signal_14720), .B1_t (new_AGEMA_signal_14721), .B1_f (new_AGEMA_signal_14722), .Z0_t (MixColumnsOutput[5]), .Z0_f (new_AGEMA_signal_16112), .Z1_t (new_AGEMA_signal_16113), .Z1_f (new_AGEMA_signal_16114) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U87 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n178), .A0_f (new_AGEMA_signal_14759), .A1_t (new_AGEMA_signal_14760), .A1_f (new_AGEMA_signal_14761), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13835), .B1_t (new_AGEMA_signal_13836), .B1_f (new_AGEMA_signal_13837), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n180), .Z0_f (new_AGEMA_signal_15362), .Z1_t (new_AGEMA_signal_15363), .Z1_f (new_AGEMA_signal_15364) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U86 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n177), .A0_f (new_AGEMA_signal_16115), .A1_t (new_AGEMA_signal_16116), .A1_f (new_AGEMA_signal_16117), .B0_t (MixColumnsIns_MixOneColumnInst_3_n176), .B0_f (new_AGEMA_signal_15377), .B1_t (new_AGEMA_signal_15378), .B1_f (new_AGEMA_signal_15379), .Z0_t (MixColumnsOutput[4]), .Z0_f (new_AGEMA_signal_16922), .Z1_t (new_AGEMA_signal_16923), .Z1_f (new_AGEMA_signal_16924) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U85 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n175), .A0_f (new_AGEMA_signal_15434), .A1_t (new_AGEMA_signal_15435), .A1_f (new_AGEMA_signal_15436), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13838), .B1_t (new_AGEMA_signal_13839), .B1_f (new_AGEMA_signal_13840), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n177), .Z0_f (new_AGEMA_signal_16115), .Z1_t (new_AGEMA_signal_16116), .Z1_f (new_AGEMA_signal_16117) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U84 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n174), .A0_f (new_AGEMA_signal_16118), .A1_t (new_AGEMA_signal_16119), .A1_f (new_AGEMA_signal_16120), .B0_t (MixColumnsIns_MixOneColumnInst_3_n173), .B0_f (new_AGEMA_signal_15380), .B1_t (new_AGEMA_signal_15381), .B1_f (new_AGEMA_signal_15382), .Z0_t (MixColumnsOutput[3]), .Z0_f (new_AGEMA_signal_16925), .Z1_t (new_AGEMA_signal_16926), .Z1_f (new_AGEMA_signal_16927) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U83 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n172), .A0_f (new_AGEMA_signal_15440), .A1_t (new_AGEMA_signal_15441), .A1_f (new_AGEMA_signal_15442), .B0_t (MixColumnsInput[11]), .B0_f (new_AGEMA_signal_13841), .B1_t (new_AGEMA_signal_13842), .B1_f (new_AGEMA_signal_13843), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n174), .Z0_f (new_AGEMA_signal_16118), .Z1_t (new_AGEMA_signal_16119), .Z1_f (new_AGEMA_signal_16120) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U82 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n171), .A0_f (new_AGEMA_signal_15365), .A1_t (new_AGEMA_signal_15366), .A1_f (new_AGEMA_signal_15367), .B0_t (MixColumnsIns_MixOneColumnInst_3_n185), .B0_f (new_AGEMA_signal_14714), .B1_t (new_AGEMA_signal_14715), .B1_f (new_AGEMA_signal_14716), .Z0_t (MixColumnsOutput[31]), .Z0_f (new_AGEMA_signal_16121), .Z1_t (new_AGEMA_signal_16122), .Z1_f (new_AGEMA_signal_16123) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U81 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13934), .A1_t (new_AGEMA_signal_13935), .A1_f (new_AGEMA_signal_13936), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13706), .B1_t (new_AGEMA_signal_13707), .B1_f (new_AGEMA_signal_13708), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n185), .Z0_f (new_AGEMA_signal_14714), .Z1_t (new_AGEMA_signal_14715), .Z1_f (new_AGEMA_signal_14716) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U80 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13724), .A1_t (new_AGEMA_signal_13725), .A1_f (new_AGEMA_signal_13726), .B0_t (MixColumnsIns_MixOneColumnInst_3_n170), .B0_f (new_AGEMA_signal_14726), .B1_t (new_AGEMA_signal_14727), .B1_f (new_AGEMA_signal_14728), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n171), .Z0_f (new_AGEMA_signal_15365), .Z1_t (new_AGEMA_signal_15366), .Z1_f (new_AGEMA_signal_15367) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U79 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n169), .A0_f (new_AGEMA_signal_15368), .A1_t (new_AGEMA_signal_15369), .A1_f (new_AGEMA_signal_15370), .B0_t (MixColumnsIns_MixOneColumnInst_3_n182), .B0_f (new_AGEMA_signal_14717), .B1_t (new_AGEMA_signal_14718), .B1_f (new_AGEMA_signal_14719), .Z0_t (MixColumnsOutput[30]), .Z0_f (new_AGEMA_signal_16124), .Z1_t (new_AGEMA_signal_16125), .Z1_f (new_AGEMA_signal_16126) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U78 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .A0_f (new_AGEMA_signal_13937), .A1_t (new_AGEMA_signal_13938), .A1_f (new_AGEMA_signal_13939), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13709), .B1_t (new_AGEMA_signal_13710), .B1_f (new_AGEMA_signal_13711), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n182), .Z0_f (new_AGEMA_signal_14717), .Z1_t (new_AGEMA_signal_14718), .Z1_f (new_AGEMA_signal_14719) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U77 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13727), .A1_t (new_AGEMA_signal_13728), .A1_f (new_AGEMA_signal_13729), .B0_t (MixColumnsIns_MixOneColumnInst_3_n168), .B0_f (new_AGEMA_signal_14729), .B1_t (new_AGEMA_signal_14730), .B1_f (new_AGEMA_signal_14731), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n169), .Z0_f (new_AGEMA_signal_15368), .Z1_t (new_AGEMA_signal_15369), .Z1_f (new_AGEMA_signal_15370) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U76 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n167), .A0_f (new_AGEMA_signal_15371), .A1_t (new_AGEMA_signal_15372), .A1_f (new_AGEMA_signal_15373), .B0_t (MixColumnsIns_MixOneColumnInst_3_n166), .B0_f (new_AGEMA_signal_14723), .B1_t (new_AGEMA_signal_14724), .B1_f (new_AGEMA_signal_14725), .Z0_t (MixColumnsOutput[2]), .Z0_f (new_AGEMA_signal_16127), .Z1_t (new_AGEMA_signal_16128), .Z1_f (new_AGEMA_signal_16129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U75 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n165), .A0_f (new_AGEMA_signal_14765), .A1_t (new_AGEMA_signal_14766), .A1_f (new_AGEMA_signal_14767), .B0_t (MixColumnsInput[10]), .B0_f (new_AGEMA_signal_13844), .B1_t (new_AGEMA_signal_13845), .B1_f (new_AGEMA_signal_13846), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n167), .Z0_f (new_AGEMA_signal_15371), .Z1_t (new_AGEMA_signal_15372), .Z1_f (new_AGEMA_signal_15373) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U74 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n164), .A0_f (new_AGEMA_signal_15374), .A1_t (new_AGEMA_signal_15375), .A1_f (new_AGEMA_signal_15376), .B0_t (MixColumnsIns_MixOneColumnInst_3_n179), .B0_f (new_AGEMA_signal_14720), .B1_t (new_AGEMA_signal_14721), .B1_f (new_AGEMA_signal_14722), .Z0_t (MixColumnsOutput[29]), .Z0_f (new_AGEMA_signal_16130), .Z1_t (new_AGEMA_signal_16131), .Z1_f (new_AGEMA_signal_16132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U73 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .A0_f (new_AGEMA_signal_13940), .A1_t (new_AGEMA_signal_13941), .A1_f (new_AGEMA_signal_13942), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13712), .B1_t (new_AGEMA_signal_13713), .B1_f (new_AGEMA_signal_13714), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n179), .Z0_f (new_AGEMA_signal_14720), .Z1_t (new_AGEMA_signal_14721), .Z1_f (new_AGEMA_signal_14722) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U72 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13730), .A1_t (new_AGEMA_signal_13731), .A1_f (new_AGEMA_signal_13732), .B0_t (MixColumnsIns_MixOneColumnInst_3_n163), .B0_f (new_AGEMA_signal_14732), .B1_t (new_AGEMA_signal_14733), .B1_f (new_AGEMA_signal_14734), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n164), .Z0_f (new_AGEMA_signal_15374), .Z1_t (new_AGEMA_signal_15375), .Z1_f (new_AGEMA_signal_15376) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U71 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n162), .A0_f (new_AGEMA_signal_16133), .A1_t (new_AGEMA_signal_16134), .A1_f (new_AGEMA_signal_16135), .B0_t (MixColumnsIns_MixOneColumnInst_3_n176), .B0_f (new_AGEMA_signal_15377), .B1_t (new_AGEMA_signal_15378), .B1_f (new_AGEMA_signal_15379), .Z0_t (MixColumnsOutput[28]), .Z0_f (new_AGEMA_signal_16928), .Z1_t (new_AGEMA_signal_16929), .Z1_f (new_AGEMA_signal_16930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U70 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .A0_f (new_AGEMA_signal_13943), .A1_t (new_AGEMA_signal_13944), .A1_f (new_AGEMA_signal_13945), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]), .B0_f (new_AGEMA_signal_14774), .B1_t (new_AGEMA_signal_14775), .B1_f (new_AGEMA_signal_14776), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n176), .Z0_f (new_AGEMA_signal_15377), .Z1_t (new_AGEMA_signal_15378), .Z1_f (new_AGEMA_signal_15379) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U69 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13733), .A1_t (new_AGEMA_signal_13734), .A1_f (new_AGEMA_signal_13735), .B0_t (MixColumnsIns_MixOneColumnInst_3_n161), .B0_f (new_AGEMA_signal_15398), .B1_t (new_AGEMA_signal_15399), .B1_f (new_AGEMA_signal_15400), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n162), .Z0_f (new_AGEMA_signal_16133), .Z1_t (new_AGEMA_signal_16134), .Z1_f (new_AGEMA_signal_16135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U68 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n160), .A0_f (new_AGEMA_signal_16136), .A1_t (new_AGEMA_signal_16137), .A1_f (new_AGEMA_signal_16138), .B0_t (MixColumnsIns_MixOneColumnInst_3_n173), .B0_f (new_AGEMA_signal_15380), .B1_t (new_AGEMA_signal_15381), .B1_f (new_AGEMA_signal_15382), .Z0_t (MixColumnsOutput[27]), .Z0_f (new_AGEMA_signal_16931), .Z1_t (new_AGEMA_signal_16932), .Z1_f (new_AGEMA_signal_16933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U67 ( .A0_t (MixColumnsInput[19]), .A0_f (new_AGEMA_signal_13946), .A1_t (new_AGEMA_signal_13947), .A1_f (new_AGEMA_signal_13948), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]), .B0_f (new_AGEMA_signal_14777), .B1_t (new_AGEMA_signal_14778), .B1_f (new_AGEMA_signal_14779), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n173), .Z0_f (new_AGEMA_signal_15380), .Z1_t (new_AGEMA_signal_15381), .Z1_f (new_AGEMA_signal_15382) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U66 ( .A0_t (MixColumnsInput[3]), .A0_f (new_AGEMA_signal_13736), .A1_t (new_AGEMA_signal_13737), .A1_f (new_AGEMA_signal_13738), .B0_t (MixColumnsIns_MixOneColumnInst_3_n159), .B0_f (new_AGEMA_signal_15407), .B1_t (new_AGEMA_signal_15408), .B1_f (new_AGEMA_signal_15409), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n160), .Z0_f (new_AGEMA_signal_16136), .Z1_t (new_AGEMA_signal_16137), .Z1_f (new_AGEMA_signal_16138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U65 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n158), .A0_f (new_AGEMA_signal_15383), .A1_t (new_AGEMA_signal_15384), .A1_f (new_AGEMA_signal_15385), .B0_t (MixColumnsIns_MixOneColumnInst_3_n166), .B0_f (new_AGEMA_signal_14723), .B1_t (new_AGEMA_signal_14724), .B1_f (new_AGEMA_signal_14725), .Z0_t (MixColumnsOutput[26]), .Z0_f (new_AGEMA_signal_16139), .Z1_t (new_AGEMA_signal_16140), .Z1_f (new_AGEMA_signal_16141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U64 ( .A0_t (MixColumnsInput[18]), .A0_f (new_AGEMA_signal_13949), .A1_t (new_AGEMA_signal_13950), .A1_f (new_AGEMA_signal_13951), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13721), .B1_t (new_AGEMA_signal_13722), .B1_f (new_AGEMA_signal_13723), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n166), .Z0_f (new_AGEMA_signal_14723), .Z1_t (new_AGEMA_signal_14724), .Z1_f (new_AGEMA_signal_14725) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U63 ( .A0_t (MixColumnsInput[2]), .A0_f (new_AGEMA_signal_13739), .A1_t (new_AGEMA_signal_13740), .A1_f (new_AGEMA_signal_13741), .B0_t (MixColumnsIns_MixOneColumnInst_3_n157), .B0_f (new_AGEMA_signal_14735), .B1_t (new_AGEMA_signal_14736), .B1_f (new_AGEMA_signal_14737), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n158), .Z0_f (new_AGEMA_signal_15383), .Z1_t (new_AGEMA_signal_15384), .Z1_f (new_AGEMA_signal_15385) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U62 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n156), .A0_f (new_AGEMA_signal_16142), .A1_t (new_AGEMA_signal_16143), .A1_f (new_AGEMA_signal_16144), .B0_t (MixColumnsIns_MixOneColumnInst_3_n155), .B0_f (new_AGEMA_signal_15401), .B1_t (new_AGEMA_signal_15402), .B1_f (new_AGEMA_signal_15403), .Z0_t (MixColumnsOutput[25]), .Z0_f (new_AGEMA_signal_16934), .Z1_t (new_AGEMA_signal_16935), .Z1_f (new_AGEMA_signal_16936) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U61 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .A0_f (new_AGEMA_signal_13742), .A1_t (new_AGEMA_signal_13743), .A1_f (new_AGEMA_signal_13744), .B0_t (MixColumnsIns_MixOneColumnInst_3_n154), .B0_f (new_AGEMA_signal_15413), .B1_t (new_AGEMA_signal_15414), .B1_f (new_AGEMA_signal_15415), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n156), .Z0_f (new_AGEMA_signal_16142), .Z1_t (new_AGEMA_signal_16143), .Z1_f (new_AGEMA_signal_16144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U60 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n153), .A0_f (new_AGEMA_signal_15386), .A1_t (new_AGEMA_signal_15387), .A1_f (new_AGEMA_signal_15388), .B0_t (MixColumnsIns_MixOneColumnInst_3_n152), .B0_f (new_AGEMA_signal_14738), .B1_t (new_AGEMA_signal_14739), .B1_f (new_AGEMA_signal_14740), .Z0_t (MixColumnsOutput[24]), .Z0_f (new_AGEMA_signal_16145), .Z1_t (new_AGEMA_signal_16146), .Z1_f (new_AGEMA_signal_16147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U59 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n151), .A0_f (new_AGEMA_signal_14768), .A1_t (new_AGEMA_signal_14769), .A1_f (new_AGEMA_signal_14770), .B0_t (MixColumnsInput[0]), .B0_f (new_AGEMA_signal_13130), .B1_t (new_AGEMA_signal_13131), .B1_f (new_AGEMA_signal_13132), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n153), .Z0_f (new_AGEMA_signal_15386), .Z1_t (new_AGEMA_signal_15387), .Z1_f (new_AGEMA_signal_15388) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U58 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n150), .A0_f (new_AGEMA_signal_15389), .A1_t (new_AGEMA_signal_15390), .A1_f (new_AGEMA_signal_15391), .B0_t (MixColumnsIns_MixOneColumnInst_3_n170), .B0_f (new_AGEMA_signal_14726), .B1_t (new_AGEMA_signal_14727), .B1_f (new_AGEMA_signal_14728), .Z0_t (MixColumnsOutput[23]), .Z0_f (new_AGEMA_signal_16148), .Z1_t (new_AGEMA_signal_16149), .Z1_f (new_AGEMA_signal_16150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U57 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13829), .A1_t (new_AGEMA_signal_13830), .A1_f (new_AGEMA_signal_13831), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13937), .B1_t (new_AGEMA_signal_13938), .B1_f (new_AGEMA_signal_13939), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n170), .Z0_f (new_AGEMA_signal_14726), .Z1_t (new_AGEMA_signal_14727), .Z1_f (new_AGEMA_signal_14728) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U56 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13703), .A1_t (new_AGEMA_signal_13704), .A1_f (new_AGEMA_signal_13705), .B0_t (MixColumnsIns_MixOneColumnInst_3_n149), .B0_f (new_AGEMA_signal_14744), .B1_t (new_AGEMA_signal_14745), .B1_f (new_AGEMA_signal_14746), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n150), .Z0_f (new_AGEMA_signal_15389), .Z1_t (new_AGEMA_signal_15390), .Z1_f (new_AGEMA_signal_15391) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U55 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n148), .A0_f (new_AGEMA_signal_15392), .A1_t (new_AGEMA_signal_15393), .A1_f (new_AGEMA_signal_15394), .B0_t (MixColumnsIns_MixOneColumnInst_3_n168), .B0_f (new_AGEMA_signal_14729), .B1_t (new_AGEMA_signal_14730), .B1_f (new_AGEMA_signal_14731), .Z0_t (MixColumnsOutput[22]), .Z0_f (new_AGEMA_signal_16151), .Z1_t (new_AGEMA_signal_16152), .Z1_f (new_AGEMA_signal_16153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U54 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .A0_f (new_AGEMA_signal_13832), .A1_t (new_AGEMA_signal_13833), .A1_f (new_AGEMA_signal_13834), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13940), .B1_t (new_AGEMA_signal_13941), .B1_f (new_AGEMA_signal_13942), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n168), .Z0_f (new_AGEMA_signal_14729), .Z1_t (new_AGEMA_signal_14730), .Z1_f (new_AGEMA_signal_14731) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U53 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .A0_f (new_AGEMA_signal_13706), .A1_t (new_AGEMA_signal_13707), .A1_f (new_AGEMA_signal_13708), .B0_t (MixColumnsIns_MixOneColumnInst_3_n147), .B0_f (new_AGEMA_signal_14750), .B1_t (new_AGEMA_signal_14751), .B1_f (new_AGEMA_signal_14752), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n148), .Z0_f (new_AGEMA_signal_15392), .Z1_t (new_AGEMA_signal_15393), .Z1_f (new_AGEMA_signal_15394) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U52 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n146), .A0_f (new_AGEMA_signal_15395), .A1_t (new_AGEMA_signal_15396), .A1_f (new_AGEMA_signal_15397), .B0_t (MixColumnsIns_MixOneColumnInst_3_n163), .B0_f (new_AGEMA_signal_14732), .B1_t (new_AGEMA_signal_14733), .B1_f (new_AGEMA_signal_14734), .Z0_t (MixColumnsOutput[21]), .Z0_f (new_AGEMA_signal_16154), .Z1_t (new_AGEMA_signal_16155), .Z1_f (new_AGEMA_signal_16156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U51 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .A0_f (new_AGEMA_signal_13835), .A1_t (new_AGEMA_signal_13836), .A1_f (new_AGEMA_signal_13837), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13943), .B1_t (new_AGEMA_signal_13944), .B1_f (new_AGEMA_signal_13945), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n163), .Z0_f (new_AGEMA_signal_14732), .Z1_t (new_AGEMA_signal_14733), .Z1_f (new_AGEMA_signal_14734) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U50 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .A0_f (new_AGEMA_signal_13709), .A1_t (new_AGEMA_signal_13710), .A1_f (new_AGEMA_signal_13711), .B0_t (MixColumnsIns_MixOneColumnInst_3_n145), .B0_f (new_AGEMA_signal_14756), .B1_t (new_AGEMA_signal_14757), .B1_f (new_AGEMA_signal_14758), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n146), .Z0_f (new_AGEMA_signal_15395), .Z1_t (new_AGEMA_signal_15396), .Z1_f (new_AGEMA_signal_15397) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U49 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n144), .A0_f (new_AGEMA_signal_16157), .A1_t (new_AGEMA_signal_16158), .A1_f (new_AGEMA_signal_16159), .B0_t (MixColumnsIns_MixOneColumnInst_3_n161), .B0_f (new_AGEMA_signal_15398), .B1_t (new_AGEMA_signal_15399), .B1_f (new_AGEMA_signal_15400), .Z0_t (MixColumnsOutput[20]), .Z0_f (new_AGEMA_signal_16937), .Z1_t (new_AGEMA_signal_16938), .Z1_f (new_AGEMA_signal_16939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U48 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .A0_f (new_AGEMA_signal_13838), .A1_t (new_AGEMA_signal_13839), .A1_f (new_AGEMA_signal_13840), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]), .B0_f (new_AGEMA_signal_14783), .B1_t (new_AGEMA_signal_14784), .B1_f (new_AGEMA_signal_14785), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n161), .Z0_f (new_AGEMA_signal_15398), .Z1_t (new_AGEMA_signal_15399), .Z1_f (new_AGEMA_signal_15400) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U47 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .A0_f (new_AGEMA_signal_13712), .A1_t (new_AGEMA_signal_13713), .A1_f (new_AGEMA_signal_13714), .B0_t (MixColumnsIns_MixOneColumnInst_3_n143), .B0_f (new_AGEMA_signal_15431), .B1_t (new_AGEMA_signal_15432), .B1_f (new_AGEMA_signal_15433), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n144), .Z0_f (new_AGEMA_signal_16157), .Z1_t (new_AGEMA_signal_16158), .Z1_f (new_AGEMA_signal_16159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U46 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n142), .A0_f (new_AGEMA_signal_16160), .A1_t (new_AGEMA_signal_16161), .A1_f (new_AGEMA_signal_16162), .B0_t (MixColumnsIns_MixOneColumnInst_3_n155), .B0_f (new_AGEMA_signal_15401), .B1_t (new_AGEMA_signal_15402), .B1_f (new_AGEMA_signal_15403), .Z0_t (MixColumnsOutput[1]), .Z0_f (new_AGEMA_signal_16940), .Z1_t (new_AGEMA_signal_16941), .Z1_f (new_AGEMA_signal_16942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U45 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .A0_f (new_AGEMA_signal_13952), .A1_t (new_AGEMA_signal_13953), .A1_f (new_AGEMA_signal_13954), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]), .B0_f (new_AGEMA_signal_14780), .B1_t (new_AGEMA_signal_14781), .B1_f (new_AGEMA_signal_14782), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n155), .Z0_f (new_AGEMA_signal_15401), .Z1_t (new_AGEMA_signal_15402), .Z1_f (new_AGEMA_signal_15403) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U44 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .A0_f (new_AGEMA_signal_13847), .A1_t (new_AGEMA_signal_13848), .A1_f (new_AGEMA_signal_13849), .B0_t (MixColumnsIns_MixOneColumnInst_3_n190), .B0_f (new_AGEMA_signal_15404), .B1_t (new_AGEMA_signal_15405), .B1_f (new_AGEMA_signal_15406), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n142), .Z0_f (new_AGEMA_signal_16160), .Z1_t (new_AGEMA_signal_16161), .Z1_f (new_AGEMA_signal_16162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U43 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .A0_f (new_AGEMA_signal_13721), .A1_t (new_AGEMA_signal_13722), .A1_f (new_AGEMA_signal_13723), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]), .B0_f (new_AGEMA_signal_14807), .B1_t (new_AGEMA_signal_14808), .B1_f (new_AGEMA_signal_14809), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n190), .Z0_f (new_AGEMA_signal_15404), .Z1_t (new_AGEMA_signal_15405), .Z1_f (new_AGEMA_signal_15406) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U42 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n141), .A0_f (new_AGEMA_signal_16163), .A1_t (new_AGEMA_signal_16164), .A1_f (new_AGEMA_signal_16165), .B0_t (MixColumnsIns_MixOneColumnInst_3_n159), .B0_f (new_AGEMA_signal_15407), .B1_t (new_AGEMA_signal_15408), .B1_f (new_AGEMA_signal_15409), .Z0_t (MixColumnsOutput[19]), .Z0_f (new_AGEMA_signal_16943), .Z1_t (new_AGEMA_signal_16944), .Z1_f (new_AGEMA_signal_16945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U41 ( .A0_t (MixColumnsInput[11]), .A0_f (new_AGEMA_signal_13841), .A1_t (new_AGEMA_signal_13842), .A1_f (new_AGEMA_signal_13843), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]), .B0_f (new_AGEMA_signal_14786), .B1_t (new_AGEMA_signal_14787), .B1_f (new_AGEMA_signal_14788), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n159), .Z0_f (new_AGEMA_signal_15407), .Z1_t (new_AGEMA_signal_15408), .Z1_f (new_AGEMA_signal_15409) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U40 ( .A0_t (MixColumnsInput[27]), .A0_f (new_AGEMA_signal_13715), .A1_t (new_AGEMA_signal_13716), .A1_f (new_AGEMA_signal_13717), .B0_t (MixColumnsIns_MixOneColumnInst_3_n140), .B0_f (new_AGEMA_signal_15437), .B1_t (new_AGEMA_signal_15438), .B1_f (new_AGEMA_signal_15439), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n141), .Z0_f (new_AGEMA_signal_16163), .Z1_t (new_AGEMA_signal_16164), .Z1_f (new_AGEMA_signal_16165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U39 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n139), .A0_f (new_AGEMA_signal_15410), .A1_t (new_AGEMA_signal_15411), .A1_f (new_AGEMA_signal_15412), .B0_t (MixColumnsIns_MixOneColumnInst_3_n157), .B0_f (new_AGEMA_signal_14735), .B1_t (new_AGEMA_signal_14736), .B1_f (new_AGEMA_signal_14737), .Z0_t (MixColumnsOutput[18]), .Z0_f (new_AGEMA_signal_16166), .Z1_t (new_AGEMA_signal_16167), .Z1_f (new_AGEMA_signal_16168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U38 ( .A0_t (MixColumnsInput[10]), .A0_f (new_AGEMA_signal_13844), .A1_t (new_AGEMA_signal_13845), .A1_f (new_AGEMA_signal_13846), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .B0_f (new_AGEMA_signal_13952), .B1_t (new_AGEMA_signal_13953), .B1_f (new_AGEMA_signal_13954), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n157), .Z0_f (new_AGEMA_signal_14735), .Z1_t (new_AGEMA_signal_14736), .Z1_f (new_AGEMA_signal_14737) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U37 ( .A0_t (MixColumnsInput[26]), .A0_f (new_AGEMA_signal_13718), .A1_t (new_AGEMA_signal_13719), .A1_f (new_AGEMA_signal_13720), .B0_t (MixColumnsIns_MixOneColumnInst_3_n138), .B0_f (new_AGEMA_signal_14762), .B1_t (new_AGEMA_signal_14763), .B1_f (new_AGEMA_signal_14764), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n139), .Z0_f (new_AGEMA_signal_15410), .Z1_t (new_AGEMA_signal_15411), .Z1_f (new_AGEMA_signal_15412) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U36 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n137), .A0_f (new_AGEMA_signal_16169), .A1_t (new_AGEMA_signal_16170), .A1_f (new_AGEMA_signal_16171), .B0_t (MixColumnsIns_MixOneColumnInst_3_n154), .B0_f (new_AGEMA_signal_15413), .B1_t (new_AGEMA_signal_15414), .B1_f (new_AGEMA_signal_15415), .Z0_t (MixColumnsOutput[17]), .Z0_f (new_AGEMA_signal_16946), .Z1_t (new_AGEMA_signal_16947), .Z1_f (new_AGEMA_signal_16948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U35 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]), .A0_f (new_AGEMA_signal_14789), .A1_t (new_AGEMA_signal_14790), .A1_f (new_AGEMA_signal_14791), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13847), .B1_t (new_AGEMA_signal_13848), .B1_f (new_AGEMA_signal_13849), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n154), .Z0_f (new_AGEMA_signal_15413), .Z1_t (new_AGEMA_signal_15414), .Z1_f (new_AGEMA_signal_15415) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U34 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n191), .A0_f (new_AGEMA_signal_15416), .A1_t (new_AGEMA_signal_15417), .A1_f (new_AGEMA_signal_15418), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .B0_f (new_AGEMA_signal_13721), .B1_t (new_AGEMA_signal_13722), .B1_f (new_AGEMA_signal_13723), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n137), .Z0_f (new_AGEMA_signal_16169), .Z1_t (new_AGEMA_signal_16170), .Z1_f (new_AGEMA_signal_16171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U33 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]), .A0_f (new_AGEMA_signal_14798), .A1_t (new_AGEMA_signal_14799), .A1_f (new_AGEMA_signal_14800), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .B0_f (new_AGEMA_signal_13742), .B1_t (new_AGEMA_signal_13743), .B1_f (new_AGEMA_signal_13744), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n191), .Z0_f (new_AGEMA_signal_15416), .Z1_t (new_AGEMA_signal_15417), .Z1_f (new_AGEMA_signal_15418) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U32 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n136), .A0_f (new_AGEMA_signal_15419), .A1_t (new_AGEMA_signal_15420), .A1_f (new_AGEMA_signal_15421), .B0_t (MixColumnsIns_MixOneColumnInst_3_n152), .B0_f (new_AGEMA_signal_14738), .B1_t (new_AGEMA_signal_14739), .B1_f (new_AGEMA_signal_14740), .Z0_t (MixColumnsOutput[16]), .Z0_f (new_AGEMA_signal_16172), .Z1_t (new_AGEMA_signal_16173), .Z1_f (new_AGEMA_signal_16174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U31 ( .A0_t (MixColumnsInput[8]), .A0_f (new_AGEMA_signal_13295), .A1_t (new_AGEMA_signal_13296), .A1_f (new_AGEMA_signal_13297), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13934), .B1_t (new_AGEMA_signal_13935), .B1_f (new_AGEMA_signal_13936), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n152), .Z0_f (new_AGEMA_signal_14738), .Z1_t (new_AGEMA_signal_14739), .Z1_f (new_AGEMA_signal_14740) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U30 ( .A0_t (MixColumnsInput[24]), .A0_f (new_AGEMA_signal_13097), .A1_t (new_AGEMA_signal_13098), .A1_f (new_AGEMA_signal_13099), .B0_t (MixColumnsIns_MixOneColumnInst_3_n188), .B0_f (new_AGEMA_signal_14741), .B1_t (new_AGEMA_signal_14742), .B1_f (new_AGEMA_signal_14743), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n136), .Z0_f (new_AGEMA_signal_15419), .Z1_t (new_AGEMA_signal_15420), .Z1_f (new_AGEMA_signal_15421) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U29 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13829), .A1_t (new_AGEMA_signal_13830), .A1_f (new_AGEMA_signal_13831), .B0_t (MixColumnsInput[0]), .B0_f (new_AGEMA_signal_13130), .B1_t (new_AGEMA_signal_13131), .B1_f (new_AGEMA_signal_13132), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n188), .Z0_f (new_AGEMA_signal_14741), .Z1_t (new_AGEMA_signal_14742), .Z1_f (new_AGEMA_signal_14743) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U28 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n135), .A0_f (new_AGEMA_signal_15422), .A1_t (new_AGEMA_signal_15423), .A1_f (new_AGEMA_signal_15424), .B0_t (MixColumnsIns_MixOneColumnInst_3_n149), .B0_f (new_AGEMA_signal_14744), .B1_t (new_AGEMA_signal_14745), .B1_f (new_AGEMA_signal_14746), .Z0_t (MixColumnsOutput[15]), .Z0_f (new_AGEMA_signal_16175), .Z1_t (new_AGEMA_signal_16176), .Z1_f (new_AGEMA_signal_16177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U27 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13724), .A1_t (new_AGEMA_signal_13725), .A1_f (new_AGEMA_signal_13726), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .B0_f (new_AGEMA_signal_13832), .B1_t (new_AGEMA_signal_13833), .B1_f (new_AGEMA_signal_13834), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n149), .Z0_f (new_AGEMA_signal_14744), .Z1_t (new_AGEMA_signal_14745), .Z1_f (new_AGEMA_signal_14746) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U26 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n184), .A0_f (new_AGEMA_signal_14747), .A1_t (new_AGEMA_signal_14748), .A1_f (new_AGEMA_signal_14749), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B0_f (new_AGEMA_signal_13934), .B1_t (new_AGEMA_signal_13935), .B1_f (new_AGEMA_signal_13936), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n135), .Z0_f (new_AGEMA_signal_15422), .Z1_t (new_AGEMA_signal_15423), .Z1_f (new_AGEMA_signal_15424) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U25 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13727), .A1_t (new_AGEMA_signal_13728), .A1_f (new_AGEMA_signal_13729), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13703), .B1_t (new_AGEMA_signal_13704), .B1_f (new_AGEMA_signal_13705), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n184), .Z0_f (new_AGEMA_signal_14747), .Z1_t (new_AGEMA_signal_14748), .Z1_f (new_AGEMA_signal_14749) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U24 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n134), .A0_f (new_AGEMA_signal_15425), .A1_t (new_AGEMA_signal_15426), .A1_f (new_AGEMA_signal_15427), .B0_t (MixColumnsIns_MixOneColumnInst_3_n147), .B0_f (new_AGEMA_signal_14750), .B1_t (new_AGEMA_signal_14751), .B1_f (new_AGEMA_signal_14752), .Z0_t (MixColumnsOutput[14]), .Z0_f (new_AGEMA_signal_16178), .Z1_t (new_AGEMA_signal_16179), .Z1_f (new_AGEMA_signal_16180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U23 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .A0_f (new_AGEMA_signal_13727), .A1_t (new_AGEMA_signal_13728), .A1_f (new_AGEMA_signal_13729), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .B0_f (new_AGEMA_signal_13835), .B1_t (new_AGEMA_signal_13836), .B1_f (new_AGEMA_signal_13837), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n147), .Z0_f (new_AGEMA_signal_14750), .Z1_t (new_AGEMA_signal_14751), .Z1_f (new_AGEMA_signal_14752) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U22 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n181), .A0_f (new_AGEMA_signal_14753), .A1_t (new_AGEMA_signal_14754), .A1_f (new_AGEMA_signal_14755), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .B0_f (new_AGEMA_signal_13937), .B1_t (new_AGEMA_signal_13938), .B1_f (new_AGEMA_signal_13939), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n134), .Z0_f (new_AGEMA_signal_15425), .Z1_t (new_AGEMA_signal_15426), .Z1_f (new_AGEMA_signal_15427) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U21 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13730), .A1_t (new_AGEMA_signal_13731), .A1_f (new_AGEMA_signal_13732), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .B0_f (new_AGEMA_signal_13706), .B1_t (new_AGEMA_signal_13707), .B1_f (new_AGEMA_signal_13708), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n181), .Z0_f (new_AGEMA_signal_14753), .Z1_t (new_AGEMA_signal_14754), .Z1_f (new_AGEMA_signal_14755) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U20 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n133), .A0_f (new_AGEMA_signal_15428), .A1_t (new_AGEMA_signal_15429), .A1_f (new_AGEMA_signal_15430), .B0_t (MixColumnsIns_MixOneColumnInst_3_n145), .B0_f (new_AGEMA_signal_14756), .B1_t (new_AGEMA_signal_14757), .B1_f (new_AGEMA_signal_14758), .Z0_t (MixColumnsOutput[13]), .Z0_f (new_AGEMA_signal_16181), .Z1_t (new_AGEMA_signal_16182), .Z1_f (new_AGEMA_signal_16183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U19 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .A0_f (new_AGEMA_signal_13730), .A1_t (new_AGEMA_signal_13731), .A1_f (new_AGEMA_signal_13732), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .B0_f (new_AGEMA_signal_13838), .B1_t (new_AGEMA_signal_13839), .B1_f (new_AGEMA_signal_13840), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n145), .Z0_f (new_AGEMA_signal_14756), .Z1_t (new_AGEMA_signal_14757), .Z1_f (new_AGEMA_signal_14758) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U18 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n178), .A0_f (new_AGEMA_signal_14759), .A1_t (new_AGEMA_signal_14760), .A1_f (new_AGEMA_signal_14761), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .B0_f (new_AGEMA_signal_13940), .B1_t (new_AGEMA_signal_13941), .B1_f (new_AGEMA_signal_13942), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n133), .Z0_f (new_AGEMA_signal_15428), .Z1_t (new_AGEMA_signal_15429), .Z1_f (new_AGEMA_signal_15430) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U17 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13733), .A1_t (new_AGEMA_signal_13734), .A1_f (new_AGEMA_signal_13735), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .B0_f (new_AGEMA_signal_13709), .B1_t (new_AGEMA_signal_13710), .B1_f (new_AGEMA_signal_13711), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n178), .Z0_f (new_AGEMA_signal_14759), .Z1_t (new_AGEMA_signal_14760), .Z1_f (new_AGEMA_signal_14761) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U16 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n132), .A0_f (new_AGEMA_signal_16184), .A1_t (new_AGEMA_signal_16185), .A1_f (new_AGEMA_signal_16186), .B0_t (MixColumnsIns_MixOneColumnInst_3_n143), .B0_f (new_AGEMA_signal_15431), .B1_t (new_AGEMA_signal_15432), .B1_f (new_AGEMA_signal_15433), .Z0_t (MixColumnsOutput[12]), .Z0_f (new_AGEMA_signal_16949), .Z1_t (new_AGEMA_signal_16950), .Z1_f (new_AGEMA_signal_16951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U15 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .A0_f (new_AGEMA_signal_13733), .A1_t (new_AGEMA_signal_13734), .A1_f (new_AGEMA_signal_13735), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]), .B0_f (new_AGEMA_signal_14792), .B1_t (new_AGEMA_signal_14793), .B1_f (new_AGEMA_signal_14794), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n143), .Z0_f (new_AGEMA_signal_15431), .Z1_t (new_AGEMA_signal_15432), .Z1_f (new_AGEMA_signal_15433) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U14 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n175), .A0_f (new_AGEMA_signal_15434), .A1_t (new_AGEMA_signal_15435), .A1_f (new_AGEMA_signal_15436), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .B0_f (new_AGEMA_signal_13943), .B1_t (new_AGEMA_signal_13944), .B1_f (new_AGEMA_signal_13945), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n132), .Z0_f (new_AGEMA_signal_16184), .Z1_t (new_AGEMA_signal_16185), .Z1_f (new_AGEMA_signal_16186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U13 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]), .A0_f (new_AGEMA_signal_14801), .A1_t (new_AGEMA_signal_14802), .A1_f (new_AGEMA_signal_14803), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .B0_f (new_AGEMA_signal_13712), .B1_t (new_AGEMA_signal_13713), .B1_f (new_AGEMA_signal_13714), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n175), .Z0_f (new_AGEMA_signal_15434), .Z1_t (new_AGEMA_signal_15435), .Z1_f (new_AGEMA_signal_15436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U12 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n131), .A0_f (new_AGEMA_signal_16187), .A1_t (new_AGEMA_signal_16188), .A1_f (new_AGEMA_signal_16189), .B0_t (MixColumnsIns_MixOneColumnInst_3_n140), .B0_f (new_AGEMA_signal_15437), .B1_t (new_AGEMA_signal_15438), .B1_f (new_AGEMA_signal_15439), .Z0_t (MixColumnsOutput[11]), .Z0_f (new_AGEMA_signal_16952), .Z1_t (new_AGEMA_signal_16953), .Z1_f (new_AGEMA_signal_16954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U11 ( .A0_t (MixColumnsInput[3]), .A0_f (new_AGEMA_signal_13736), .A1_t (new_AGEMA_signal_13737), .A1_f (new_AGEMA_signal_13738), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]), .B0_f (new_AGEMA_signal_14795), .B1_t (new_AGEMA_signal_14796), .B1_f (new_AGEMA_signal_14797), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n140), .Z0_f (new_AGEMA_signal_15437), .Z1_t (new_AGEMA_signal_15438), .Z1_f (new_AGEMA_signal_15439) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U10 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n172), .A0_f (new_AGEMA_signal_15440), .A1_t (new_AGEMA_signal_15441), .A1_f (new_AGEMA_signal_15442), .B0_t (MixColumnsInput[19]), .B0_f (new_AGEMA_signal_13946), .B1_t (new_AGEMA_signal_13947), .B1_f (new_AGEMA_signal_13948), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n131), .Z0_f (new_AGEMA_signal_16187), .Z1_t (new_AGEMA_signal_16188), .Z1_f (new_AGEMA_signal_16189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U9 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]), .A0_f (new_AGEMA_signal_14804), .A1_t (new_AGEMA_signal_14805), .A1_f (new_AGEMA_signal_14806), .B0_t (MixColumnsInput[27]), .B0_f (new_AGEMA_signal_13715), .B1_t (new_AGEMA_signal_13716), .B1_f (new_AGEMA_signal_13717), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n172), .Z0_f (new_AGEMA_signal_15440), .Z1_t (new_AGEMA_signal_15441), .Z1_f (new_AGEMA_signal_15442) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U8 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n130), .A0_f (new_AGEMA_signal_15443), .A1_t (new_AGEMA_signal_15444), .A1_f (new_AGEMA_signal_15445), .B0_t (MixColumnsIns_MixOneColumnInst_3_n138), .B0_f (new_AGEMA_signal_14762), .B1_t (new_AGEMA_signal_14763), .B1_f (new_AGEMA_signal_14764), .Z0_t (MixColumnsOutput[10]), .Z0_f (new_AGEMA_signal_16190), .Z1_t (new_AGEMA_signal_16191), .Z1_f (new_AGEMA_signal_16192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U7 ( .A0_t (MixColumnsInput[2]), .A0_f (new_AGEMA_signal_13739), .A1_t (new_AGEMA_signal_13740), .A1_f (new_AGEMA_signal_13741), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .B0_f (new_AGEMA_signal_13847), .B1_t (new_AGEMA_signal_13848), .B1_f (new_AGEMA_signal_13849), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n138), .Z0_f (new_AGEMA_signal_14762), .Z1_t (new_AGEMA_signal_14763), .Z1_f (new_AGEMA_signal_14764) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U6 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n165), .A0_f (new_AGEMA_signal_14765), .A1_t (new_AGEMA_signal_14766), .A1_f (new_AGEMA_signal_14767), .B0_t (MixColumnsInput[18]), .B0_f (new_AGEMA_signal_13949), .B1_t (new_AGEMA_signal_13950), .B1_f (new_AGEMA_signal_13951), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n130), .Z0_f (new_AGEMA_signal_15443), .Z1_t (new_AGEMA_signal_15444), .Z1_f (new_AGEMA_signal_15445) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U5 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .A0_f (new_AGEMA_signal_13742), .A1_t (new_AGEMA_signal_13743), .A1_f (new_AGEMA_signal_13744), .B0_t (MixColumnsInput[26]), .B0_f (new_AGEMA_signal_13718), .B1_t (new_AGEMA_signal_13719), .B1_f (new_AGEMA_signal_13720), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n165), .Z0_f (new_AGEMA_signal_14765), .Z1_t (new_AGEMA_signal_14766), .Z1_f (new_AGEMA_signal_14767) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n129), .A0_f (new_AGEMA_signal_15446), .A1_t (new_AGEMA_signal_15447), .A1_f (new_AGEMA_signal_15448), .B0_t (MixColumnsInput[8]), .B0_f (new_AGEMA_signal_13295), .B1_t (new_AGEMA_signal_13296), .B1_f (new_AGEMA_signal_13297), .Z0_t (MixColumnsOutput[0]), .Z0_f (new_AGEMA_signal_16193), .Z1_t (new_AGEMA_signal_16194), .Z1_f (new_AGEMA_signal_16195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n187), .A0_f (new_AGEMA_signal_14771), .A1_t (new_AGEMA_signal_14772), .A1_f (new_AGEMA_signal_14773), .B0_t (MixColumnsIns_MixOneColumnInst_3_n151), .B0_f (new_AGEMA_signal_14768), .B1_t (new_AGEMA_signal_14769), .B1_f (new_AGEMA_signal_14770), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n129), .Z0_f (new_AGEMA_signal_15446), .Z1_t (new_AGEMA_signal_15447), .Z1_f (new_AGEMA_signal_15448) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U2 ( .A0_t (MixColumnsInput[16]), .A0_f (new_AGEMA_signal_13460), .A1_t (new_AGEMA_signal_13461), .A1_f (new_AGEMA_signal_13462), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B0_f (new_AGEMA_signal_13703), .B1_t (new_AGEMA_signal_13704), .B1_f (new_AGEMA_signal_13705), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n151), .Z0_f (new_AGEMA_signal_14768), .Z1_t (new_AGEMA_signal_14769), .Z1_f (new_AGEMA_signal_14770) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U1 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13724), .A1_t (new_AGEMA_signal_13725), .A1_f (new_AGEMA_signal_13726), .B0_t (MixColumnsInput[24]), .B0_f (new_AGEMA_signal_13097), .B1_t (new_AGEMA_signal_13098), .B1_f (new_AGEMA_signal_13099), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n187), .Z0_f (new_AGEMA_signal_14771), .Z1_t (new_AGEMA_signal_14772), .Z1_f (new_AGEMA_signal_14773) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13703), .A1_t (new_AGEMA_signal_13704), .A1_f (new_AGEMA_signal_13705), .B0_t (MixColumnsInput[27]), .B0_f (new_AGEMA_signal_13715), .B1_t (new_AGEMA_signal_13716), .B1_f (new_AGEMA_signal_13717), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]), .Z0_f (new_AGEMA_signal_14774), .Z1_t (new_AGEMA_signal_14775), .Z1_f (new_AGEMA_signal_14776) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13703), .A1_t (new_AGEMA_signal_13704), .A1_f (new_AGEMA_signal_13705), .B0_t (MixColumnsInput[26]), .B0_f (new_AGEMA_signal_13718), .B1_t (new_AGEMA_signal_13719), .B1_f (new_AGEMA_signal_13720), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]), .Z0_f (new_AGEMA_signal_14777), .Z1_t (new_AGEMA_signal_14778), .Z1_f (new_AGEMA_signal_14779) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .A0_f (new_AGEMA_signal_13703), .A1_t (new_AGEMA_signal_13704), .A1_f (new_AGEMA_signal_13705), .B0_t (MixColumnsInput[24]), .B0_f (new_AGEMA_signal_13097), .B1_t (new_AGEMA_signal_13098), .B1_f (new_AGEMA_signal_13099), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]), .Z0_f (new_AGEMA_signal_14780), .Z1_t (new_AGEMA_signal_14781), .Z1_f (new_AGEMA_signal_14782) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13934), .A1_t (new_AGEMA_signal_13935), .A1_f (new_AGEMA_signal_13936), .B0_t (MixColumnsInput[19]), .B0_f (new_AGEMA_signal_13946), .B1_t (new_AGEMA_signal_13947), .B1_f (new_AGEMA_signal_13948), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]), .Z0_f (new_AGEMA_signal_14783), .Z1_t (new_AGEMA_signal_14784), .Z1_f (new_AGEMA_signal_14785) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13934), .A1_t (new_AGEMA_signal_13935), .A1_f (new_AGEMA_signal_13936), .B0_t (MixColumnsInput[18]), .B0_f (new_AGEMA_signal_13949), .B1_t (new_AGEMA_signal_13950), .B1_f (new_AGEMA_signal_13951), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]), .Z0_f (new_AGEMA_signal_14786), .Z1_t (new_AGEMA_signal_14787), .Z1_f (new_AGEMA_signal_14788) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .A0_f (new_AGEMA_signal_13934), .A1_t (new_AGEMA_signal_13935), .A1_f (new_AGEMA_signal_13936), .B0_t (MixColumnsInput[16]), .B0_f (new_AGEMA_signal_13460), .B1_t (new_AGEMA_signal_13461), .B1_f (new_AGEMA_signal_13462), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]), .Z0_f (new_AGEMA_signal_14789), .Z1_t (new_AGEMA_signal_14790), .Z1_f (new_AGEMA_signal_14791) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13829), .A1_t (new_AGEMA_signal_13830), .A1_f (new_AGEMA_signal_13831), .B0_t (MixColumnsInput[11]), .B0_f (new_AGEMA_signal_13841), .B1_t (new_AGEMA_signal_13842), .B1_f (new_AGEMA_signal_13843), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]), .Z0_f (new_AGEMA_signal_14792), .Z1_t (new_AGEMA_signal_14793), .Z1_f (new_AGEMA_signal_14794) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13829), .A1_t (new_AGEMA_signal_13830), .A1_f (new_AGEMA_signal_13831), .B0_t (MixColumnsInput[10]), .B0_f (new_AGEMA_signal_13844), .B1_t (new_AGEMA_signal_13845), .B1_f (new_AGEMA_signal_13846), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]), .Z0_f (new_AGEMA_signal_14795), .Z1_t (new_AGEMA_signal_14796), .Z1_f (new_AGEMA_signal_14797) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .A0_f (new_AGEMA_signal_13829), .A1_t (new_AGEMA_signal_13830), .A1_f (new_AGEMA_signal_13831), .B0_t (MixColumnsInput[8]), .B0_f (new_AGEMA_signal_13295), .B1_t (new_AGEMA_signal_13296), .B1_f (new_AGEMA_signal_13297), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]), .Z0_f (new_AGEMA_signal_14798), .Z1_t (new_AGEMA_signal_14799), .Z1_f (new_AGEMA_signal_14800) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13724), .A1_t (new_AGEMA_signal_13725), .A1_f (new_AGEMA_signal_13726), .B0_t (MixColumnsInput[3]), .B0_f (new_AGEMA_signal_13736), .B1_t (new_AGEMA_signal_13737), .B1_f (new_AGEMA_signal_13738), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]), .Z0_f (new_AGEMA_signal_14801), .Z1_t (new_AGEMA_signal_14802), .Z1_f (new_AGEMA_signal_14803) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13724), .A1_t (new_AGEMA_signal_13725), .A1_f (new_AGEMA_signal_13726), .B0_t (MixColumnsInput[2]), .B0_f (new_AGEMA_signal_13739), .B1_t (new_AGEMA_signal_13740), .B1_f (new_AGEMA_signal_13741), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]), .Z0_f (new_AGEMA_signal_14804), .Z1_t (new_AGEMA_signal_14805), .Z1_f (new_AGEMA_signal_14806) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .A0_f (new_AGEMA_signal_13724), .A1_t (new_AGEMA_signal_13725), .A1_f (new_AGEMA_signal_13726), .B0_t (MixColumnsInput[0]), .B0_f (new_AGEMA_signal_13130), .B1_t (new_AGEMA_signal_13131), .B1_f (new_AGEMA_signal_13132), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]), .Z0_f (new_AGEMA_signal_14807), .Z1_t (new_AGEMA_signal_14808), .Z1_f (new_AGEMA_signal_14809) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_0_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[0]), .A0_f (new_AGEMA_signal_15809), .A1_t (new_AGEMA_signal_15810), .A1_f (new_AGEMA_signal_15811), .B0_t (key_s0_t[0]), .B0_f (key_s0_f[0]), .B1_t (key_s1_t[0]), .B1_f (key_s1_f[0]), .Z0_t (KeyReg_Inst_ff_SDE_0_MUX_inst_X), .Z0_f (new_AGEMA_signal_16199), .Z1_t (new_AGEMA_signal_16200), .Z1_f (new_AGEMA_signal_16201) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_0_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_0_MUX_inst_X), .B0_f (new_AGEMA_signal_16199), .B1_t (new_AGEMA_signal_16200), .B1_f (new_AGEMA_signal_16201), .Z0_t (KeyReg_Inst_ff_SDE_0_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16955), .Z1_t (new_AGEMA_signal_16956), .Z1_f (new_AGEMA_signal_16957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_0_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_0_MUX_inst_Y), .A0_f (new_AGEMA_signal_16955), .A1_t (new_AGEMA_signal_16956), .A1_f (new_AGEMA_signal_16957), .B0_t (KeyExpansionOutput[0]), .B0_f (new_AGEMA_signal_15809), .B1_t (new_AGEMA_signal_15810), .B1_f (new_AGEMA_signal_15811), .Z0_t (RoundKey[0]), .Z0_f (new_AGEMA_signal_5063), .Z1_t (new_AGEMA_signal_5064), .Z1_f (new_AGEMA_signal_5065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_1_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[1]), .A0_f (new_AGEMA_signal_16541), .A1_t (new_AGEMA_signal_16542), .A1_f (new_AGEMA_signal_16543), .B0_t (key_s0_t[1]), .B0_f (key_s0_f[1]), .B1_t (key_s1_t[1]), .B1_f (key_s1_f[1]), .Z0_t (KeyReg_Inst_ff_SDE_1_MUX_inst_X), .Z0_f (new_AGEMA_signal_16961), .Z1_t (new_AGEMA_signal_16962), .Z1_f (new_AGEMA_signal_16963) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_1_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_1_MUX_inst_X), .B0_f (new_AGEMA_signal_16961), .B1_t (new_AGEMA_signal_16962), .B1_f (new_AGEMA_signal_16963), .Z0_t (KeyReg_Inst_ff_SDE_1_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17630), .Z1_t (new_AGEMA_signal_17631), .Z1_f (new_AGEMA_signal_17632) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_1_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_1_MUX_inst_Y), .A0_f (new_AGEMA_signal_17630), .A1_t (new_AGEMA_signal_17631), .A1_f (new_AGEMA_signal_17632), .B0_t (KeyExpansionOutput[1]), .B0_f (new_AGEMA_signal_16541), .B1_t (new_AGEMA_signal_16542), .B1_f (new_AGEMA_signal_16543), .Z0_t (RoundKey[1]), .Z0_f (new_AGEMA_signal_5414), .Z1_t (new_AGEMA_signal_5415), .Z1_f (new_AGEMA_signal_5416) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_2_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[2]), .A0_f (new_AGEMA_signal_16508), .A1_t (new_AGEMA_signal_16509), .A1_f (new_AGEMA_signal_16510), .B0_t (key_s0_t[2]), .B0_f (key_s0_f[2]), .B1_t (key_s1_t[2]), .B1_f (key_s1_f[2]), .Z0_t (KeyReg_Inst_ff_SDE_2_MUX_inst_X), .Z0_f (new_AGEMA_signal_16967), .Z1_t (new_AGEMA_signal_16968), .Z1_f (new_AGEMA_signal_16969) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_2_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_2_MUX_inst_X), .B0_f (new_AGEMA_signal_16967), .B1_t (new_AGEMA_signal_16968), .B1_f (new_AGEMA_signal_16969), .Z0_t (KeyReg_Inst_ff_SDE_2_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17633), .Z1_t (new_AGEMA_signal_17634), .Z1_f (new_AGEMA_signal_17635) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_2_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_2_MUX_inst_Y), .A0_f (new_AGEMA_signal_17633), .A1_t (new_AGEMA_signal_17634), .A1_f (new_AGEMA_signal_17635), .B0_t (KeyExpansionOutput[2]), .B0_f (new_AGEMA_signal_16508), .B1_t (new_AGEMA_signal_16509), .B1_f (new_AGEMA_signal_16510), .Z0_t (RoundKey[2]), .Z0_f (new_AGEMA_signal_5513), .Z1_t (new_AGEMA_signal_5514), .Z1_f (new_AGEMA_signal_5515) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_3_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[3]), .A0_f (new_AGEMA_signal_16499), .A1_t (new_AGEMA_signal_16500), .A1_f (new_AGEMA_signal_16501), .B0_t (key_s0_t[3]), .B0_f (key_s0_f[3]), .B1_t (key_s1_t[3]), .B1_f (key_s1_f[3]), .Z0_t (KeyReg_Inst_ff_SDE_3_MUX_inst_X), .Z0_f (new_AGEMA_signal_16973), .Z1_t (new_AGEMA_signal_16974), .Z1_f (new_AGEMA_signal_16975) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_3_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_3_MUX_inst_X), .B0_f (new_AGEMA_signal_16973), .B1_t (new_AGEMA_signal_16974), .B1_f (new_AGEMA_signal_16975), .Z0_t (KeyReg_Inst_ff_SDE_3_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17636), .Z1_t (new_AGEMA_signal_17637), .Z1_f (new_AGEMA_signal_17638) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_3_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_3_MUX_inst_Y), .A0_f (new_AGEMA_signal_17636), .A1_t (new_AGEMA_signal_17637), .A1_f (new_AGEMA_signal_17638), .B0_t (KeyExpansionOutput[3]), .B0_f (new_AGEMA_signal_16499), .B1_t (new_AGEMA_signal_16500), .B1_f (new_AGEMA_signal_16501), .Z0_t (RoundKey[3]), .Z0_f (new_AGEMA_signal_5612), .Z1_t (new_AGEMA_signal_5613), .Z1_f (new_AGEMA_signal_5614) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_4_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[4]), .A0_f (new_AGEMA_signal_16496), .A1_t (new_AGEMA_signal_16497), .A1_f (new_AGEMA_signal_16498), .B0_t (key_s0_t[4]), .B0_f (key_s0_f[4]), .B1_t (key_s1_t[4]), .B1_f (key_s1_f[4]), .Z0_t (KeyReg_Inst_ff_SDE_4_MUX_inst_X), .Z0_f (new_AGEMA_signal_16979), .Z1_t (new_AGEMA_signal_16980), .Z1_f (new_AGEMA_signal_16981) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_4_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_4_MUX_inst_X), .B0_f (new_AGEMA_signal_16979), .B1_t (new_AGEMA_signal_16980), .B1_f (new_AGEMA_signal_16981), .Z0_t (KeyReg_Inst_ff_SDE_4_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17639), .Z1_t (new_AGEMA_signal_17640), .Z1_f (new_AGEMA_signal_17641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_4_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_4_MUX_inst_Y), .A0_f (new_AGEMA_signal_17639), .A1_t (new_AGEMA_signal_17640), .A1_f (new_AGEMA_signal_17641), .B0_t (KeyExpansionOutput[4]), .B0_f (new_AGEMA_signal_16496), .B1_t (new_AGEMA_signal_16497), .B1_f (new_AGEMA_signal_16498), .Z0_t (RoundKey[4]), .Z0_f (new_AGEMA_signal_5711), .Z1_t (new_AGEMA_signal_5712), .Z1_f (new_AGEMA_signal_5713) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_5_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[5]), .A0_f (new_AGEMA_signal_16493), .A1_t (new_AGEMA_signal_16494), .A1_f (new_AGEMA_signal_16495), .B0_t (key_s0_t[5]), .B0_f (key_s0_f[5]), .B1_t (key_s1_t[5]), .B1_f (key_s1_f[5]), .Z0_t (KeyReg_Inst_ff_SDE_5_MUX_inst_X), .Z0_f (new_AGEMA_signal_16985), .Z1_t (new_AGEMA_signal_16986), .Z1_f (new_AGEMA_signal_16987) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_5_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_5_MUX_inst_X), .B0_f (new_AGEMA_signal_16985), .B1_t (new_AGEMA_signal_16986), .B1_f (new_AGEMA_signal_16987), .Z0_t (KeyReg_Inst_ff_SDE_5_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17642), .Z1_t (new_AGEMA_signal_17643), .Z1_f (new_AGEMA_signal_17644) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_5_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_5_MUX_inst_Y), .A0_f (new_AGEMA_signal_17642), .A1_t (new_AGEMA_signal_17643), .A1_f (new_AGEMA_signal_17644), .B0_t (KeyExpansionOutput[5]), .B0_f (new_AGEMA_signal_16493), .B1_t (new_AGEMA_signal_16494), .B1_f (new_AGEMA_signal_16495), .Z0_t (RoundKey[5]), .Z0_f (new_AGEMA_signal_5810), .Z1_t (new_AGEMA_signal_5811), .Z1_f (new_AGEMA_signal_5812) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_6_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[6]), .A0_f (new_AGEMA_signal_16490), .A1_t (new_AGEMA_signal_16491), .A1_f (new_AGEMA_signal_16492), .B0_t (key_s0_t[6]), .B0_f (key_s0_f[6]), .B1_t (key_s1_t[6]), .B1_f (key_s1_f[6]), .Z0_t (KeyReg_Inst_ff_SDE_6_MUX_inst_X), .Z0_f (new_AGEMA_signal_16991), .Z1_t (new_AGEMA_signal_16992), .Z1_f (new_AGEMA_signal_16993) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_6_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_6_MUX_inst_X), .B0_f (new_AGEMA_signal_16991), .B1_t (new_AGEMA_signal_16992), .B1_f (new_AGEMA_signal_16993), .Z0_t (KeyReg_Inst_ff_SDE_6_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17645), .Z1_t (new_AGEMA_signal_17646), .Z1_f (new_AGEMA_signal_17647) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_6_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_6_MUX_inst_Y), .A0_f (new_AGEMA_signal_17645), .A1_t (new_AGEMA_signal_17646), .A1_f (new_AGEMA_signal_17647), .B0_t (KeyExpansionOutput[6]), .B0_f (new_AGEMA_signal_16490), .B1_t (new_AGEMA_signal_16491), .B1_f (new_AGEMA_signal_16492), .Z0_t (RoundKey[6]), .Z0_f (new_AGEMA_signal_5909), .Z1_t (new_AGEMA_signal_5910), .Z1_f (new_AGEMA_signal_5911) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_7_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[7]), .A0_f (new_AGEMA_signal_16487), .A1_t (new_AGEMA_signal_16488), .A1_f (new_AGEMA_signal_16489), .B0_t (key_s0_t[7]), .B0_f (key_s0_f[7]), .B1_t (key_s1_t[7]), .B1_f (key_s1_f[7]), .Z0_t (KeyReg_Inst_ff_SDE_7_MUX_inst_X), .Z0_f (new_AGEMA_signal_16997), .Z1_t (new_AGEMA_signal_16998), .Z1_f (new_AGEMA_signal_16999) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_7_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_7_MUX_inst_X), .B0_f (new_AGEMA_signal_16997), .B1_t (new_AGEMA_signal_16998), .B1_f (new_AGEMA_signal_16999), .Z0_t (KeyReg_Inst_ff_SDE_7_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17648), .Z1_t (new_AGEMA_signal_17649), .Z1_f (new_AGEMA_signal_17650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_7_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_7_MUX_inst_Y), .A0_f (new_AGEMA_signal_17648), .A1_t (new_AGEMA_signal_17649), .A1_f (new_AGEMA_signal_17650), .B0_t (KeyExpansionOutput[7]), .B0_f (new_AGEMA_signal_16487), .B1_t (new_AGEMA_signal_16488), .B1_f (new_AGEMA_signal_16489), .Z0_t (RoundKey[7]), .Z0_f (new_AGEMA_signal_6008), .Z1_t (new_AGEMA_signal_6009), .Z1_f (new_AGEMA_signal_6010) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_8_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[8]), .A0_f (new_AGEMA_signal_15716), .A1_t (new_AGEMA_signal_15717), .A1_f (new_AGEMA_signal_15718), .B0_t (key_s0_t[8]), .B0_f (key_s0_f[8]), .B1_t (key_s1_t[8]), .B1_f (key_s1_f[8]), .Z0_t (KeyReg_Inst_ff_SDE_8_MUX_inst_X), .Z0_f (new_AGEMA_signal_16205), .Z1_t (new_AGEMA_signal_16206), .Z1_f (new_AGEMA_signal_16207) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_8_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_8_MUX_inst_X), .B0_f (new_AGEMA_signal_16205), .B1_t (new_AGEMA_signal_16206), .B1_f (new_AGEMA_signal_16207), .Z0_t (KeyReg_Inst_ff_SDE_8_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17000), .Z1_t (new_AGEMA_signal_17001), .Z1_f (new_AGEMA_signal_17002) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_8_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_8_MUX_inst_Y), .A0_f (new_AGEMA_signal_17000), .A1_t (new_AGEMA_signal_17001), .A1_f (new_AGEMA_signal_17002), .B0_t (KeyExpansionOutput[8]), .B0_f (new_AGEMA_signal_15716), .B1_t (new_AGEMA_signal_15717), .B1_f (new_AGEMA_signal_15718), .Z0_t (RoundKey[8]), .Z0_f (new_AGEMA_signal_6107), .Z1_t (new_AGEMA_signal_6108), .Z1_f (new_AGEMA_signal_6109) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_9_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[9]), .A0_f (new_AGEMA_signal_16484), .A1_t (new_AGEMA_signal_16485), .A1_f (new_AGEMA_signal_16486), .B0_t (key_s0_t[9]), .B0_f (key_s0_f[9]), .B1_t (key_s1_t[9]), .B1_f (key_s1_f[9]), .Z0_t (KeyReg_Inst_ff_SDE_9_MUX_inst_X), .Z0_f (new_AGEMA_signal_17006), .Z1_t (new_AGEMA_signal_17007), .Z1_f (new_AGEMA_signal_17008) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_9_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_9_MUX_inst_X), .B0_f (new_AGEMA_signal_17006), .B1_t (new_AGEMA_signal_17007), .B1_f (new_AGEMA_signal_17008), .Z0_t (KeyReg_Inst_ff_SDE_9_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17651), .Z1_t (new_AGEMA_signal_17652), .Z1_f (new_AGEMA_signal_17653) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_9_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_9_MUX_inst_Y), .A0_f (new_AGEMA_signal_17651), .A1_t (new_AGEMA_signal_17652), .A1_f (new_AGEMA_signal_17653), .B0_t (KeyExpansionOutput[9]), .B0_f (new_AGEMA_signal_16484), .B1_t (new_AGEMA_signal_16485), .B1_f (new_AGEMA_signal_16486), .Z0_t (RoundKey[9]), .Z0_f (new_AGEMA_signal_6206), .Z1_t (new_AGEMA_signal_6207), .Z1_f (new_AGEMA_signal_6208) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_10_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[10]), .A0_f (new_AGEMA_signal_16568), .A1_t (new_AGEMA_signal_16569), .A1_f (new_AGEMA_signal_16570), .B0_t (key_s0_t[10]), .B0_f (key_s0_f[10]), .B1_t (key_s1_t[10]), .B1_f (key_s1_f[10]), .Z0_t (KeyReg_Inst_ff_SDE_10_MUX_inst_X), .Z0_f (new_AGEMA_signal_17012), .Z1_t (new_AGEMA_signal_17013), .Z1_f (new_AGEMA_signal_17014) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_10_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_10_MUX_inst_X), .B0_f (new_AGEMA_signal_17012), .B1_t (new_AGEMA_signal_17013), .B1_f (new_AGEMA_signal_17014), .Z0_t (KeyReg_Inst_ff_SDE_10_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17654), .Z1_t (new_AGEMA_signal_17655), .Z1_f (new_AGEMA_signal_17656) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_10_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_10_MUX_inst_Y), .A0_f (new_AGEMA_signal_17654), .A1_t (new_AGEMA_signal_17655), .A1_f (new_AGEMA_signal_17656), .B0_t (KeyExpansionOutput[10]), .B0_f (new_AGEMA_signal_16568), .B1_t (new_AGEMA_signal_16569), .B1_f (new_AGEMA_signal_16570), .Z0_t (RoundKey[10]), .Z0_f (new_AGEMA_signal_5162), .Z1_t (new_AGEMA_signal_5163), .Z1_f (new_AGEMA_signal_5164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_11_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[11]), .A0_f (new_AGEMA_signal_16565), .A1_t (new_AGEMA_signal_16566), .A1_f (new_AGEMA_signal_16567), .B0_t (key_s0_t[11]), .B0_f (key_s0_f[11]), .B1_t (key_s1_t[11]), .B1_f (key_s1_f[11]), .Z0_t (KeyReg_Inst_ff_SDE_11_MUX_inst_X), .Z0_f (new_AGEMA_signal_17018), .Z1_t (new_AGEMA_signal_17019), .Z1_f (new_AGEMA_signal_17020) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_11_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_11_MUX_inst_X), .B0_f (new_AGEMA_signal_17018), .B1_t (new_AGEMA_signal_17019), .B1_f (new_AGEMA_signal_17020), .Z0_t (KeyReg_Inst_ff_SDE_11_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17657), .Z1_t (new_AGEMA_signal_17658), .Z1_f (new_AGEMA_signal_17659) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_11_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_11_MUX_inst_Y), .A0_f (new_AGEMA_signal_17657), .A1_t (new_AGEMA_signal_17658), .A1_f (new_AGEMA_signal_17659), .B0_t (KeyExpansionOutput[11]), .B0_f (new_AGEMA_signal_16565), .B1_t (new_AGEMA_signal_16566), .B1_f (new_AGEMA_signal_16567), .Z0_t (RoundKey[11]), .Z0_f (new_AGEMA_signal_5261), .Z1_t (new_AGEMA_signal_5262), .Z1_f (new_AGEMA_signal_5263) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_12_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[12]), .A0_f (new_AGEMA_signal_16562), .A1_t (new_AGEMA_signal_16563), .A1_f (new_AGEMA_signal_16564), .B0_t (key_s0_t[12]), .B0_f (key_s0_f[12]), .B1_t (key_s1_t[12]), .B1_f (key_s1_f[12]), .Z0_t (KeyReg_Inst_ff_SDE_12_MUX_inst_X), .Z0_f (new_AGEMA_signal_17024), .Z1_t (new_AGEMA_signal_17025), .Z1_f (new_AGEMA_signal_17026) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_12_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_12_MUX_inst_X), .B0_f (new_AGEMA_signal_17024), .B1_t (new_AGEMA_signal_17025), .B1_f (new_AGEMA_signal_17026), .Z0_t (KeyReg_Inst_ff_SDE_12_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17660), .Z1_t (new_AGEMA_signal_17661), .Z1_f (new_AGEMA_signal_17662) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_12_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_12_MUX_inst_Y), .A0_f (new_AGEMA_signal_17660), .A1_t (new_AGEMA_signal_17661), .A1_f (new_AGEMA_signal_17662), .B0_t (KeyExpansionOutput[12]), .B0_f (new_AGEMA_signal_16562), .B1_t (new_AGEMA_signal_16563), .B1_f (new_AGEMA_signal_16564), .Z0_t (RoundKey[12]), .Z0_f (new_AGEMA_signal_5342), .Z1_t (new_AGEMA_signal_5343), .Z1_f (new_AGEMA_signal_5344) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_13_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[13]), .A0_f (new_AGEMA_signal_16559), .A1_t (new_AGEMA_signal_16560), .A1_f (new_AGEMA_signal_16561), .B0_t (key_s0_t[13]), .B0_f (key_s0_f[13]), .B1_t (key_s1_t[13]), .B1_f (key_s1_f[13]), .Z0_t (KeyReg_Inst_ff_SDE_13_MUX_inst_X), .Z0_f (new_AGEMA_signal_17030), .Z1_t (new_AGEMA_signal_17031), .Z1_f (new_AGEMA_signal_17032) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_13_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_13_MUX_inst_X), .B0_f (new_AGEMA_signal_17030), .B1_t (new_AGEMA_signal_17031), .B1_f (new_AGEMA_signal_17032), .Z0_t (KeyReg_Inst_ff_SDE_13_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17663), .Z1_t (new_AGEMA_signal_17664), .Z1_f (new_AGEMA_signal_17665) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_13_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_13_MUX_inst_Y), .A0_f (new_AGEMA_signal_17663), .A1_t (new_AGEMA_signal_17664), .A1_f (new_AGEMA_signal_17665), .B0_t (KeyExpansionOutput[13]), .B0_f (new_AGEMA_signal_16559), .B1_t (new_AGEMA_signal_16560), .B1_f (new_AGEMA_signal_16561), .Z0_t (RoundKey[13]), .Z0_f (new_AGEMA_signal_5351), .Z1_t (new_AGEMA_signal_5352), .Z1_f (new_AGEMA_signal_5353) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_14_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[14]), .A0_f (new_AGEMA_signal_16556), .A1_t (new_AGEMA_signal_16557), .A1_f (new_AGEMA_signal_16558), .B0_t (key_s0_t[14]), .B0_f (key_s0_f[14]), .B1_t (key_s1_t[14]), .B1_f (key_s1_f[14]), .Z0_t (KeyReg_Inst_ff_SDE_14_MUX_inst_X), .Z0_f (new_AGEMA_signal_17036), .Z1_t (new_AGEMA_signal_17037), .Z1_f (new_AGEMA_signal_17038) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_14_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_14_MUX_inst_X), .B0_f (new_AGEMA_signal_17036), .B1_t (new_AGEMA_signal_17037), .B1_f (new_AGEMA_signal_17038), .Z0_t (KeyReg_Inst_ff_SDE_14_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17666), .Z1_t (new_AGEMA_signal_17667), .Z1_f (new_AGEMA_signal_17668) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_14_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_14_MUX_inst_Y), .A0_f (new_AGEMA_signal_17666), .A1_t (new_AGEMA_signal_17667), .A1_f (new_AGEMA_signal_17668), .B0_t (KeyExpansionOutput[14]), .B0_f (new_AGEMA_signal_16556), .B1_t (new_AGEMA_signal_16557), .B1_f (new_AGEMA_signal_16558), .Z0_t (RoundKey[14]), .Z0_f (new_AGEMA_signal_5360), .Z1_t (new_AGEMA_signal_5361), .Z1_f (new_AGEMA_signal_5362) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_15_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[15]), .A0_f (new_AGEMA_signal_16553), .A1_t (new_AGEMA_signal_16554), .A1_f (new_AGEMA_signal_16555), .B0_t (key_s0_t[15]), .B0_f (key_s0_f[15]), .B1_t (key_s1_t[15]), .B1_f (key_s1_f[15]), .Z0_t (KeyReg_Inst_ff_SDE_15_MUX_inst_X), .Z0_f (new_AGEMA_signal_17042), .Z1_t (new_AGEMA_signal_17043), .Z1_f (new_AGEMA_signal_17044) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_15_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_15_MUX_inst_X), .B0_f (new_AGEMA_signal_17042), .B1_t (new_AGEMA_signal_17043), .B1_f (new_AGEMA_signal_17044), .Z0_t (KeyReg_Inst_ff_SDE_15_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17669), .Z1_t (new_AGEMA_signal_17670), .Z1_f (new_AGEMA_signal_17671) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_15_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_15_MUX_inst_Y), .A0_f (new_AGEMA_signal_17669), .A1_t (new_AGEMA_signal_17670), .A1_f (new_AGEMA_signal_17671), .B0_t (KeyExpansionOutput[15]), .B0_f (new_AGEMA_signal_16553), .B1_t (new_AGEMA_signal_16554), .B1_f (new_AGEMA_signal_16555), .Z0_t (RoundKey[15]), .Z0_f (new_AGEMA_signal_5369), .Z1_t (new_AGEMA_signal_5370), .Z1_f (new_AGEMA_signal_5371) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_16_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[16]), .A0_f (new_AGEMA_signal_15788), .A1_t (new_AGEMA_signal_15789), .A1_f (new_AGEMA_signal_15790), .B0_t (key_s0_t[16]), .B0_f (key_s0_f[16]), .B1_t (key_s1_t[16]), .B1_f (key_s1_f[16]), .Z0_t (KeyReg_Inst_ff_SDE_16_MUX_inst_X), .Z0_f (new_AGEMA_signal_16211), .Z1_t (new_AGEMA_signal_16212), .Z1_f (new_AGEMA_signal_16213) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_16_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_16_MUX_inst_X), .B0_f (new_AGEMA_signal_16211), .B1_t (new_AGEMA_signal_16212), .B1_f (new_AGEMA_signal_16213), .Z0_t (KeyReg_Inst_ff_SDE_16_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17045), .Z1_t (new_AGEMA_signal_17046), .Z1_f (new_AGEMA_signal_17047) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_16_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_16_MUX_inst_Y), .A0_f (new_AGEMA_signal_17045), .A1_t (new_AGEMA_signal_17046), .A1_f (new_AGEMA_signal_17047), .B0_t (KeyExpansionOutput[16]), .B0_f (new_AGEMA_signal_15788), .B1_t (new_AGEMA_signal_15789), .B1_f (new_AGEMA_signal_15790), .Z0_t (RoundKey[16]), .Z0_f (new_AGEMA_signal_5378), .Z1_t (new_AGEMA_signal_5379), .Z1_f (new_AGEMA_signal_5380) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_17_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[17]), .A0_f (new_AGEMA_signal_16550), .A1_t (new_AGEMA_signal_16551), .A1_f (new_AGEMA_signal_16552), .B0_t (key_s0_t[17]), .B0_f (key_s0_f[17]), .B1_t (key_s1_t[17]), .B1_f (key_s1_f[17]), .Z0_t (KeyReg_Inst_ff_SDE_17_MUX_inst_X), .Z0_f (new_AGEMA_signal_17051), .Z1_t (new_AGEMA_signal_17052), .Z1_f (new_AGEMA_signal_17053) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_17_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_17_MUX_inst_X), .B0_f (new_AGEMA_signal_17051), .B1_t (new_AGEMA_signal_17052), .B1_f (new_AGEMA_signal_17053), .Z0_t (KeyReg_Inst_ff_SDE_17_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17672), .Z1_t (new_AGEMA_signal_17673), .Z1_f (new_AGEMA_signal_17674) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_17_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_17_MUX_inst_Y), .A0_f (new_AGEMA_signal_17672), .A1_t (new_AGEMA_signal_17673), .A1_f (new_AGEMA_signal_17674), .B0_t (KeyExpansionOutput[17]), .B0_f (new_AGEMA_signal_16550), .B1_t (new_AGEMA_signal_16551), .B1_f (new_AGEMA_signal_16552), .Z0_t (RoundKey[17]), .Z0_f (new_AGEMA_signal_5387), .Z1_t (new_AGEMA_signal_5388), .Z1_f (new_AGEMA_signal_5389) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_18_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[18]), .A0_f (new_AGEMA_signal_16547), .A1_t (new_AGEMA_signal_16548), .A1_f (new_AGEMA_signal_16549), .B0_t (key_s0_t[18]), .B0_f (key_s0_f[18]), .B1_t (key_s1_t[18]), .B1_f (key_s1_f[18]), .Z0_t (KeyReg_Inst_ff_SDE_18_MUX_inst_X), .Z0_f (new_AGEMA_signal_17057), .Z1_t (new_AGEMA_signal_17058), .Z1_f (new_AGEMA_signal_17059) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_18_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_18_MUX_inst_X), .B0_f (new_AGEMA_signal_17057), .B1_t (new_AGEMA_signal_17058), .B1_f (new_AGEMA_signal_17059), .Z0_t (KeyReg_Inst_ff_SDE_18_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17675), .Z1_t (new_AGEMA_signal_17676), .Z1_f (new_AGEMA_signal_17677) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_18_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_18_MUX_inst_Y), .A0_f (new_AGEMA_signal_17675), .A1_t (new_AGEMA_signal_17676), .A1_f (new_AGEMA_signal_17677), .B0_t (KeyExpansionOutput[18]), .B0_f (new_AGEMA_signal_16547), .B1_t (new_AGEMA_signal_16548), .B1_f (new_AGEMA_signal_16549), .Z0_t (RoundKey[18]), .Z0_f (new_AGEMA_signal_5396), .Z1_t (new_AGEMA_signal_5397), .Z1_f (new_AGEMA_signal_5398) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_19_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[19]), .A0_f (new_AGEMA_signal_16544), .A1_t (new_AGEMA_signal_16545), .A1_f (new_AGEMA_signal_16546), .B0_t (key_s0_t[19]), .B0_f (key_s0_f[19]), .B1_t (key_s1_t[19]), .B1_f (key_s1_f[19]), .Z0_t (KeyReg_Inst_ff_SDE_19_MUX_inst_X), .Z0_f (new_AGEMA_signal_17063), .Z1_t (new_AGEMA_signal_17064), .Z1_f (new_AGEMA_signal_17065) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_19_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_19_MUX_inst_X), .B0_f (new_AGEMA_signal_17063), .B1_t (new_AGEMA_signal_17064), .B1_f (new_AGEMA_signal_17065), .Z0_t (KeyReg_Inst_ff_SDE_19_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17678), .Z1_t (new_AGEMA_signal_17679), .Z1_f (new_AGEMA_signal_17680) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_19_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_19_MUX_inst_Y), .A0_f (new_AGEMA_signal_17678), .A1_t (new_AGEMA_signal_17679), .A1_f (new_AGEMA_signal_17680), .B0_t (KeyExpansionOutput[19]), .B0_f (new_AGEMA_signal_16544), .B1_t (new_AGEMA_signal_16545), .B1_f (new_AGEMA_signal_16546), .Z0_t (RoundKey[19]), .Z0_f (new_AGEMA_signal_5405), .Z1_t (new_AGEMA_signal_5406), .Z1_f (new_AGEMA_signal_5407) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_20_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[20]), .A0_f (new_AGEMA_signal_16538), .A1_t (new_AGEMA_signal_16539), .A1_f (new_AGEMA_signal_16540), .B0_t (key_s0_t[20]), .B0_f (key_s0_f[20]), .B1_t (key_s1_t[20]), .B1_f (key_s1_f[20]), .Z0_t (KeyReg_Inst_ff_SDE_20_MUX_inst_X), .Z0_f (new_AGEMA_signal_17069), .Z1_t (new_AGEMA_signal_17070), .Z1_f (new_AGEMA_signal_17071) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_20_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_20_MUX_inst_X), .B0_f (new_AGEMA_signal_17069), .B1_t (new_AGEMA_signal_17070), .B1_f (new_AGEMA_signal_17071), .Z0_t (KeyReg_Inst_ff_SDE_20_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17681), .Z1_t (new_AGEMA_signal_17682), .Z1_f (new_AGEMA_signal_17683) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_20_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_20_MUX_inst_Y), .A0_f (new_AGEMA_signal_17681), .A1_t (new_AGEMA_signal_17682), .A1_f (new_AGEMA_signal_17683), .B0_t (KeyExpansionOutput[20]), .B0_f (new_AGEMA_signal_16538), .B1_t (new_AGEMA_signal_16539), .B1_f (new_AGEMA_signal_16540), .Z0_t (RoundKey[20]), .Z0_f (new_AGEMA_signal_5423), .Z1_t (new_AGEMA_signal_5424), .Z1_f (new_AGEMA_signal_5425) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_21_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[21]), .A0_f (new_AGEMA_signal_16535), .A1_t (new_AGEMA_signal_16536), .A1_f (new_AGEMA_signal_16537), .B0_t (key_s0_t[21]), .B0_f (key_s0_f[21]), .B1_t (key_s1_t[21]), .B1_f (key_s1_f[21]), .Z0_t (KeyReg_Inst_ff_SDE_21_MUX_inst_X), .Z0_f (new_AGEMA_signal_17075), .Z1_t (new_AGEMA_signal_17076), .Z1_f (new_AGEMA_signal_17077) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_21_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_21_MUX_inst_X), .B0_f (new_AGEMA_signal_17075), .B1_t (new_AGEMA_signal_17076), .B1_f (new_AGEMA_signal_17077), .Z0_t (KeyReg_Inst_ff_SDE_21_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17684), .Z1_t (new_AGEMA_signal_17685), .Z1_f (new_AGEMA_signal_17686) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_21_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_21_MUX_inst_Y), .A0_f (new_AGEMA_signal_17684), .A1_t (new_AGEMA_signal_17685), .A1_f (new_AGEMA_signal_17686), .B0_t (KeyExpansionOutput[21]), .B0_f (new_AGEMA_signal_16535), .B1_t (new_AGEMA_signal_16536), .B1_f (new_AGEMA_signal_16537), .Z0_t (RoundKey[21]), .Z0_f (new_AGEMA_signal_5432), .Z1_t (new_AGEMA_signal_5433), .Z1_f (new_AGEMA_signal_5434) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_22_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[22]), .A0_f (new_AGEMA_signal_16532), .A1_t (new_AGEMA_signal_16533), .A1_f (new_AGEMA_signal_16534), .B0_t (key_s0_t[22]), .B0_f (key_s0_f[22]), .B1_t (key_s1_t[22]), .B1_f (key_s1_f[22]), .Z0_t (KeyReg_Inst_ff_SDE_22_MUX_inst_X), .Z0_f (new_AGEMA_signal_17081), .Z1_t (new_AGEMA_signal_17082), .Z1_f (new_AGEMA_signal_17083) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_22_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_22_MUX_inst_X), .B0_f (new_AGEMA_signal_17081), .B1_t (new_AGEMA_signal_17082), .B1_f (new_AGEMA_signal_17083), .Z0_t (KeyReg_Inst_ff_SDE_22_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17687), .Z1_t (new_AGEMA_signal_17688), .Z1_f (new_AGEMA_signal_17689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_22_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_22_MUX_inst_Y), .A0_f (new_AGEMA_signal_17687), .A1_t (new_AGEMA_signal_17688), .A1_f (new_AGEMA_signal_17689), .B0_t (KeyExpansionOutput[22]), .B0_f (new_AGEMA_signal_16532), .B1_t (new_AGEMA_signal_16533), .B1_f (new_AGEMA_signal_16534), .Z0_t (RoundKey[22]), .Z0_f (new_AGEMA_signal_5441), .Z1_t (new_AGEMA_signal_5442), .Z1_f (new_AGEMA_signal_5443) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_23_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[23]), .A0_f (new_AGEMA_signal_16529), .A1_t (new_AGEMA_signal_16530), .A1_f (new_AGEMA_signal_16531), .B0_t (key_s0_t[23]), .B0_f (key_s0_f[23]), .B1_t (key_s1_t[23]), .B1_f (key_s1_f[23]), .Z0_t (KeyReg_Inst_ff_SDE_23_MUX_inst_X), .Z0_f (new_AGEMA_signal_17087), .Z1_t (new_AGEMA_signal_17088), .Z1_f (new_AGEMA_signal_17089) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_23_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_23_MUX_inst_X), .B0_f (new_AGEMA_signal_17087), .B1_t (new_AGEMA_signal_17088), .B1_f (new_AGEMA_signal_17089), .Z0_t (KeyReg_Inst_ff_SDE_23_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17690), .Z1_t (new_AGEMA_signal_17691), .Z1_f (new_AGEMA_signal_17692) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_23_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_23_MUX_inst_Y), .A0_f (new_AGEMA_signal_17690), .A1_t (new_AGEMA_signal_17691), .A1_f (new_AGEMA_signal_17692), .B0_t (KeyExpansionOutput[23]), .B0_f (new_AGEMA_signal_16529), .B1_t (new_AGEMA_signal_16530), .B1_f (new_AGEMA_signal_16531), .Z0_t (RoundKey[23]), .Z0_f (new_AGEMA_signal_5450), .Z1_t (new_AGEMA_signal_5451), .Z1_f (new_AGEMA_signal_5452) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_24_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[24]), .A0_f (new_AGEMA_signal_16526), .A1_t (new_AGEMA_signal_16527), .A1_f (new_AGEMA_signal_16528), .B0_t (key_s0_t[24]), .B0_f (key_s0_f[24]), .B1_t (key_s1_t[24]), .B1_f (key_s1_f[24]), .Z0_t (KeyReg_Inst_ff_SDE_24_MUX_inst_X), .Z0_f (new_AGEMA_signal_17093), .Z1_t (new_AGEMA_signal_17094), .Z1_f (new_AGEMA_signal_17095) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_24_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_24_MUX_inst_X), .B0_f (new_AGEMA_signal_17093), .B1_t (new_AGEMA_signal_17094), .B1_f (new_AGEMA_signal_17095), .Z0_t (KeyReg_Inst_ff_SDE_24_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17693), .Z1_t (new_AGEMA_signal_17694), .Z1_f (new_AGEMA_signal_17695) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_24_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_24_MUX_inst_Y), .A0_f (new_AGEMA_signal_17693), .A1_t (new_AGEMA_signal_17694), .A1_f (new_AGEMA_signal_17695), .B0_t (KeyExpansionOutput[24]), .B0_f (new_AGEMA_signal_16526), .B1_t (new_AGEMA_signal_16527), .B1_f (new_AGEMA_signal_16528), .Z0_t (RoundKey[24]), .Z0_f (new_AGEMA_signal_5459), .Z1_t (new_AGEMA_signal_5460), .Z1_f (new_AGEMA_signal_5461) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_25_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[25]), .A0_f (new_AGEMA_signal_17243), .A1_t (new_AGEMA_signal_17244), .A1_f (new_AGEMA_signal_17245), .B0_t (key_s0_t[25]), .B0_f (key_s0_f[25]), .B1_t (key_s1_t[25]), .B1_f (key_s1_f[25]), .Z0_t (KeyReg_Inst_ff_SDE_25_MUX_inst_X), .Z0_f (new_AGEMA_signal_17699), .Z1_t (new_AGEMA_signal_17700), .Z1_f (new_AGEMA_signal_17701) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_25_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_25_MUX_inst_X), .B0_f (new_AGEMA_signal_17699), .B1_t (new_AGEMA_signal_17700), .B1_f (new_AGEMA_signal_17701), .Z0_t (KeyReg_Inst_ff_SDE_25_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18383), .Z1_t (new_AGEMA_signal_18384), .Z1_f (new_AGEMA_signal_18385) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_25_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_25_MUX_inst_Y), .A0_f (new_AGEMA_signal_18383), .A1_t (new_AGEMA_signal_18384), .A1_f (new_AGEMA_signal_18385), .B0_t (KeyExpansionOutput[25]), .B0_f (new_AGEMA_signal_17243), .B1_t (new_AGEMA_signal_17244), .B1_f (new_AGEMA_signal_17245), .Z0_t (RoundKey[25]), .Z0_f (new_AGEMA_signal_5468), .Z1_t (new_AGEMA_signal_5469), .Z1_f (new_AGEMA_signal_5470) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_26_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[26]), .A0_f (new_AGEMA_signal_17240), .A1_t (new_AGEMA_signal_17241), .A1_f (new_AGEMA_signal_17242), .B0_t (key_s0_t[26]), .B0_f (key_s0_f[26]), .B1_t (key_s1_t[26]), .B1_f (key_s1_f[26]), .Z0_t (KeyReg_Inst_ff_SDE_26_MUX_inst_X), .Z0_f (new_AGEMA_signal_17705), .Z1_t (new_AGEMA_signal_17706), .Z1_f (new_AGEMA_signal_17707) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_26_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_26_MUX_inst_X), .B0_f (new_AGEMA_signal_17705), .B1_t (new_AGEMA_signal_17706), .B1_f (new_AGEMA_signal_17707), .Z0_t (KeyReg_Inst_ff_SDE_26_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18386), .Z1_t (new_AGEMA_signal_18387), .Z1_f (new_AGEMA_signal_18388) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_26_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_26_MUX_inst_Y), .A0_f (new_AGEMA_signal_18386), .A1_t (new_AGEMA_signal_18387), .A1_f (new_AGEMA_signal_18388), .B0_t (KeyExpansionOutput[26]), .B0_f (new_AGEMA_signal_17240), .B1_t (new_AGEMA_signal_17241), .B1_f (new_AGEMA_signal_17242), .Z0_t (RoundKey[26]), .Z0_f (new_AGEMA_signal_5477), .Z1_t (new_AGEMA_signal_5478), .Z1_f (new_AGEMA_signal_5479) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_27_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[27]), .A0_f (new_AGEMA_signal_17237), .A1_t (new_AGEMA_signal_17238), .A1_f (new_AGEMA_signal_17239), .B0_t (key_s0_t[27]), .B0_f (key_s0_f[27]), .B1_t (key_s1_t[27]), .B1_f (key_s1_f[27]), .Z0_t (KeyReg_Inst_ff_SDE_27_MUX_inst_X), .Z0_f (new_AGEMA_signal_17711), .Z1_t (new_AGEMA_signal_17712), .Z1_f (new_AGEMA_signal_17713) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_27_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_27_MUX_inst_X), .B0_f (new_AGEMA_signal_17711), .B1_t (new_AGEMA_signal_17712), .B1_f (new_AGEMA_signal_17713), .Z0_t (KeyReg_Inst_ff_SDE_27_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18389), .Z1_t (new_AGEMA_signal_18390), .Z1_f (new_AGEMA_signal_18391) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_27_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_27_MUX_inst_Y), .A0_f (new_AGEMA_signal_18389), .A1_t (new_AGEMA_signal_18390), .A1_f (new_AGEMA_signal_18391), .B0_t (KeyExpansionOutput[27]), .B0_f (new_AGEMA_signal_17237), .B1_t (new_AGEMA_signal_17238), .B1_f (new_AGEMA_signal_17239), .Z0_t (RoundKey[27]), .Z0_f (new_AGEMA_signal_5486), .Z1_t (new_AGEMA_signal_5487), .Z1_f (new_AGEMA_signal_5488) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_28_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[28]), .A0_f (new_AGEMA_signal_17234), .A1_t (new_AGEMA_signal_17235), .A1_f (new_AGEMA_signal_17236), .B0_t (key_s0_t[28]), .B0_f (key_s0_f[28]), .B1_t (key_s1_t[28]), .B1_f (key_s1_f[28]), .Z0_t (KeyReg_Inst_ff_SDE_28_MUX_inst_X), .Z0_f (new_AGEMA_signal_17717), .Z1_t (new_AGEMA_signal_17718), .Z1_f (new_AGEMA_signal_17719) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_28_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_28_MUX_inst_X), .B0_f (new_AGEMA_signal_17717), .B1_t (new_AGEMA_signal_17718), .B1_f (new_AGEMA_signal_17719), .Z0_t (KeyReg_Inst_ff_SDE_28_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18392), .Z1_t (new_AGEMA_signal_18393), .Z1_f (new_AGEMA_signal_18394) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_28_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_28_MUX_inst_Y), .A0_f (new_AGEMA_signal_18392), .A1_t (new_AGEMA_signal_18393), .A1_f (new_AGEMA_signal_18394), .B0_t (KeyExpansionOutput[28]), .B0_f (new_AGEMA_signal_17234), .B1_t (new_AGEMA_signal_17235), .B1_f (new_AGEMA_signal_17236), .Z0_t (RoundKey[28]), .Z0_f (new_AGEMA_signal_5495), .Z1_t (new_AGEMA_signal_5496), .Z1_f (new_AGEMA_signal_5497) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_29_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[29]), .A0_f (new_AGEMA_signal_17231), .A1_t (new_AGEMA_signal_17232), .A1_f (new_AGEMA_signal_17233), .B0_t (key_s0_t[29]), .B0_f (key_s0_f[29]), .B1_t (key_s1_t[29]), .B1_f (key_s1_f[29]), .Z0_t (KeyReg_Inst_ff_SDE_29_MUX_inst_X), .Z0_f (new_AGEMA_signal_17723), .Z1_t (new_AGEMA_signal_17724), .Z1_f (new_AGEMA_signal_17725) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_29_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_29_MUX_inst_X), .B0_f (new_AGEMA_signal_17723), .B1_t (new_AGEMA_signal_17724), .B1_f (new_AGEMA_signal_17725), .Z0_t (KeyReg_Inst_ff_SDE_29_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18395), .Z1_t (new_AGEMA_signal_18396), .Z1_f (new_AGEMA_signal_18397) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_29_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_29_MUX_inst_Y), .A0_f (new_AGEMA_signal_18395), .A1_t (new_AGEMA_signal_18396), .A1_f (new_AGEMA_signal_18397), .B0_t (KeyExpansionOutput[29]), .B0_f (new_AGEMA_signal_17231), .B1_t (new_AGEMA_signal_17232), .B1_f (new_AGEMA_signal_17233), .Z0_t (RoundKey[29]), .Z0_f (new_AGEMA_signal_5504), .Z1_t (new_AGEMA_signal_5505), .Z1_f (new_AGEMA_signal_5506) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_30_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[30]), .A0_f (new_AGEMA_signal_17228), .A1_t (new_AGEMA_signal_17229), .A1_f (new_AGEMA_signal_17230), .B0_t (key_s0_t[30]), .B0_f (key_s0_f[30]), .B1_t (key_s1_t[30]), .B1_f (key_s1_f[30]), .Z0_t (KeyReg_Inst_ff_SDE_30_MUX_inst_X), .Z0_f (new_AGEMA_signal_17729), .Z1_t (new_AGEMA_signal_17730), .Z1_f (new_AGEMA_signal_17731) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_30_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_30_MUX_inst_X), .B0_f (new_AGEMA_signal_17729), .B1_t (new_AGEMA_signal_17730), .B1_f (new_AGEMA_signal_17731), .Z0_t (KeyReg_Inst_ff_SDE_30_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18398), .Z1_t (new_AGEMA_signal_18399), .Z1_f (new_AGEMA_signal_18400) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_30_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_30_MUX_inst_Y), .A0_f (new_AGEMA_signal_18398), .A1_t (new_AGEMA_signal_18399), .A1_f (new_AGEMA_signal_18400), .B0_t (KeyExpansionOutput[30]), .B0_f (new_AGEMA_signal_17228), .B1_t (new_AGEMA_signal_17229), .B1_f (new_AGEMA_signal_17230), .Z0_t (RoundKey[30]), .Z0_f (new_AGEMA_signal_5522), .Z1_t (new_AGEMA_signal_5523), .Z1_f (new_AGEMA_signal_5524) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_31_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[31]), .A0_f (new_AGEMA_signal_17225), .A1_t (new_AGEMA_signal_17226), .A1_f (new_AGEMA_signal_17227), .B0_t (key_s0_t[31]), .B0_f (key_s0_f[31]), .B1_t (key_s1_t[31]), .B1_f (key_s1_f[31]), .Z0_t (KeyReg_Inst_ff_SDE_31_MUX_inst_X), .Z0_f (new_AGEMA_signal_17735), .Z1_t (new_AGEMA_signal_17736), .Z1_f (new_AGEMA_signal_17737) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_31_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_31_MUX_inst_X), .B0_f (new_AGEMA_signal_17735), .B1_t (new_AGEMA_signal_17736), .B1_f (new_AGEMA_signal_17737), .Z0_t (KeyReg_Inst_ff_SDE_31_MUX_inst_Y), .Z0_f (new_AGEMA_signal_18401), .Z1_t (new_AGEMA_signal_18402), .Z1_f (new_AGEMA_signal_18403) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_31_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_31_MUX_inst_Y), .A0_f (new_AGEMA_signal_18401), .A1_t (new_AGEMA_signal_18402), .A1_f (new_AGEMA_signal_18403), .B0_t (KeyExpansionOutput[31]), .B0_f (new_AGEMA_signal_17225), .B1_t (new_AGEMA_signal_17226), .B1_f (new_AGEMA_signal_17227), .Z0_t (RoundKey[31]), .Z0_f (new_AGEMA_signal_5531), .Z1_t (new_AGEMA_signal_5532), .Z1_f (new_AGEMA_signal_5533) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_32_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[32]), .A0_f (new_AGEMA_signal_15062), .A1_t (new_AGEMA_signal_15063), .A1_f (new_AGEMA_signal_15064), .B0_t (key_s0_t[32]), .B0_f (key_s0_f[32]), .B1_t (key_s1_t[32]), .B1_f (key_s1_f[32]), .Z0_t (KeyReg_Inst_ff_SDE_32_MUX_inst_X), .Z0_f (new_AGEMA_signal_15452), .Z1_t (new_AGEMA_signal_15453), .Z1_f (new_AGEMA_signal_15454) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_32_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_32_MUX_inst_X), .B0_f (new_AGEMA_signal_15452), .B1_t (new_AGEMA_signal_15453), .B1_f (new_AGEMA_signal_15454), .Z0_t (KeyReg_Inst_ff_SDE_32_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16214), .Z1_t (new_AGEMA_signal_16215), .Z1_f (new_AGEMA_signal_16216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_32_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_32_MUX_inst_Y), .A0_f (new_AGEMA_signal_16214), .A1_t (new_AGEMA_signal_16215), .A1_f (new_AGEMA_signal_16216), .B0_t (KeyExpansionOutput[32]), .B0_f (new_AGEMA_signal_15062), .B1_t (new_AGEMA_signal_15063), .B1_f (new_AGEMA_signal_15064), .Z0_t (RoundKey[32]), .Z0_f (new_AGEMA_signal_5540), .Z1_t (new_AGEMA_signal_5541), .Z1_f (new_AGEMA_signal_5542) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_33_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[33]), .A0_f (new_AGEMA_signal_15776), .A1_t (new_AGEMA_signal_15777), .A1_f (new_AGEMA_signal_15778), .B0_t (key_s0_t[33]), .B0_f (key_s0_f[33]), .B1_t (key_s1_t[33]), .B1_f (key_s1_f[33]), .Z0_t (KeyReg_Inst_ff_SDE_33_MUX_inst_X), .Z0_f (new_AGEMA_signal_16220), .Z1_t (new_AGEMA_signal_16221), .Z1_f (new_AGEMA_signal_16222) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_33_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_33_MUX_inst_X), .B0_f (new_AGEMA_signal_16220), .B1_t (new_AGEMA_signal_16221), .B1_f (new_AGEMA_signal_16222), .Z0_t (KeyReg_Inst_ff_SDE_33_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17096), .Z1_t (new_AGEMA_signal_17097), .Z1_f (new_AGEMA_signal_17098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_33_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_33_MUX_inst_Y), .A0_f (new_AGEMA_signal_17096), .A1_t (new_AGEMA_signal_17097), .A1_f (new_AGEMA_signal_17098), .B0_t (KeyExpansionOutput[33]), .B0_f (new_AGEMA_signal_15776), .B1_t (new_AGEMA_signal_15777), .B1_f (new_AGEMA_signal_15778), .Z0_t (RoundKey[33]), .Z0_f (new_AGEMA_signal_5549), .Z1_t (new_AGEMA_signal_5550), .Z1_f (new_AGEMA_signal_5551) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_34_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[34]), .A0_f (new_AGEMA_signal_15743), .A1_t (new_AGEMA_signal_15744), .A1_f (new_AGEMA_signal_15745), .B0_t (key_s0_t[34]), .B0_f (key_s0_f[34]), .B1_t (key_s1_t[34]), .B1_f (key_s1_f[34]), .Z0_t (KeyReg_Inst_ff_SDE_34_MUX_inst_X), .Z0_f (new_AGEMA_signal_16226), .Z1_t (new_AGEMA_signal_16227), .Z1_f (new_AGEMA_signal_16228) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_34_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_34_MUX_inst_X), .B0_f (new_AGEMA_signal_16226), .B1_t (new_AGEMA_signal_16227), .B1_f (new_AGEMA_signal_16228), .Z0_t (KeyReg_Inst_ff_SDE_34_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17099), .Z1_t (new_AGEMA_signal_17100), .Z1_f (new_AGEMA_signal_17101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_34_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_34_MUX_inst_Y), .A0_f (new_AGEMA_signal_17099), .A1_t (new_AGEMA_signal_17100), .A1_f (new_AGEMA_signal_17101), .B0_t (KeyExpansionOutput[34]), .B0_f (new_AGEMA_signal_15743), .B1_t (new_AGEMA_signal_15744), .B1_f (new_AGEMA_signal_15745), .Z0_t (RoundKey[34]), .Z0_f (new_AGEMA_signal_5558), .Z1_t (new_AGEMA_signal_5559), .Z1_f (new_AGEMA_signal_5560) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_35_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[35]), .A0_f (new_AGEMA_signal_15734), .A1_t (new_AGEMA_signal_15735), .A1_f (new_AGEMA_signal_15736), .B0_t (key_s0_t[35]), .B0_f (key_s0_f[35]), .B1_t (key_s1_t[35]), .B1_f (key_s1_f[35]), .Z0_t (KeyReg_Inst_ff_SDE_35_MUX_inst_X), .Z0_f (new_AGEMA_signal_16232), .Z1_t (new_AGEMA_signal_16233), .Z1_f (new_AGEMA_signal_16234) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_35_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_35_MUX_inst_X), .B0_f (new_AGEMA_signal_16232), .B1_t (new_AGEMA_signal_16233), .B1_f (new_AGEMA_signal_16234), .Z0_t (KeyReg_Inst_ff_SDE_35_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17102), .Z1_t (new_AGEMA_signal_17103), .Z1_f (new_AGEMA_signal_17104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_35_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_35_MUX_inst_Y), .A0_f (new_AGEMA_signal_17102), .A1_t (new_AGEMA_signal_17103), .A1_f (new_AGEMA_signal_17104), .B0_t (KeyExpansionOutput[35]), .B0_f (new_AGEMA_signal_15734), .B1_t (new_AGEMA_signal_15735), .B1_f (new_AGEMA_signal_15736), .Z0_t (RoundKey[35]), .Z0_f (new_AGEMA_signal_5567), .Z1_t (new_AGEMA_signal_5568), .Z1_f (new_AGEMA_signal_5569) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_36_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[36]), .A0_f (new_AGEMA_signal_15731), .A1_t (new_AGEMA_signal_15732), .A1_f (new_AGEMA_signal_15733), .B0_t (key_s0_t[36]), .B0_f (key_s0_f[36]), .B1_t (key_s1_t[36]), .B1_f (key_s1_f[36]), .Z0_t (KeyReg_Inst_ff_SDE_36_MUX_inst_X), .Z0_f (new_AGEMA_signal_16238), .Z1_t (new_AGEMA_signal_16239), .Z1_f (new_AGEMA_signal_16240) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_36_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_36_MUX_inst_X), .B0_f (new_AGEMA_signal_16238), .B1_t (new_AGEMA_signal_16239), .B1_f (new_AGEMA_signal_16240), .Z0_t (KeyReg_Inst_ff_SDE_36_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17105), .Z1_t (new_AGEMA_signal_17106), .Z1_f (new_AGEMA_signal_17107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_36_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_36_MUX_inst_Y), .A0_f (new_AGEMA_signal_17105), .A1_t (new_AGEMA_signal_17106), .A1_f (new_AGEMA_signal_17107), .B0_t (KeyExpansionOutput[36]), .B0_f (new_AGEMA_signal_15731), .B1_t (new_AGEMA_signal_15732), .B1_f (new_AGEMA_signal_15733), .Z0_t (RoundKey[36]), .Z0_f (new_AGEMA_signal_5576), .Z1_t (new_AGEMA_signal_5577), .Z1_f (new_AGEMA_signal_5578) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_37_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[37]), .A0_f (new_AGEMA_signal_15728), .A1_t (new_AGEMA_signal_15729), .A1_f (new_AGEMA_signal_15730), .B0_t (key_s0_t[37]), .B0_f (key_s0_f[37]), .B1_t (key_s1_t[37]), .B1_f (key_s1_f[37]), .Z0_t (KeyReg_Inst_ff_SDE_37_MUX_inst_X), .Z0_f (new_AGEMA_signal_16244), .Z1_t (new_AGEMA_signal_16245), .Z1_f (new_AGEMA_signal_16246) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_37_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_37_MUX_inst_X), .B0_f (new_AGEMA_signal_16244), .B1_t (new_AGEMA_signal_16245), .B1_f (new_AGEMA_signal_16246), .Z0_t (KeyReg_Inst_ff_SDE_37_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17108), .Z1_t (new_AGEMA_signal_17109), .Z1_f (new_AGEMA_signal_17110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_37_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_37_MUX_inst_Y), .A0_f (new_AGEMA_signal_17108), .A1_t (new_AGEMA_signal_17109), .A1_f (new_AGEMA_signal_17110), .B0_t (KeyExpansionOutput[37]), .B0_f (new_AGEMA_signal_15728), .B1_t (new_AGEMA_signal_15729), .B1_f (new_AGEMA_signal_15730), .Z0_t (RoundKey[37]), .Z0_f (new_AGEMA_signal_5585), .Z1_t (new_AGEMA_signal_5586), .Z1_f (new_AGEMA_signal_5587) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_38_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[38]), .A0_f (new_AGEMA_signal_15725), .A1_t (new_AGEMA_signal_15726), .A1_f (new_AGEMA_signal_15727), .B0_t (key_s0_t[38]), .B0_f (key_s0_f[38]), .B1_t (key_s1_t[38]), .B1_f (key_s1_f[38]), .Z0_t (KeyReg_Inst_ff_SDE_38_MUX_inst_X), .Z0_f (new_AGEMA_signal_16250), .Z1_t (new_AGEMA_signal_16251), .Z1_f (new_AGEMA_signal_16252) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_38_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_38_MUX_inst_X), .B0_f (new_AGEMA_signal_16250), .B1_t (new_AGEMA_signal_16251), .B1_f (new_AGEMA_signal_16252), .Z0_t (KeyReg_Inst_ff_SDE_38_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17111), .Z1_t (new_AGEMA_signal_17112), .Z1_f (new_AGEMA_signal_17113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_38_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_38_MUX_inst_Y), .A0_f (new_AGEMA_signal_17111), .A1_t (new_AGEMA_signal_17112), .A1_f (new_AGEMA_signal_17113), .B0_t (KeyExpansionOutput[38]), .B0_f (new_AGEMA_signal_15725), .B1_t (new_AGEMA_signal_15726), .B1_f (new_AGEMA_signal_15727), .Z0_t (RoundKey[38]), .Z0_f (new_AGEMA_signal_5594), .Z1_t (new_AGEMA_signal_5595), .Z1_f (new_AGEMA_signal_5596) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_39_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[39]), .A0_f (new_AGEMA_signal_15722), .A1_t (new_AGEMA_signal_15723), .A1_f (new_AGEMA_signal_15724), .B0_t (key_s0_t[39]), .B0_f (key_s0_f[39]), .B1_t (key_s1_t[39]), .B1_f (key_s1_f[39]), .Z0_t (KeyReg_Inst_ff_SDE_39_MUX_inst_X), .Z0_f (new_AGEMA_signal_16256), .Z1_t (new_AGEMA_signal_16257), .Z1_f (new_AGEMA_signal_16258) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_39_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_39_MUX_inst_X), .B0_f (new_AGEMA_signal_16256), .B1_t (new_AGEMA_signal_16257), .B1_f (new_AGEMA_signal_16258), .Z0_t (KeyReg_Inst_ff_SDE_39_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17114), .Z1_t (new_AGEMA_signal_17115), .Z1_f (new_AGEMA_signal_17116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_39_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_39_MUX_inst_Y), .A0_f (new_AGEMA_signal_17114), .A1_t (new_AGEMA_signal_17115), .A1_f (new_AGEMA_signal_17116), .B0_t (KeyExpansionOutput[39]), .B0_f (new_AGEMA_signal_15722), .B1_t (new_AGEMA_signal_15723), .B1_f (new_AGEMA_signal_15724), .Z0_t (RoundKey[39]), .Z0_f (new_AGEMA_signal_5603), .Z1_t (new_AGEMA_signal_5604), .Z1_f (new_AGEMA_signal_5605) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_40_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[40]), .A0_f (new_AGEMA_signal_14972), .A1_t (new_AGEMA_signal_14973), .A1_f (new_AGEMA_signal_14974), .B0_t (key_s0_t[40]), .B0_f (key_s0_f[40]), .B1_t (key_s1_t[40]), .B1_f (key_s1_f[40]), .Z0_t (KeyReg_Inst_ff_SDE_40_MUX_inst_X), .Z0_f (new_AGEMA_signal_15458), .Z1_t (new_AGEMA_signal_15459), .Z1_f (new_AGEMA_signal_15460) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_40_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_40_MUX_inst_X), .B0_f (new_AGEMA_signal_15458), .B1_t (new_AGEMA_signal_15459), .B1_f (new_AGEMA_signal_15460), .Z0_t (KeyReg_Inst_ff_SDE_40_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16259), .Z1_t (new_AGEMA_signal_16260), .Z1_f (new_AGEMA_signal_16261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_40_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_40_MUX_inst_Y), .A0_f (new_AGEMA_signal_16259), .A1_t (new_AGEMA_signal_16260), .A1_f (new_AGEMA_signal_16261), .B0_t (KeyExpansionOutput[40]), .B0_f (new_AGEMA_signal_14972), .B1_t (new_AGEMA_signal_14973), .B1_f (new_AGEMA_signal_14974), .Z0_t (RoundKey[40]), .Z0_f (new_AGEMA_signal_5621), .Z1_t (new_AGEMA_signal_5622), .Z1_f (new_AGEMA_signal_5623) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_41_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[41]), .A0_f (new_AGEMA_signal_15719), .A1_t (new_AGEMA_signal_15720), .A1_f (new_AGEMA_signal_15721), .B0_t (key_s0_t[41]), .B0_f (key_s0_f[41]), .B1_t (key_s1_t[41]), .B1_f (key_s1_f[41]), .Z0_t (KeyReg_Inst_ff_SDE_41_MUX_inst_X), .Z0_f (new_AGEMA_signal_16265), .Z1_t (new_AGEMA_signal_16266), .Z1_f (new_AGEMA_signal_16267) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_41_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_41_MUX_inst_X), .B0_f (new_AGEMA_signal_16265), .B1_t (new_AGEMA_signal_16266), .B1_f (new_AGEMA_signal_16267), .Z0_t (KeyReg_Inst_ff_SDE_41_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17117), .Z1_t (new_AGEMA_signal_17118), .Z1_f (new_AGEMA_signal_17119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_41_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_41_MUX_inst_Y), .A0_f (new_AGEMA_signal_17117), .A1_t (new_AGEMA_signal_17118), .A1_f (new_AGEMA_signal_17119), .B0_t (KeyExpansionOutput[41]), .B0_f (new_AGEMA_signal_15719), .B1_t (new_AGEMA_signal_15720), .B1_f (new_AGEMA_signal_15721), .Z0_t (RoundKey[41]), .Z0_f (new_AGEMA_signal_5630), .Z1_t (new_AGEMA_signal_5631), .Z1_f (new_AGEMA_signal_5632) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_42_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[42]), .A0_f (new_AGEMA_signal_15806), .A1_t (new_AGEMA_signal_15807), .A1_f (new_AGEMA_signal_15808), .B0_t (key_s0_t[42]), .B0_f (key_s0_f[42]), .B1_t (key_s1_t[42]), .B1_f (key_s1_f[42]), .Z0_t (KeyReg_Inst_ff_SDE_42_MUX_inst_X), .Z0_f (new_AGEMA_signal_16271), .Z1_t (new_AGEMA_signal_16272), .Z1_f (new_AGEMA_signal_16273) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_42_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_42_MUX_inst_X), .B0_f (new_AGEMA_signal_16271), .B1_t (new_AGEMA_signal_16272), .B1_f (new_AGEMA_signal_16273), .Z0_t (KeyReg_Inst_ff_SDE_42_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17120), .Z1_t (new_AGEMA_signal_17121), .Z1_f (new_AGEMA_signal_17122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_42_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_42_MUX_inst_Y), .A0_f (new_AGEMA_signal_17120), .A1_t (new_AGEMA_signal_17121), .A1_f (new_AGEMA_signal_17122), .B0_t (KeyExpansionOutput[42]), .B0_f (new_AGEMA_signal_15806), .B1_t (new_AGEMA_signal_15807), .B1_f (new_AGEMA_signal_15808), .Z0_t (RoundKey[42]), .Z0_f (new_AGEMA_signal_5639), .Z1_t (new_AGEMA_signal_5640), .Z1_f (new_AGEMA_signal_5641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_43_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[43]), .A0_f (new_AGEMA_signal_15803), .A1_t (new_AGEMA_signal_15804), .A1_f (new_AGEMA_signal_15805), .B0_t (key_s0_t[43]), .B0_f (key_s0_f[43]), .B1_t (key_s1_t[43]), .B1_f (key_s1_f[43]), .Z0_t (KeyReg_Inst_ff_SDE_43_MUX_inst_X), .Z0_f (new_AGEMA_signal_16277), .Z1_t (new_AGEMA_signal_16278), .Z1_f (new_AGEMA_signal_16279) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_43_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_43_MUX_inst_X), .B0_f (new_AGEMA_signal_16277), .B1_t (new_AGEMA_signal_16278), .B1_f (new_AGEMA_signal_16279), .Z0_t (KeyReg_Inst_ff_SDE_43_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17123), .Z1_t (new_AGEMA_signal_17124), .Z1_f (new_AGEMA_signal_17125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_43_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_43_MUX_inst_Y), .A0_f (new_AGEMA_signal_17123), .A1_t (new_AGEMA_signal_17124), .A1_f (new_AGEMA_signal_17125), .B0_t (KeyExpansionOutput[43]), .B0_f (new_AGEMA_signal_15803), .B1_t (new_AGEMA_signal_15804), .B1_f (new_AGEMA_signal_15805), .Z0_t (RoundKey[43]), .Z0_f (new_AGEMA_signal_5648), .Z1_t (new_AGEMA_signal_5649), .Z1_f (new_AGEMA_signal_5650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_44_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[44]), .A0_f (new_AGEMA_signal_15800), .A1_t (new_AGEMA_signal_15801), .A1_f (new_AGEMA_signal_15802), .B0_t (key_s0_t[44]), .B0_f (key_s0_f[44]), .B1_t (key_s1_t[44]), .B1_f (key_s1_f[44]), .Z0_t (KeyReg_Inst_ff_SDE_44_MUX_inst_X), .Z0_f (new_AGEMA_signal_16283), .Z1_t (new_AGEMA_signal_16284), .Z1_f (new_AGEMA_signal_16285) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_44_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_44_MUX_inst_X), .B0_f (new_AGEMA_signal_16283), .B1_t (new_AGEMA_signal_16284), .B1_f (new_AGEMA_signal_16285), .Z0_t (KeyReg_Inst_ff_SDE_44_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17126), .Z1_t (new_AGEMA_signal_17127), .Z1_f (new_AGEMA_signal_17128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_44_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_44_MUX_inst_Y), .A0_f (new_AGEMA_signal_17126), .A1_t (new_AGEMA_signal_17127), .A1_f (new_AGEMA_signal_17128), .B0_t (KeyExpansionOutput[44]), .B0_f (new_AGEMA_signal_15800), .B1_t (new_AGEMA_signal_15801), .B1_f (new_AGEMA_signal_15802), .Z0_t (RoundKey[44]), .Z0_f (new_AGEMA_signal_5657), .Z1_t (new_AGEMA_signal_5658), .Z1_f (new_AGEMA_signal_5659) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_45_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[45]), .A0_f (new_AGEMA_signal_15797), .A1_t (new_AGEMA_signal_15798), .A1_f (new_AGEMA_signal_15799), .B0_t (key_s0_t[45]), .B0_f (key_s0_f[45]), .B1_t (key_s1_t[45]), .B1_f (key_s1_f[45]), .Z0_t (KeyReg_Inst_ff_SDE_45_MUX_inst_X), .Z0_f (new_AGEMA_signal_16289), .Z1_t (new_AGEMA_signal_16290), .Z1_f (new_AGEMA_signal_16291) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_45_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_45_MUX_inst_X), .B0_f (new_AGEMA_signal_16289), .B1_t (new_AGEMA_signal_16290), .B1_f (new_AGEMA_signal_16291), .Z0_t (KeyReg_Inst_ff_SDE_45_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17129), .Z1_t (new_AGEMA_signal_17130), .Z1_f (new_AGEMA_signal_17131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_45_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_45_MUX_inst_Y), .A0_f (new_AGEMA_signal_17129), .A1_t (new_AGEMA_signal_17130), .A1_f (new_AGEMA_signal_17131), .B0_t (KeyExpansionOutput[45]), .B0_f (new_AGEMA_signal_15797), .B1_t (new_AGEMA_signal_15798), .B1_f (new_AGEMA_signal_15799), .Z0_t (RoundKey[45]), .Z0_f (new_AGEMA_signal_5666), .Z1_t (new_AGEMA_signal_5667), .Z1_f (new_AGEMA_signal_5668) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_46_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[46]), .A0_f (new_AGEMA_signal_15794), .A1_t (new_AGEMA_signal_15795), .A1_f (new_AGEMA_signal_15796), .B0_t (key_s0_t[46]), .B0_f (key_s0_f[46]), .B1_t (key_s1_t[46]), .B1_f (key_s1_f[46]), .Z0_t (KeyReg_Inst_ff_SDE_46_MUX_inst_X), .Z0_f (new_AGEMA_signal_16295), .Z1_t (new_AGEMA_signal_16296), .Z1_f (new_AGEMA_signal_16297) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_46_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_46_MUX_inst_X), .B0_f (new_AGEMA_signal_16295), .B1_t (new_AGEMA_signal_16296), .B1_f (new_AGEMA_signal_16297), .Z0_t (KeyReg_Inst_ff_SDE_46_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17132), .Z1_t (new_AGEMA_signal_17133), .Z1_f (new_AGEMA_signal_17134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_46_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_46_MUX_inst_Y), .A0_f (new_AGEMA_signal_17132), .A1_t (new_AGEMA_signal_17133), .A1_f (new_AGEMA_signal_17134), .B0_t (KeyExpansionOutput[46]), .B0_f (new_AGEMA_signal_15794), .B1_t (new_AGEMA_signal_15795), .B1_f (new_AGEMA_signal_15796), .Z0_t (RoundKey[46]), .Z0_f (new_AGEMA_signal_5675), .Z1_t (new_AGEMA_signal_5676), .Z1_f (new_AGEMA_signal_5677) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_47_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[47]), .A0_f (new_AGEMA_signal_15791), .A1_t (new_AGEMA_signal_15792), .A1_f (new_AGEMA_signal_15793), .B0_t (key_s0_t[47]), .B0_f (key_s0_f[47]), .B1_t (key_s1_t[47]), .B1_f (key_s1_f[47]), .Z0_t (KeyReg_Inst_ff_SDE_47_MUX_inst_X), .Z0_f (new_AGEMA_signal_16301), .Z1_t (new_AGEMA_signal_16302), .Z1_f (new_AGEMA_signal_16303) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_47_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_47_MUX_inst_X), .B0_f (new_AGEMA_signal_16301), .B1_t (new_AGEMA_signal_16302), .B1_f (new_AGEMA_signal_16303), .Z0_t (KeyReg_Inst_ff_SDE_47_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17135), .Z1_t (new_AGEMA_signal_17136), .Z1_f (new_AGEMA_signal_17137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_47_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_47_MUX_inst_Y), .A0_f (new_AGEMA_signal_17135), .A1_t (new_AGEMA_signal_17136), .A1_f (new_AGEMA_signal_17137), .B0_t (KeyExpansionOutput[47]), .B0_f (new_AGEMA_signal_15791), .B1_t (new_AGEMA_signal_15792), .B1_f (new_AGEMA_signal_15793), .Z0_t (RoundKey[47]), .Z0_f (new_AGEMA_signal_5684), .Z1_t (new_AGEMA_signal_5685), .Z1_f (new_AGEMA_signal_5686) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_48_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[48]), .A0_f (new_AGEMA_signal_15020), .A1_t (new_AGEMA_signal_15021), .A1_f (new_AGEMA_signal_15022), .B0_t (key_s0_t[48]), .B0_f (key_s0_f[48]), .B1_t (key_s1_t[48]), .B1_f (key_s1_f[48]), .Z0_t (KeyReg_Inst_ff_SDE_48_MUX_inst_X), .Z0_f (new_AGEMA_signal_15464), .Z1_t (new_AGEMA_signal_15465), .Z1_f (new_AGEMA_signal_15466) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_48_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_48_MUX_inst_X), .B0_f (new_AGEMA_signal_15464), .B1_t (new_AGEMA_signal_15465), .B1_f (new_AGEMA_signal_15466), .Z0_t (KeyReg_Inst_ff_SDE_48_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16304), .Z1_t (new_AGEMA_signal_16305), .Z1_f (new_AGEMA_signal_16306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_48_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_48_MUX_inst_Y), .A0_f (new_AGEMA_signal_16304), .A1_t (new_AGEMA_signal_16305), .A1_f (new_AGEMA_signal_16306), .B0_t (KeyExpansionOutput[48]), .B0_f (new_AGEMA_signal_15020), .B1_t (new_AGEMA_signal_15021), .B1_f (new_AGEMA_signal_15022), .Z0_t (RoundKey[48]), .Z0_f (new_AGEMA_signal_5693), .Z1_t (new_AGEMA_signal_5694), .Z1_f (new_AGEMA_signal_5695) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_49_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[49]), .A0_f (new_AGEMA_signal_15785), .A1_t (new_AGEMA_signal_15786), .A1_f (new_AGEMA_signal_15787), .B0_t (key_s0_t[49]), .B0_f (key_s0_f[49]), .B1_t (key_s1_t[49]), .B1_f (key_s1_f[49]), .Z0_t (KeyReg_Inst_ff_SDE_49_MUX_inst_X), .Z0_f (new_AGEMA_signal_16310), .Z1_t (new_AGEMA_signal_16311), .Z1_f (new_AGEMA_signal_16312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_49_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_49_MUX_inst_X), .B0_f (new_AGEMA_signal_16310), .B1_t (new_AGEMA_signal_16311), .B1_f (new_AGEMA_signal_16312), .Z0_t (KeyReg_Inst_ff_SDE_49_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17138), .Z1_t (new_AGEMA_signal_17139), .Z1_f (new_AGEMA_signal_17140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_49_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_49_MUX_inst_Y), .A0_f (new_AGEMA_signal_17138), .A1_t (new_AGEMA_signal_17139), .A1_f (new_AGEMA_signal_17140), .B0_t (KeyExpansionOutput[49]), .B0_f (new_AGEMA_signal_15785), .B1_t (new_AGEMA_signal_15786), .B1_f (new_AGEMA_signal_15787), .Z0_t (RoundKey[49]), .Z0_f (new_AGEMA_signal_5702), .Z1_t (new_AGEMA_signal_5703), .Z1_f (new_AGEMA_signal_5704) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_50_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[50]), .A0_f (new_AGEMA_signal_15782), .A1_t (new_AGEMA_signal_15783), .A1_f (new_AGEMA_signal_15784), .B0_t (key_s0_t[50]), .B0_f (key_s0_f[50]), .B1_t (key_s1_t[50]), .B1_f (key_s1_f[50]), .Z0_t (KeyReg_Inst_ff_SDE_50_MUX_inst_X), .Z0_f (new_AGEMA_signal_16316), .Z1_t (new_AGEMA_signal_16317), .Z1_f (new_AGEMA_signal_16318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_50_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_50_MUX_inst_X), .B0_f (new_AGEMA_signal_16316), .B1_t (new_AGEMA_signal_16317), .B1_f (new_AGEMA_signal_16318), .Z0_t (KeyReg_Inst_ff_SDE_50_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17141), .Z1_t (new_AGEMA_signal_17142), .Z1_f (new_AGEMA_signal_17143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_50_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_50_MUX_inst_Y), .A0_f (new_AGEMA_signal_17141), .A1_t (new_AGEMA_signal_17142), .A1_f (new_AGEMA_signal_17143), .B0_t (KeyExpansionOutput[50]), .B0_f (new_AGEMA_signal_15782), .B1_t (new_AGEMA_signal_15783), .B1_f (new_AGEMA_signal_15784), .Z0_t (RoundKey[50]), .Z0_f (new_AGEMA_signal_5720), .Z1_t (new_AGEMA_signal_5721), .Z1_f (new_AGEMA_signal_5722) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_51_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[51]), .A0_f (new_AGEMA_signal_15779), .A1_t (new_AGEMA_signal_15780), .A1_f (new_AGEMA_signal_15781), .B0_t (key_s0_t[51]), .B0_f (key_s0_f[51]), .B1_t (key_s1_t[51]), .B1_f (key_s1_f[51]), .Z0_t (KeyReg_Inst_ff_SDE_51_MUX_inst_X), .Z0_f (new_AGEMA_signal_16322), .Z1_t (new_AGEMA_signal_16323), .Z1_f (new_AGEMA_signal_16324) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_51_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_51_MUX_inst_X), .B0_f (new_AGEMA_signal_16322), .B1_t (new_AGEMA_signal_16323), .B1_f (new_AGEMA_signal_16324), .Z0_t (KeyReg_Inst_ff_SDE_51_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17144), .Z1_t (new_AGEMA_signal_17145), .Z1_f (new_AGEMA_signal_17146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_51_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_51_MUX_inst_Y), .A0_f (new_AGEMA_signal_17144), .A1_t (new_AGEMA_signal_17145), .A1_f (new_AGEMA_signal_17146), .B0_t (KeyExpansionOutput[51]), .B0_f (new_AGEMA_signal_15779), .B1_t (new_AGEMA_signal_15780), .B1_f (new_AGEMA_signal_15781), .Z0_t (RoundKey[51]), .Z0_f (new_AGEMA_signal_5729), .Z1_t (new_AGEMA_signal_5730), .Z1_f (new_AGEMA_signal_5731) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_52_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[52]), .A0_f (new_AGEMA_signal_15773), .A1_t (new_AGEMA_signal_15774), .A1_f (new_AGEMA_signal_15775), .B0_t (key_s0_t[52]), .B0_f (key_s0_f[52]), .B1_t (key_s1_t[52]), .B1_f (key_s1_f[52]), .Z0_t (KeyReg_Inst_ff_SDE_52_MUX_inst_X), .Z0_f (new_AGEMA_signal_16328), .Z1_t (new_AGEMA_signal_16329), .Z1_f (new_AGEMA_signal_16330) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_52_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_52_MUX_inst_X), .B0_f (new_AGEMA_signal_16328), .B1_t (new_AGEMA_signal_16329), .B1_f (new_AGEMA_signal_16330), .Z0_t (KeyReg_Inst_ff_SDE_52_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17147), .Z1_t (new_AGEMA_signal_17148), .Z1_f (new_AGEMA_signal_17149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_52_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_52_MUX_inst_Y), .A0_f (new_AGEMA_signal_17147), .A1_t (new_AGEMA_signal_17148), .A1_f (new_AGEMA_signal_17149), .B0_t (KeyExpansionOutput[52]), .B0_f (new_AGEMA_signal_15773), .B1_t (new_AGEMA_signal_15774), .B1_f (new_AGEMA_signal_15775), .Z0_t (RoundKey[52]), .Z0_f (new_AGEMA_signal_5738), .Z1_t (new_AGEMA_signal_5739), .Z1_f (new_AGEMA_signal_5740) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_53_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[53]), .A0_f (new_AGEMA_signal_15770), .A1_t (new_AGEMA_signal_15771), .A1_f (new_AGEMA_signal_15772), .B0_t (key_s0_t[53]), .B0_f (key_s0_f[53]), .B1_t (key_s1_t[53]), .B1_f (key_s1_f[53]), .Z0_t (KeyReg_Inst_ff_SDE_53_MUX_inst_X), .Z0_f (new_AGEMA_signal_16334), .Z1_t (new_AGEMA_signal_16335), .Z1_f (new_AGEMA_signal_16336) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_53_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_53_MUX_inst_X), .B0_f (new_AGEMA_signal_16334), .B1_t (new_AGEMA_signal_16335), .B1_f (new_AGEMA_signal_16336), .Z0_t (KeyReg_Inst_ff_SDE_53_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17150), .Z1_t (new_AGEMA_signal_17151), .Z1_f (new_AGEMA_signal_17152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_53_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_53_MUX_inst_Y), .A0_f (new_AGEMA_signal_17150), .A1_t (new_AGEMA_signal_17151), .A1_f (new_AGEMA_signal_17152), .B0_t (KeyExpansionOutput[53]), .B0_f (new_AGEMA_signal_15770), .B1_t (new_AGEMA_signal_15771), .B1_f (new_AGEMA_signal_15772), .Z0_t (RoundKey[53]), .Z0_f (new_AGEMA_signal_5747), .Z1_t (new_AGEMA_signal_5748), .Z1_f (new_AGEMA_signal_5749) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_54_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[54]), .A0_f (new_AGEMA_signal_15767), .A1_t (new_AGEMA_signal_15768), .A1_f (new_AGEMA_signal_15769), .B0_t (key_s0_t[54]), .B0_f (key_s0_f[54]), .B1_t (key_s1_t[54]), .B1_f (key_s1_f[54]), .Z0_t (KeyReg_Inst_ff_SDE_54_MUX_inst_X), .Z0_f (new_AGEMA_signal_16340), .Z1_t (new_AGEMA_signal_16341), .Z1_f (new_AGEMA_signal_16342) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_54_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_54_MUX_inst_X), .B0_f (new_AGEMA_signal_16340), .B1_t (new_AGEMA_signal_16341), .B1_f (new_AGEMA_signal_16342), .Z0_t (KeyReg_Inst_ff_SDE_54_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17153), .Z1_t (new_AGEMA_signal_17154), .Z1_f (new_AGEMA_signal_17155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_54_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_54_MUX_inst_Y), .A0_f (new_AGEMA_signal_17153), .A1_t (new_AGEMA_signal_17154), .A1_f (new_AGEMA_signal_17155), .B0_t (KeyExpansionOutput[54]), .B0_f (new_AGEMA_signal_15767), .B1_t (new_AGEMA_signal_15768), .B1_f (new_AGEMA_signal_15769), .Z0_t (RoundKey[54]), .Z0_f (new_AGEMA_signal_5756), .Z1_t (new_AGEMA_signal_5757), .Z1_f (new_AGEMA_signal_5758) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_55_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[55]), .A0_f (new_AGEMA_signal_15764), .A1_t (new_AGEMA_signal_15765), .A1_f (new_AGEMA_signal_15766), .B0_t (key_s0_t[55]), .B0_f (key_s0_f[55]), .B1_t (key_s1_t[55]), .B1_f (key_s1_f[55]), .Z0_t (KeyReg_Inst_ff_SDE_55_MUX_inst_X), .Z0_f (new_AGEMA_signal_16346), .Z1_t (new_AGEMA_signal_16347), .Z1_f (new_AGEMA_signal_16348) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_55_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_55_MUX_inst_X), .B0_f (new_AGEMA_signal_16346), .B1_t (new_AGEMA_signal_16347), .B1_f (new_AGEMA_signal_16348), .Z0_t (KeyReg_Inst_ff_SDE_55_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17156), .Z1_t (new_AGEMA_signal_17157), .Z1_f (new_AGEMA_signal_17158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_55_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_55_MUX_inst_Y), .A0_f (new_AGEMA_signal_17156), .A1_t (new_AGEMA_signal_17157), .A1_f (new_AGEMA_signal_17158), .B0_t (KeyExpansionOutput[55]), .B0_f (new_AGEMA_signal_15764), .B1_t (new_AGEMA_signal_15765), .B1_f (new_AGEMA_signal_15766), .Z0_t (RoundKey[55]), .Z0_f (new_AGEMA_signal_5765), .Z1_t (new_AGEMA_signal_5766), .Z1_f (new_AGEMA_signal_5767) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_56_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[56]), .A0_f (new_AGEMA_signal_15761), .A1_t (new_AGEMA_signal_15762), .A1_f (new_AGEMA_signal_15763), .B0_t (key_s0_t[56]), .B0_f (key_s0_f[56]), .B1_t (key_s1_t[56]), .B1_f (key_s1_f[56]), .Z0_t (KeyReg_Inst_ff_SDE_56_MUX_inst_X), .Z0_f (new_AGEMA_signal_16352), .Z1_t (new_AGEMA_signal_16353), .Z1_f (new_AGEMA_signal_16354) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_56_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_56_MUX_inst_X), .B0_f (new_AGEMA_signal_16352), .B1_t (new_AGEMA_signal_16353), .B1_f (new_AGEMA_signal_16354), .Z0_t (KeyReg_Inst_ff_SDE_56_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17159), .Z1_t (new_AGEMA_signal_17160), .Z1_f (new_AGEMA_signal_17161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_56_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_56_MUX_inst_Y), .A0_f (new_AGEMA_signal_17159), .A1_t (new_AGEMA_signal_17160), .A1_f (new_AGEMA_signal_17161), .B0_t (KeyExpansionOutput[56]), .B0_f (new_AGEMA_signal_15761), .B1_t (new_AGEMA_signal_15762), .B1_f (new_AGEMA_signal_15763), .Z0_t (RoundKey[56]), .Z0_f (new_AGEMA_signal_5774), .Z1_t (new_AGEMA_signal_5775), .Z1_f (new_AGEMA_signal_5776) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_57_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[57]), .A0_f (new_AGEMA_signal_16523), .A1_t (new_AGEMA_signal_16524), .A1_f (new_AGEMA_signal_16525), .B0_t (key_s0_t[57]), .B0_f (key_s0_f[57]), .B1_t (key_s1_t[57]), .B1_f (key_s1_f[57]), .Z0_t (KeyReg_Inst_ff_SDE_57_MUX_inst_X), .Z0_f (new_AGEMA_signal_17165), .Z1_t (new_AGEMA_signal_17166), .Z1_f (new_AGEMA_signal_17167) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_57_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_57_MUX_inst_X), .B0_f (new_AGEMA_signal_17165), .B1_t (new_AGEMA_signal_17166), .B1_f (new_AGEMA_signal_17167), .Z0_t (KeyReg_Inst_ff_SDE_57_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17738), .Z1_t (new_AGEMA_signal_17739), .Z1_f (new_AGEMA_signal_17740) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_57_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_57_MUX_inst_Y), .A0_f (new_AGEMA_signal_17738), .A1_t (new_AGEMA_signal_17739), .A1_f (new_AGEMA_signal_17740), .B0_t (KeyExpansionOutput[57]), .B0_f (new_AGEMA_signal_16523), .B1_t (new_AGEMA_signal_16524), .B1_f (new_AGEMA_signal_16525), .Z0_t (RoundKey[57]), .Z0_f (new_AGEMA_signal_5783), .Z1_t (new_AGEMA_signal_5784), .Z1_f (new_AGEMA_signal_5785) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_58_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[58]), .A0_f (new_AGEMA_signal_16520), .A1_t (new_AGEMA_signal_16521), .A1_f (new_AGEMA_signal_16522), .B0_t (key_s0_t[58]), .B0_f (key_s0_f[58]), .B1_t (key_s1_t[58]), .B1_f (key_s1_f[58]), .Z0_t (KeyReg_Inst_ff_SDE_58_MUX_inst_X), .Z0_f (new_AGEMA_signal_17171), .Z1_t (new_AGEMA_signal_17172), .Z1_f (new_AGEMA_signal_17173) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_58_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_58_MUX_inst_X), .B0_f (new_AGEMA_signal_17171), .B1_t (new_AGEMA_signal_17172), .B1_f (new_AGEMA_signal_17173), .Z0_t (KeyReg_Inst_ff_SDE_58_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17741), .Z1_t (new_AGEMA_signal_17742), .Z1_f (new_AGEMA_signal_17743) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_58_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_58_MUX_inst_Y), .A0_f (new_AGEMA_signal_17741), .A1_t (new_AGEMA_signal_17742), .A1_f (new_AGEMA_signal_17743), .B0_t (KeyExpansionOutput[58]), .B0_f (new_AGEMA_signal_16520), .B1_t (new_AGEMA_signal_16521), .B1_f (new_AGEMA_signal_16522), .Z0_t (RoundKey[58]), .Z0_f (new_AGEMA_signal_5792), .Z1_t (new_AGEMA_signal_5793), .Z1_f (new_AGEMA_signal_5794) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_59_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[59]), .A0_f (new_AGEMA_signal_16517), .A1_t (new_AGEMA_signal_16518), .A1_f (new_AGEMA_signal_16519), .B0_t (key_s0_t[59]), .B0_f (key_s0_f[59]), .B1_t (key_s1_t[59]), .B1_f (key_s1_f[59]), .Z0_t (KeyReg_Inst_ff_SDE_59_MUX_inst_X), .Z0_f (new_AGEMA_signal_17177), .Z1_t (new_AGEMA_signal_17178), .Z1_f (new_AGEMA_signal_17179) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_59_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_59_MUX_inst_X), .B0_f (new_AGEMA_signal_17177), .B1_t (new_AGEMA_signal_17178), .B1_f (new_AGEMA_signal_17179), .Z0_t (KeyReg_Inst_ff_SDE_59_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17744), .Z1_t (new_AGEMA_signal_17745), .Z1_f (new_AGEMA_signal_17746) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_59_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_59_MUX_inst_Y), .A0_f (new_AGEMA_signal_17744), .A1_t (new_AGEMA_signal_17745), .A1_f (new_AGEMA_signal_17746), .B0_t (KeyExpansionOutput[59]), .B0_f (new_AGEMA_signal_16517), .B1_t (new_AGEMA_signal_16518), .B1_f (new_AGEMA_signal_16519), .Z0_t (RoundKey[59]), .Z0_f (new_AGEMA_signal_5801), .Z1_t (new_AGEMA_signal_5802), .Z1_f (new_AGEMA_signal_5803) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_60_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[60]), .A0_f (new_AGEMA_signal_16514), .A1_t (new_AGEMA_signal_16515), .A1_f (new_AGEMA_signal_16516), .B0_t (key_s0_t[60]), .B0_f (key_s0_f[60]), .B1_t (key_s1_t[60]), .B1_f (key_s1_f[60]), .Z0_t (KeyReg_Inst_ff_SDE_60_MUX_inst_X), .Z0_f (new_AGEMA_signal_17183), .Z1_t (new_AGEMA_signal_17184), .Z1_f (new_AGEMA_signal_17185) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_60_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_60_MUX_inst_X), .B0_f (new_AGEMA_signal_17183), .B1_t (new_AGEMA_signal_17184), .B1_f (new_AGEMA_signal_17185), .Z0_t (KeyReg_Inst_ff_SDE_60_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17747), .Z1_t (new_AGEMA_signal_17748), .Z1_f (new_AGEMA_signal_17749) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_60_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_60_MUX_inst_Y), .A0_f (new_AGEMA_signal_17747), .A1_t (new_AGEMA_signal_17748), .A1_f (new_AGEMA_signal_17749), .B0_t (KeyExpansionOutput[60]), .B0_f (new_AGEMA_signal_16514), .B1_t (new_AGEMA_signal_16515), .B1_f (new_AGEMA_signal_16516), .Z0_t (RoundKey[60]), .Z0_f (new_AGEMA_signal_5819), .Z1_t (new_AGEMA_signal_5820), .Z1_f (new_AGEMA_signal_5821) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_61_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[61]), .A0_f (new_AGEMA_signal_16511), .A1_t (new_AGEMA_signal_16512), .A1_f (new_AGEMA_signal_16513), .B0_t (key_s0_t[61]), .B0_f (key_s0_f[61]), .B1_t (key_s1_t[61]), .B1_f (key_s1_f[61]), .Z0_t (KeyReg_Inst_ff_SDE_61_MUX_inst_X), .Z0_f (new_AGEMA_signal_17189), .Z1_t (new_AGEMA_signal_17190), .Z1_f (new_AGEMA_signal_17191) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_61_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_61_MUX_inst_X), .B0_f (new_AGEMA_signal_17189), .B1_t (new_AGEMA_signal_17190), .B1_f (new_AGEMA_signal_17191), .Z0_t (KeyReg_Inst_ff_SDE_61_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17750), .Z1_t (new_AGEMA_signal_17751), .Z1_f (new_AGEMA_signal_17752) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_61_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_61_MUX_inst_Y), .A0_f (new_AGEMA_signal_17750), .A1_t (new_AGEMA_signal_17751), .A1_f (new_AGEMA_signal_17752), .B0_t (KeyExpansionOutput[61]), .B0_f (new_AGEMA_signal_16511), .B1_t (new_AGEMA_signal_16512), .B1_f (new_AGEMA_signal_16513), .Z0_t (RoundKey[61]), .Z0_f (new_AGEMA_signal_5828), .Z1_t (new_AGEMA_signal_5829), .Z1_f (new_AGEMA_signal_5830) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_62_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[62]), .A0_f (new_AGEMA_signal_16505), .A1_t (new_AGEMA_signal_16506), .A1_f (new_AGEMA_signal_16507), .B0_t (key_s0_t[62]), .B0_f (key_s0_f[62]), .B1_t (key_s1_t[62]), .B1_f (key_s1_f[62]), .Z0_t (KeyReg_Inst_ff_SDE_62_MUX_inst_X), .Z0_f (new_AGEMA_signal_17195), .Z1_t (new_AGEMA_signal_17196), .Z1_f (new_AGEMA_signal_17197) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_62_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_62_MUX_inst_X), .B0_f (new_AGEMA_signal_17195), .B1_t (new_AGEMA_signal_17196), .B1_f (new_AGEMA_signal_17197), .Z0_t (KeyReg_Inst_ff_SDE_62_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17753), .Z1_t (new_AGEMA_signal_17754), .Z1_f (new_AGEMA_signal_17755) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_62_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_62_MUX_inst_Y), .A0_f (new_AGEMA_signal_17753), .A1_t (new_AGEMA_signal_17754), .A1_f (new_AGEMA_signal_17755), .B0_t (KeyExpansionOutput[62]), .B0_f (new_AGEMA_signal_16505), .B1_t (new_AGEMA_signal_16506), .B1_f (new_AGEMA_signal_16507), .Z0_t (RoundKey[62]), .Z0_f (new_AGEMA_signal_5837), .Z1_t (new_AGEMA_signal_5838), .Z1_f (new_AGEMA_signal_5839) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_63_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[63]), .A0_f (new_AGEMA_signal_16502), .A1_t (new_AGEMA_signal_16503), .A1_f (new_AGEMA_signal_16504), .B0_t (key_s0_t[63]), .B0_f (key_s0_f[63]), .B1_t (key_s1_t[63]), .B1_f (key_s1_f[63]), .Z0_t (KeyReg_Inst_ff_SDE_63_MUX_inst_X), .Z0_f (new_AGEMA_signal_17201), .Z1_t (new_AGEMA_signal_17202), .Z1_f (new_AGEMA_signal_17203) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_63_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_63_MUX_inst_X), .B0_f (new_AGEMA_signal_17201), .B1_t (new_AGEMA_signal_17202), .B1_f (new_AGEMA_signal_17203), .Z0_t (KeyReg_Inst_ff_SDE_63_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17756), .Z1_t (new_AGEMA_signal_17757), .Z1_f (new_AGEMA_signal_17758) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_63_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_63_MUX_inst_Y), .A0_f (new_AGEMA_signal_17756), .A1_t (new_AGEMA_signal_17757), .A1_f (new_AGEMA_signal_17758), .B0_t (KeyExpansionOutput[63]), .B0_f (new_AGEMA_signal_16502), .B1_t (new_AGEMA_signal_16503), .B1_f (new_AGEMA_signal_16504), .Z0_t (RoundKey[63]), .Z0_f (new_AGEMA_signal_5846), .Z1_t (new_AGEMA_signal_5847), .Z1_f (new_AGEMA_signal_5848) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_64_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[64]), .A0_f (new_AGEMA_signal_14066), .A1_t (new_AGEMA_signal_14067), .A1_f (new_AGEMA_signal_14068), .B0_t (key_s0_t[64]), .B0_f (key_s0_f[64]), .B1_t (key_s1_t[64]), .B1_f (key_s1_f[64]), .Z0_t (KeyReg_Inst_ff_SDE_64_MUX_inst_X), .Z0_f (new_AGEMA_signal_14813), .Z1_t (new_AGEMA_signal_14814), .Z1_f (new_AGEMA_signal_14815) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_64_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_64_MUX_inst_X), .B0_f (new_AGEMA_signal_14813), .B1_t (new_AGEMA_signal_14814), .B1_f (new_AGEMA_signal_14815), .Z0_t (KeyReg_Inst_ff_SDE_64_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15467), .Z1_t (new_AGEMA_signal_15468), .Z1_f (new_AGEMA_signal_15469) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_64_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_64_MUX_inst_Y), .A0_f (new_AGEMA_signal_15467), .A1_t (new_AGEMA_signal_15468), .A1_f (new_AGEMA_signal_15469), .B0_t (KeyExpansionOutput[64]), .B0_f (new_AGEMA_signal_14066), .B1_t (new_AGEMA_signal_14067), .B1_f (new_AGEMA_signal_14068), .Z0_t (RoundKey[64]), .Z0_f (new_AGEMA_signal_5855), .Z1_t (new_AGEMA_signal_5856), .Z1_f (new_AGEMA_signal_5857) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_65_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[65]), .A0_f (new_AGEMA_signal_15008), .A1_t (new_AGEMA_signal_15009), .A1_f (new_AGEMA_signal_15010), .B0_t (key_s0_t[65]), .B0_f (key_s0_f[65]), .B1_t (key_s1_t[65]), .B1_f (key_s1_f[65]), .Z0_t (KeyReg_Inst_ff_SDE_65_MUX_inst_X), .Z0_f (new_AGEMA_signal_15473), .Z1_t (new_AGEMA_signal_15474), .Z1_f (new_AGEMA_signal_15475) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_65_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_65_MUX_inst_X), .B0_f (new_AGEMA_signal_15473), .B1_t (new_AGEMA_signal_15474), .B1_f (new_AGEMA_signal_15475), .Z0_t (KeyReg_Inst_ff_SDE_65_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16355), .Z1_t (new_AGEMA_signal_16356), .Z1_f (new_AGEMA_signal_16357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_65_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_65_MUX_inst_Y), .A0_f (new_AGEMA_signal_16355), .A1_t (new_AGEMA_signal_16356), .A1_f (new_AGEMA_signal_16357), .B0_t (KeyExpansionOutput[65]), .B0_f (new_AGEMA_signal_15008), .B1_t (new_AGEMA_signal_15009), .B1_f (new_AGEMA_signal_15010), .Z0_t (RoundKey[65]), .Z0_f (new_AGEMA_signal_5864), .Z1_t (new_AGEMA_signal_5865), .Z1_f (new_AGEMA_signal_5866) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_66_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[66]), .A0_f (new_AGEMA_signal_14990), .A1_t (new_AGEMA_signal_14991), .A1_f (new_AGEMA_signal_14992), .B0_t (key_s0_t[66]), .B0_f (key_s0_f[66]), .B1_t (key_s1_t[66]), .B1_f (key_s1_f[66]), .Z0_t (KeyReg_Inst_ff_SDE_66_MUX_inst_X), .Z0_f (new_AGEMA_signal_15479), .Z1_t (new_AGEMA_signal_15480), .Z1_f (new_AGEMA_signal_15481) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_66_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_66_MUX_inst_X), .B0_f (new_AGEMA_signal_15479), .B1_t (new_AGEMA_signal_15480), .B1_f (new_AGEMA_signal_15481), .Z0_t (KeyReg_Inst_ff_SDE_66_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16358), .Z1_t (new_AGEMA_signal_16359), .Z1_f (new_AGEMA_signal_16360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_66_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_66_MUX_inst_Y), .A0_f (new_AGEMA_signal_16358), .A1_t (new_AGEMA_signal_16359), .A1_f (new_AGEMA_signal_16360), .B0_t (KeyExpansionOutput[66]), .B0_f (new_AGEMA_signal_14990), .B1_t (new_AGEMA_signal_14991), .B1_f (new_AGEMA_signal_14992), .Z0_t (RoundKey[66]), .Z0_f (new_AGEMA_signal_5873), .Z1_t (new_AGEMA_signal_5874), .Z1_f (new_AGEMA_signal_5875) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_67_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[67]), .A0_f (new_AGEMA_signal_14987), .A1_t (new_AGEMA_signal_14988), .A1_f (new_AGEMA_signal_14989), .B0_t (key_s0_t[67]), .B0_f (key_s0_f[67]), .B1_t (key_s1_t[67]), .B1_f (key_s1_f[67]), .Z0_t (KeyReg_Inst_ff_SDE_67_MUX_inst_X), .Z0_f (new_AGEMA_signal_15485), .Z1_t (new_AGEMA_signal_15486), .Z1_f (new_AGEMA_signal_15487) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_67_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_67_MUX_inst_X), .B0_f (new_AGEMA_signal_15485), .B1_t (new_AGEMA_signal_15486), .B1_f (new_AGEMA_signal_15487), .Z0_t (KeyReg_Inst_ff_SDE_67_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16361), .Z1_t (new_AGEMA_signal_16362), .Z1_f (new_AGEMA_signal_16363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_67_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_67_MUX_inst_Y), .A0_f (new_AGEMA_signal_16361), .A1_t (new_AGEMA_signal_16362), .A1_f (new_AGEMA_signal_16363), .B0_t (KeyExpansionOutput[67]), .B0_f (new_AGEMA_signal_14987), .B1_t (new_AGEMA_signal_14988), .B1_f (new_AGEMA_signal_14989), .Z0_t (RoundKey[67]), .Z0_f (new_AGEMA_signal_5882), .Z1_t (new_AGEMA_signal_5883), .Z1_f (new_AGEMA_signal_5884) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_68_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[68]), .A0_f (new_AGEMA_signal_14984), .A1_t (new_AGEMA_signal_14985), .A1_f (new_AGEMA_signal_14986), .B0_t (key_s0_t[68]), .B0_f (key_s0_f[68]), .B1_t (key_s1_t[68]), .B1_f (key_s1_f[68]), .Z0_t (KeyReg_Inst_ff_SDE_68_MUX_inst_X), .Z0_f (new_AGEMA_signal_15491), .Z1_t (new_AGEMA_signal_15492), .Z1_f (new_AGEMA_signal_15493) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_68_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_68_MUX_inst_X), .B0_f (new_AGEMA_signal_15491), .B1_t (new_AGEMA_signal_15492), .B1_f (new_AGEMA_signal_15493), .Z0_t (KeyReg_Inst_ff_SDE_68_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16364), .Z1_t (new_AGEMA_signal_16365), .Z1_f (new_AGEMA_signal_16366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_68_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_68_MUX_inst_Y), .A0_f (new_AGEMA_signal_16364), .A1_t (new_AGEMA_signal_16365), .A1_f (new_AGEMA_signal_16366), .B0_t (KeyExpansionOutput[68]), .B0_f (new_AGEMA_signal_14984), .B1_t (new_AGEMA_signal_14985), .B1_f (new_AGEMA_signal_14986), .Z0_t (RoundKey[68]), .Z0_f (new_AGEMA_signal_5891), .Z1_t (new_AGEMA_signal_5892), .Z1_f (new_AGEMA_signal_5893) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_69_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[69]), .A0_f (new_AGEMA_signal_14981), .A1_t (new_AGEMA_signal_14982), .A1_f (new_AGEMA_signal_14983), .B0_t (key_s0_t[69]), .B0_f (key_s0_f[69]), .B1_t (key_s1_t[69]), .B1_f (key_s1_f[69]), .Z0_t (KeyReg_Inst_ff_SDE_69_MUX_inst_X), .Z0_f (new_AGEMA_signal_15497), .Z1_t (new_AGEMA_signal_15498), .Z1_f (new_AGEMA_signal_15499) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_69_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_69_MUX_inst_X), .B0_f (new_AGEMA_signal_15497), .B1_t (new_AGEMA_signal_15498), .B1_f (new_AGEMA_signal_15499), .Z0_t (KeyReg_Inst_ff_SDE_69_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16367), .Z1_t (new_AGEMA_signal_16368), .Z1_f (new_AGEMA_signal_16369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_69_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_69_MUX_inst_Y), .A0_f (new_AGEMA_signal_16367), .A1_t (new_AGEMA_signal_16368), .A1_f (new_AGEMA_signal_16369), .B0_t (KeyExpansionOutput[69]), .B0_f (new_AGEMA_signal_14981), .B1_t (new_AGEMA_signal_14982), .B1_f (new_AGEMA_signal_14983), .Z0_t (RoundKey[69]), .Z0_f (new_AGEMA_signal_5900), .Z1_t (new_AGEMA_signal_5901), .Z1_f (new_AGEMA_signal_5902) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_70_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[70]), .A0_f (new_AGEMA_signal_14978), .A1_t (new_AGEMA_signal_14979), .A1_f (new_AGEMA_signal_14980), .B0_t (key_s0_t[70]), .B0_f (key_s0_f[70]), .B1_t (key_s1_t[70]), .B1_f (key_s1_f[70]), .Z0_t (KeyReg_Inst_ff_SDE_70_MUX_inst_X), .Z0_f (new_AGEMA_signal_15503), .Z1_t (new_AGEMA_signal_15504), .Z1_f (new_AGEMA_signal_15505) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_70_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_70_MUX_inst_X), .B0_f (new_AGEMA_signal_15503), .B1_t (new_AGEMA_signal_15504), .B1_f (new_AGEMA_signal_15505), .Z0_t (KeyReg_Inst_ff_SDE_70_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16370), .Z1_t (new_AGEMA_signal_16371), .Z1_f (new_AGEMA_signal_16372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_70_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_70_MUX_inst_Y), .A0_f (new_AGEMA_signal_16370), .A1_t (new_AGEMA_signal_16371), .A1_f (new_AGEMA_signal_16372), .B0_t (KeyExpansionOutput[70]), .B0_f (new_AGEMA_signal_14978), .B1_t (new_AGEMA_signal_14979), .B1_f (new_AGEMA_signal_14980), .Z0_t (RoundKey[70]), .Z0_f (new_AGEMA_signal_5918), .Z1_t (new_AGEMA_signal_5919), .Z1_f (new_AGEMA_signal_5920) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_71_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[71]), .A0_f (new_AGEMA_signal_14975), .A1_t (new_AGEMA_signal_14976), .A1_f (new_AGEMA_signal_14977), .B0_t (key_s0_t[71]), .B0_f (key_s0_f[71]), .B1_t (key_s1_t[71]), .B1_f (key_s1_f[71]), .Z0_t (KeyReg_Inst_ff_SDE_71_MUX_inst_X), .Z0_f (new_AGEMA_signal_15509), .Z1_t (new_AGEMA_signal_15510), .Z1_f (new_AGEMA_signal_15511) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_71_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_71_MUX_inst_X), .B0_f (new_AGEMA_signal_15509), .B1_t (new_AGEMA_signal_15510), .B1_f (new_AGEMA_signal_15511), .Z0_t (KeyReg_Inst_ff_SDE_71_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16373), .Z1_t (new_AGEMA_signal_16374), .Z1_f (new_AGEMA_signal_16375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_71_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_71_MUX_inst_Y), .A0_f (new_AGEMA_signal_16373), .A1_t (new_AGEMA_signal_16374), .A1_f (new_AGEMA_signal_16375), .B0_t (KeyExpansionOutput[71]), .B0_f (new_AGEMA_signal_14975), .B1_t (new_AGEMA_signal_14976), .B1_f (new_AGEMA_signal_14977), .Z0_t (RoundKey[71]), .Z0_f (new_AGEMA_signal_5927), .Z1_t (new_AGEMA_signal_5928), .Z1_f (new_AGEMA_signal_5929) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_72_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[72]), .A0_f (new_AGEMA_signal_13994), .A1_t (new_AGEMA_signal_13995), .A1_f (new_AGEMA_signal_13996), .B0_t (key_s0_t[72]), .B0_f (key_s0_f[72]), .B1_t (key_s1_t[72]), .B1_f (key_s1_f[72]), .Z0_t (KeyReg_Inst_ff_SDE_72_MUX_inst_X), .Z0_f (new_AGEMA_signal_14819), .Z1_t (new_AGEMA_signal_14820), .Z1_f (new_AGEMA_signal_14821) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_72_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_72_MUX_inst_X), .B0_f (new_AGEMA_signal_14819), .B1_t (new_AGEMA_signal_14820), .B1_f (new_AGEMA_signal_14821), .Z0_t (KeyReg_Inst_ff_SDE_72_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15512), .Z1_t (new_AGEMA_signal_15513), .Z1_f (new_AGEMA_signal_15514) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_72_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_72_MUX_inst_Y), .A0_f (new_AGEMA_signal_15512), .A1_t (new_AGEMA_signal_15513), .A1_f (new_AGEMA_signal_15514), .B0_t (KeyExpansionOutput[72]), .B0_f (new_AGEMA_signal_13994), .B1_t (new_AGEMA_signal_13995), .B1_f (new_AGEMA_signal_13996), .Z0_t (RoundKey[72]), .Z0_f (new_AGEMA_signal_5936), .Z1_t (new_AGEMA_signal_5937), .Z1_f (new_AGEMA_signal_5938) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_73_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[73]), .A0_f (new_AGEMA_signal_14969), .A1_t (new_AGEMA_signal_14970), .A1_f (new_AGEMA_signal_14971), .B0_t (key_s0_t[73]), .B0_f (key_s0_f[73]), .B1_t (key_s1_t[73]), .B1_f (key_s1_f[73]), .Z0_t (KeyReg_Inst_ff_SDE_73_MUX_inst_X), .Z0_f (new_AGEMA_signal_15518), .Z1_t (new_AGEMA_signal_15519), .Z1_f (new_AGEMA_signal_15520) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_73_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_73_MUX_inst_X), .B0_f (new_AGEMA_signal_15518), .B1_t (new_AGEMA_signal_15519), .B1_f (new_AGEMA_signal_15520), .Z0_t (KeyReg_Inst_ff_SDE_73_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16376), .Z1_t (new_AGEMA_signal_16377), .Z1_f (new_AGEMA_signal_16378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_73_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_73_MUX_inst_Y), .A0_f (new_AGEMA_signal_16376), .A1_t (new_AGEMA_signal_16377), .A1_f (new_AGEMA_signal_16378), .B0_t (KeyExpansionOutput[73]), .B0_f (new_AGEMA_signal_14969), .B1_t (new_AGEMA_signal_14970), .B1_f (new_AGEMA_signal_14971), .Z0_t (RoundKey[73]), .Z0_f (new_AGEMA_signal_5945), .Z1_t (new_AGEMA_signal_5946), .Z1_f (new_AGEMA_signal_5947) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_74_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[74]), .A0_f (new_AGEMA_signal_15059), .A1_t (new_AGEMA_signal_15060), .A1_f (new_AGEMA_signal_15061), .B0_t (key_s0_t[74]), .B0_f (key_s0_f[74]), .B1_t (key_s1_t[74]), .B1_f (key_s1_f[74]), .Z0_t (KeyReg_Inst_ff_SDE_74_MUX_inst_X), .Z0_f (new_AGEMA_signal_15524), .Z1_t (new_AGEMA_signal_15525), .Z1_f (new_AGEMA_signal_15526) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_74_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_74_MUX_inst_X), .B0_f (new_AGEMA_signal_15524), .B1_t (new_AGEMA_signal_15525), .B1_f (new_AGEMA_signal_15526), .Z0_t (KeyReg_Inst_ff_SDE_74_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16379), .Z1_t (new_AGEMA_signal_16380), .Z1_f (new_AGEMA_signal_16381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_74_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_74_MUX_inst_Y), .A0_f (new_AGEMA_signal_16379), .A1_t (new_AGEMA_signal_16380), .A1_f (new_AGEMA_signal_16381), .B0_t (KeyExpansionOutput[74]), .B0_f (new_AGEMA_signal_15059), .B1_t (new_AGEMA_signal_15060), .B1_f (new_AGEMA_signal_15061), .Z0_t (RoundKey[74]), .Z0_f (new_AGEMA_signal_5954), .Z1_t (new_AGEMA_signal_5955), .Z1_f (new_AGEMA_signal_5956) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_75_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[75]), .A0_f (new_AGEMA_signal_15056), .A1_t (new_AGEMA_signal_15057), .A1_f (new_AGEMA_signal_15058), .B0_t (key_s0_t[75]), .B0_f (key_s0_f[75]), .B1_t (key_s1_t[75]), .B1_f (key_s1_f[75]), .Z0_t (KeyReg_Inst_ff_SDE_75_MUX_inst_X), .Z0_f (new_AGEMA_signal_15530), .Z1_t (new_AGEMA_signal_15531), .Z1_f (new_AGEMA_signal_15532) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_75_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_75_MUX_inst_X), .B0_f (new_AGEMA_signal_15530), .B1_t (new_AGEMA_signal_15531), .B1_f (new_AGEMA_signal_15532), .Z0_t (KeyReg_Inst_ff_SDE_75_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16382), .Z1_t (new_AGEMA_signal_16383), .Z1_f (new_AGEMA_signal_16384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_75_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_75_MUX_inst_Y), .A0_f (new_AGEMA_signal_16382), .A1_t (new_AGEMA_signal_16383), .A1_f (new_AGEMA_signal_16384), .B0_t (KeyExpansionOutput[75]), .B0_f (new_AGEMA_signal_15056), .B1_t (new_AGEMA_signal_15057), .B1_f (new_AGEMA_signal_15058), .Z0_t (RoundKey[75]), .Z0_f (new_AGEMA_signal_5963), .Z1_t (new_AGEMA_signal_5964), .Z1_f (new_AGEMA_signal_5965) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_76_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[76]), .A0_f (new_AGEMA_signal_15032), .A1_t (new_AGEMA_signal_15033), .A1_f (new_AGEMA_signal_15034), .B0_t (key_s0_t[76]), .B0_f (key_s0_f[76]), .B1_t (key_s1_t[76]), .B1_f (key_s1_f[76]), .Z0_t (KeyReg_Inst_ff_SDE_76_MUX_inst_X), .Z0_f (new_AGEMA_signal_15536), .Z1_t (new_AGEMA_signal_15537), .Z1_f (new_AGEMA_signal_15538) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_76_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_76_MUX_inst_X), .B0_f (new_AGEMA_signal_15536), .B1_t (new_AGEMA_signal_15537), .B1_f (new_AGEMA_signal_15538), .Z0_t (KeyReg_Inst_ff_SDE_76_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16385), .Z1_t (new_AGEMA_signal_16386), .Z1_f (new_AGEMA_signal_16387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_76_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_76_MUX_inst_Y), .A0_f (new_AGEMA_signal_16385), .A1_t (new_AGEMA_signal_16386), .A1_f (new_AGEMA_signal_16387), .B0_t (KeyExpansionOutput[76]), .B0_f (new_AGEMA_signal_15032), .B1_t (new_AGEMA_signal_15033), .B1_f (new_AGEMA_signal_15034), .Z0_t (RoundKey[76]), .Z0_f (new_AGEMA_signal_5972), .Z1_t (new_AGEMA_signal_5973), .Z1_f (new_AGEMA_signal_5974) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_77_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[77]), .A0_f (new_AGEMA_signal_15029), .A1_t (new_AGEMA_signal_15030), .A1_f (new_AGEMA_signal_15031), .B0_t (key_s0_t[77]), .B0_f (key_s0_f[77]), .B1_t (key_s1_t[77]), .B1_f (key_s1_f[77]), .Z0_t (KeyReg_Inst_ff_SDE_77_MUX_inst_X), .Z0_f (new_AGEMA_signal_15542), .Z1_t (new_AGEMA_signal_15543), .Z1_f (new_AGEMA_signal_15544) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_77_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_77_MUX_inst_X), .B0_f (new_AGEMA_signal_15542), .B1_t (new_AGEMA_signal_15543), .B1_f (new_AGEMA_signal_15544), .Z0_t (KeyReg_Inst_ff_SDE_77_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16388), .Z1_t (new_AGEMA_signal_16389), .Z1_f (new_AGEMA_signal_16390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_77_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_77_MUX_inst_Y), .A0_f (new_AGEMA_signal_16388), .A1_t (new_AGEMA_signal_16389), .A1_f (new_AGEMA_signal_16390), .B0_t (KeyExpansionOutput[77]), .B0_f (new_AGEMA_signal_15029), .B1_t (new_AGEMA_signal_15030), .B1_f (new_AGEMA_signal_15031), .Z0_t (RoundKey[77]), .Z0_f (new_AGEMA_signal_5981), .Z1_t (new_AGEMA_signal_5982), .Z1_f (new_AGEMA_signal_5983) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_78_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[78]), .A0_f (new_AGEMA_signal_15026), .A1_t (new_AGEMA_signal_15027), .A1_f (new_AGEMA_signal_15028), .B0_t (key_s0_t[78]), .B0_f (key_s0_f[78]), .B1_t (key_s1_t[78]), .B1_f (key_s1_f[78]), .Z0_t (KeyReg_Inst_ff_SDE_78_MUX_inst_X), .Z0_f (new_AGEMA_signal_15548), .Z1_t (new_AGEMA_signal_15549), .Z1_f (new_AGEMA_signal_15550) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_78_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_78_MUX_inst_X), .B0_f (new_AGEMA_signal_15548), .B1_t (new_AGEMA_signal_15549), .B1_f (new_AGEMA_signal_15550), .Z0_t (KeyReg_Inst_ff_SDE_78_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16391), .Z1_t (new_AGEMA_signal_16392), .Z1_f (new_AGEMA_signal_16393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_78_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_78_MUX_inst_Y), .A0_f (new_AGEMA_signal_16391), .A1_t (new_AGEMA_signal_16392), .A1_f (new_AGEMA_signal_16393), .B0_t (KeyExpansionOutput[78]), .B0_f (new_AGEMA_signal_15026), .B1_t (new_AGEMA_signal_15027), .B1_f (new_AGEMA_signal_15028), .Z0_t (RoundKey[78]), .Z0_f (new_AGEMA_signal_5990), .Z1_t (new_AGEMA_signal_5991), .Z1_f (new_AGEMA_signal_5992) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_79_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[79]), .A0_f (new_AGEMA_signal_15023), .A1_t (new_AGEMA_signal_15024), .A1_f (new_AGEMA_signal_15025), .B0_t (key_s0_t[79]), .B0_f (key_s0_f[79]), .B1_t (key_s1_t[79]), .B1_f (key_s1_f[79]), .Z0_t (KeyReg_Inst_ff_SDE_79_MUX_inst_X), .Z0_f (new_AGEMA_signal_15554), .Z1_t (new_AGEMA_signal_15555), .Z1_f (new_AGEMA_signal_15556) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_79_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_79_MUX_inst_X), .B0_f (new_AGEMA_signal_15554), .B1_t (new_AGEMA_signal_15555), .B1_f (new_AGEMA_signal_15556), .Z0_t (KeyReg_Inst_ff_SDE_79_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16394), .Z1_t (new_AGEMA_signal_16395), .Z1_f (new_AGEMA_signal_16396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_79_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_79_MUX_inst_Y), .A0_f (new_AGEMA_signal_16394), .A1_t (new_AGEMA_signal_16395), .A1_f (new_AGEMA_signal_16396), .B0_t (KeyExpansionOutput[79]), .B0_f (new_AGEMA_signal_15023), .B1_t (new_AGEMA_signal_15024), .B1_f (new_AGEMA_signal_15025), .Z0_t (RoundKey[79]), .Z0_f (new_AGEMA_signal_5999), .Z1_t (new_AGEMA_signal_6000), .Z1_f (new_AGEMA_signal_6001) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_80_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[80]), .A0_f (new_AGEMA_signal_14006), .A1_t (new_AGEMA_signal_14007), .A1_f (new_AGEMA_signal_14008), .B0_t (key_s0_t[80]), .B0_f (key_s0_f[80]), .B1_t (key_s1_t[80]), .B1_f (key_s1_f[80]), .Z0_t (KeyReg_Inst_ff_SDE_80_MUX_inst_X), .Z0_f (new_AGEMA_signal_14825), .Z1_t (new_AGEMA_signal_14826), .Z1_f (new_AGEMA_signal_14827) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_80_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_80_MUX_inst_X), .B0_f (new_AGEMA_signal_14825), .B1_t (new_AGEMA_signal_14826), .B1_f (new_AGEMA_signal_14827), .Z0_t (KeyReg_Inst_ff_SDE_80_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15557), .Z1_t (new_AGEMA_signal_15558), .Z1_f (new_AGEMA_signal_15559) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_80_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_80_MUX_inst_Y), .A0_f (new_AGEMA_signal_15557), .A1_t (new_AGEMA_signal_15558), .A1_f (new_AGEMA_signal_15559), .B0_t (KeyExpansionOutput[80]), .B0_f (new_AGEMA_signal_14006), .B1_t (new_AGEMA_signal_14007), .B1_f (new_AGEMA_signal_14008), .Z0_t (RoundKey[80]), .Z0_f (new_AGEMA_signal_6017), .Z1_t (new_AGEMA_signal_6018), .Z1_f (new_AGEMA_signal_6019) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_81_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[81]), .A0_f (new_AGEMA_signal_15017), .A1_t (new_AGEMA_signal_15018), .A1_f (new_AGEMA_signal_15019), .B0_t (key_s0_t[81]), .B0_f (key_s0_f[81]), .B1_t (key_s1_t[81]), .B1_f (key_s1_f[81]), .Z0_t (KeyReg_Inst_ff_SDE_81_MUX_inst_X), .Z0_f (new_AGEMA_signal_15563), .Z1_t (new_AGEMA_signal_15564), .Z1_f (new_AGEMA_signal_15565) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_81_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_81_MUX_inst_X), .B0_f (new_AGEMA_signal_15563), .B1_t (new_AGEMA_signal_15564), .B1_f (new_AGEMA_signal_15565), .Z0_t (KeyReg_Inst_ff_SDE_81_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16397), .Z1_t (new_AGEMA_signal_16398), .Z1_f (new_AGEMA_signal_16399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_81_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_81_MUX_inst_Y), .A0_f (new_AGEMA_signal_16397), .A1_t (new_AGEMA_signal_16398), .A1_f (new_AGEMA_signal_16399), .B0_t (KeyExpansionOutput[81]), .B0_f (new_AGEMA_signal_15017), .B1_t (new_AGEMA_signal_15018), .B1_f (new_AGEMA_signal_15019), .Z0_t (RoundKey[81]), .Z0_f (new_AGEMA_signal_6026), .Z1_t (new_AGEMA_signal_6027), .Z1_f (new_AGEMA_signal_6028) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_82_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[82]), .A0_f (new_AGEMA_signal_15014), .A1_t (new_AGEMA_signal_15015), .A1_f (new_AGEMA_signal_15016), .B0_t (key_s0_t[82]), .B0_f (key_s0_f[82]), .B1_t (key_s1_t[82]), .B1_f (key_s1_f[82]), .Z0_t (KeyReg_Inst_ff_SDE_82_MUX_inst_X), .Z0_f (new_AGEMA_signal_15569), .Z1_t (new_AGEMA_signal_15570), .Z1_f (new_AGEMA_signal_15571) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_82_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_82_MUX_inst_X), .B0_f (new_AGEMA_signal_15569), .B1_t (new_AGEMA_signal_15570), .B1_f (new_AGEMA_signal_15571), .Z0_t (KeyReg_Inst_ff_SDE_82_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16400), .Z1_t (new_AGEMA_signal_16401), .Z1_f (new_AGEMA_signal_16402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_82_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_82_MUX_inst_Y), .A0_f (new_AGEMA_signal_16400), .A1_t (new_AGEMA_signal_16401), .A1_f (new_AGEMA_signal_16402), .B0_t (KeyExpansionOutput[82]), .B0_f (new_AGEMA_signal_15014), .B1_t (new_AGEMA_signal_15015), .B1_f (new_AGEMA_signal_15016), .Z0_t (RoundKey[82]), .Z0_f (new_AGEMA_signal_6035), .Z1_t (new_AGEMA_signal_6036), .Z1_f (new_AGEMA_signal_6037) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_83_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[83]), .A0_f (new_AGEMA_signal_15011), .A1_t (new_AGEMA_signal_15012), .A1_f (new_AGEMA_signal_15013), .B0_t (key_s0_t[83]), .B0_f (key_s0_f[83]), .B1_t (key_s1_t[83]), .B1_f (key_s1_f[83]), .Z0_t (KeyReg_Inst_ff_SDE_83_MUX_inst_X), .Z0_f (new_AGEMA_signal_15575), .Z1_t (new_AGEMA_signal_15576), .Z1_f (new_AGEMA_signal_15577) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_83_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_83_MUX_inst_X), .B0_f (new_AGEMA_signal_15575), .B1_t (new_AGEMA_signal_15576), .B1_f (new_AGEMA_signal_15577), .Z0_t (KeyReg_Inst_ff_SDE_83_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16403), .Z1_t (new_AGEMA_signal_16404), .Z1_f (new_AGEMA_signal_16405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_83_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_83_MUX_inst_Y), .A0_f (new_AGEMA_signal_16403), .A1_t (new_AGEMA_signal_16404), .A1_f (new_AGEMA_signal_16405), .B0_t (KeyExpansionOutput[83]), .B0_f (new_AGEMA_signal_15011), .B1_t (new_AGEMA_signal_15012), .B1_f (new_AGEMA_signal_15013), .Z0_t (RoundKey[83]), .Z0_f (new_AGEMA_signal_6044), .Z1_t (new_AGEMA_signal_6045), .Z1_f (new_AGEMA_signal_6046) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_84_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[84]), .A0_f (new_AGEMA_signal_15005), .A1_t (new_AGEMA_signal_15006), .A1_f (new_AGEMA_signal_15007), .B0_t (key_s0_t[84]), .B0_f (key_s0_f[84]), .B1_t (key_s1_t[84]), .B1_f (key_s1_f[84]), .Z0_t (KeyReg_Inst_ff_SDE_84_MUX_inst_X), .Z0_f (new_AGEMA_signal_15581), .Z1_t (new_AGEMA_signal_15582), .Z1_f (new_AGEMA_signal_15583) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_84_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_84_MUX_inst_X), .B0_f (new_AGEMA_signal_15581), .B1_t (new_AGEMA_signal_15582), .B1_f (new_AGEMA_signal_15583), .Z0_t (KeyReg_Inst_ff_SDE_84_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16406), .Z1_t (new_AGEMA_signal_16407), .Z1_f (new_AGEMA_signal_16408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_84_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_84_MUX_inst_Y), .A0_f (new_AGEMA_signal_16406), .A1_t (new_AGEMA_signal_16407), .A1_f (new_AGEMA_signal_16408), .B0_t (KeyExpansionOutput[84]), .B0_f (new_AGEMA_signal_15005), .B1_t (new_AGEMA_signal_15006), .B1_f (new_AGEMA_signal_15007), .Z0_t (RoundKey[84]), .Z0_f (new_AGEMA_signal_6053), .Z1_t (new_AGEMA_signal_6054), .Z1_f (new_AGEMA_signal_6055) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_85_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[85]), .A0_f (new_AGEMA_signal_15002), .A1_t (new_AGEMA_signal_15003), .A1_f (new_AGEMA_signal_15004), .B0_t (key_s0_t[85]), .B0_f (key_s0_f[85]), .B1_t (key_s1_t[85]), .B1_f (key_s1_f[85]), .Z0_t (KeyReg_Inst_ff_SDE_85_MUX_inst_X), .Z0_f (new_AGEMA_signal_15587), .Z1_t (new_AGEMA_signal_15588), .Z1_f (new_AGEMA_signal_15589) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_85_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_85_MUX_inst_X), .B0_f (new_AGEMA_signal_15587), .B1_t (new_AGEMA_signal_15588), .B1_f (new_AGEMA_signal_15589), .Z0_t (KeyReg_Inst_ff_SDE_85_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16409), .Z1_t (new_AGEMA_signal_16410), .Z1_f (new_AGEMA_signal_16411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_85_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_85_MUX_inst_Y), .A0_f (new_AGEMA_signal_16409), .A1_t (new_AGEMA_signal_16410), .A1_f (new_AGEMA_signal_16411), .B0_t (KeyExpansionOutput[85]), .B0_f (new_AGEMA_signal_15002), .B1_t (new_AGEMA_signal_15003), .B1_f (new_AGEMA_signal_15004), .Z0_t (RoundKey[85]), .Z0_f (new_AGEMA_signal_6062), .Z1_t (new_AGEMA_signal_6063), .Z1_f (new_AGEMA_signal_6064) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_86_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[86]), .A0_f (new_AGEMA_signal_14999), .A1_t (new_AGEMA_signal_15000), .A1_f (new_AGEMA_signal_15001), .B0_t (key_s0_t[86]), .B0_f (key_s0_f[86]), .B1_t (key_s1_t[86]), .B1_f (key_s1_f[86]), .Z0_t (KeyReg_Inst_ff_SDE_86_MUX_inst_X), .Z0_f (new_AGEMA_signal_15593), .Z1_t (new_AGEMA_signal_15594), .Z1_f (new_AGEMA_signal_15595) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_86_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_86_MUX_inst_X), .B0_f (new_AGEMA_signal_15593), .B1_t (new_AGEMA_signal_15594), .B1_f (new_AGEMA_signal_15595), .Z0_t (KeyReg_Inst_ff_SDE_86_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16412), .Z1_t (new_AGEMA_signal_16413), .Z1_f (new_AGEMA_signal_16414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_86_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_86_MUX_inst_Y), .A0_f (new_AGEMA_signal_16412), .A1_t (new_AGEMA_signal_16413), .A1_f (new_AGEMA_signal_16414), .B0_t (KeyExpansionOutput[86]), .B0_f (new_AGEMA_signal_14999), .B1_t (new_AGEMA_signal_15000), .B1_f (new_AGEMA_signal_15001), .Z0_t (RoundKey[86]), .Z0_f (new_AGEMA_signal_6071), .Z1_t (new_AGEMA_signal_6072), .Z1_f (new_AGEMA_signal_6073) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_87_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[87]), .A0_f (new_AGEMA_signal_14996), .A1_t (new_AGEMA_signal_14997), .A1_f (new_AGEMA_signal_14998), .B0_t (key_s0_t[87]), .B0_f (key_s0_f[87]), .B1_t (key_s1_t[87]), .B1_f (key_s1_f[87]), .Z0_t (KeyReg_Inst_ff_SDE_87_MUX_inst_X), .Z0_f (new_AGEMA_signal_15599), .Z1_t (new_AGEMA_signal_15600), .Z1_f (new_AGEMA_signal_15601) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_87_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_87_MUX_inst_X), .B0_f (new_AGEMA_signal_15599), .B1_t (new_AGEMA_signal_15600), .B1_f (new_AGEMA_signal_15601), .Z0_t (KeyReg_Inst_ff_SDE_87_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16415), .Z1_t (new_AGEMA_signal_16416), .Z1_f (new_AGEMA_signal_16417) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_87_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_87_MUX_inst_Y), .A0_f (new_AGEMA_signal_16415), .A1_t (new_AGEMA_signal_16416), .A1_f (new_AGEMA_signal_16417), .B0_t (KeyExpansionOutput[87]), .B0_f (new_AGEMA_signal_14996), .B1_t (new_AGEMA_signal_14997), .B1_f (new_AGEMA_signal_14998), .Z0_t (RoundKey[87]), .Z0_f (new_AGEMA_signal_6080), .Z1_t (new_AGEMA_signal_6081), .Z1_f (new_AGEMA_signal_6082) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_88_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[88]), .A0_f (new_AGEMA_signal_14993), .A1_t (new_AGEMA_signal_14994), .A1_f (new_AGEMA_signal_14995), .B0_t (key_s0_t[88]), .B0_f (key_s0_f[88]), .B1_t (key_s1_t[88]), .B1_f (key_s1_f[88]), .Z0_t (KeyReg_Inst_ff_SDE_88_MUX_inst_X), .Z0_f (new_AGEMA_signal_15605), .Z1_t (new_AGEMA_signal_15606), .Z1_f (new_AGEMA_signal_15607) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_88_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_88_MUX_inst_X), .B0_f (new_AGEMA_signal_15605), .B1_t (new_AGEMA_signal_15606), .B1_f (new_AGEMA_signal_15607), .Z0_t (KeyReg_Inst_ff_SDE_88_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16418), .Z1_t (new_AGEMA_signal_16419), .Z1_f (new_AGEMA_signal_16420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_88_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_88_MUX_inst_Y), .A0_f (new_AGEMA_signal_16418), .A1_t (new_AGEMA_signal_16419), .A1_f (new_AGEMA_signal_16420), .B0_t (KeyExpansionOutput[88]), .B0_f (new_AGEMA_signal_14993), .B1_t (new_AGEMA_signal_14994), .B1_f (new_AGEMA_signal_14995), .Z0_t (RoundKey[88]), .Z0_f (new_AGEMA_signal_6089), .Z1_t (new_AGEMA_signal_6090), .Z1_f (new_AGEMA_signal_6091) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_89_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[89]), .A0_f (new_AGEMA_signal_15758), .A1_t (new_AGEMA_signal_15759), .A1_f (new_AGEMA_signal_15760), .B0_t (key_s0_t[89]), .B0_f (key_s0_f[89]), .B1_t (key_s1_t[89]), .B1_f (key_s1_f[89]), .Z0_t (KeyReg_Inst_ff_SDE_89_MUX_inst_X), .Z0_f (new_AGEMA_signal_16424), .Z1_t (new_AGEMA_signal_16425), .Z1_f (new_AGEMA_signal_16426) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_89_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_89_MUX_inst_X), .B0_f (new_AGEMA_signal_16424), .B1_t (new_AGEMA_signal_16425), .B1_f (new_AGEMA_signal_16426), .Z0_t (KeyReg_Inst_ff_SDE_89_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17204), .Z1_t (new_AGEMA_signal_17205), .Z1_f (new_AGEMA_signal_17206) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_89_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_89_MUX_inst_Y), .A0_f (new_AGEMA_signal_17204), .A1_t (new_AGEMA_signal_17205), .A1_f (new_AGEMA_signal_17206), .B0_t (KeyExpansionOutput[89]), .B0_f (new_AGEMA_signal_15758), .B1_t (new_AGEMA_signal_15759), .B1_f (new_AGEMA_signal_15760), .Z0_t (RoundKey[89]), .Z0_f (new_AGEMA_signal_6098), .Z1_t (new_AGEMA_signal_6099), .Z1_f (new_AGEMA_signal_6100) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_90_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[90]), .A0_f (new_AGEMA_signal_15755), .A1_t (new_AGEMA_signal_15756), .A1_f (new_AGEMA_signal_15757), .B0_t (key_s0_t[90]), .B0_f (key_s0_f[90]), .B1_t (key_s1_t[90]), .B1_f (key_s1_f[90]), .Z0_t (KeyReg_Inst_ff_SDE_90_MUX_inst_X), .Z0_f (new_AGEMA_signal_16430), .Z1_t (new_AGEMA_signal_16431), .Z1_f (new_AGEMA_signal_16432) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_90_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_90_MUX_inst_X), .B0_f (new_AGEMA_signal_16430), .B1_t (new_AGEMA_signal_16431), .B1_f (new_AGEMA_signal_16432), .Z0_t (KeyReg_Inst_ff_SDE_90_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17207), .Z1_t (new_AGEMA_signal_17208), .Z1_f (new_AGEMA_signal_17209) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_90_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_90_MUX_inst_Y), .A0_f (new_AGEMA_signal_17207), .A1_t (new_AGEMA_signal_17208), .A1_f (new_AGEMA_signal_17209), .B0_t (KeyExpansionOutput[90]), .B0_f (new_AGEMA_signal_15755), .B1_t (new_AGEMA_signal_15756), .B1_f (new_AGEMA_signal_15757), .Z0_t (RoundKey[90]), .Z0_f (new_AGEMA_signal_6116), .Z1_t (new_AGEMA_signal_6117), .Z1_f (new_AGEMA_signal_6118) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_91_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[91]), .A0_f (new_AGEMA_signal_15752), .A1_t (new_AGEMA_signal_15753), .A1_f (new_AGEMA_signal_15754), .B0_t (key_s0_t[91]), .B0_f (key_s0_f[91]), .B1_t (key_s1_t[91]), .B1_f (key_s1_f[91]), .Z0_t (KeyReg_Inst_ff_SDE_91_MUX_inst_X), .Z0_f (new_AGEMA_signal_16436), .Z1_t (new_AGEMA_signal_16437), .Z1_f (new_AGEMA_signal_16438) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_91_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_91_MUX_inst_X), .B0_f (new_AGEMA_signal_16436), .B1_t (new_AGEMA_signal_16437), .B1_f (new_AGEMA_signal_16438), .Z0_t (KeyReg_Inst_ff_SDE_91_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17210), .Z1_t (new_AGEMA_signal_17211), .Z1_f (new_AGEMA_signal_17212) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_91_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_91_MUX_inst_Y), .A0_f (new_AGEMA_signal_17210), .A1_t (new_AGEMA_signal_17211), .A1_f (new_AGEMA_signal_17212), .B0_t (KeyExpansionOutput[91]), .B0_f (new_AGEMA_signal_15752), .B1_t (new_AGEMA_signal_15753), .B1_f (new_AGEMA_signal_15754), .Z0_t (RoundKey[91]), .Z0_f (new_AGEMA_signal_6125), .Z1_t (new_AGEMA_signal_6126), .Z1_f (new_AGEMA_signal_6127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_92_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[92]), .A0_f (new_AGEMA_signal_15749), .A1_t (new_AGEMA_signal_15750), .A1_f (new_AGEMA_signal_15751), .B0_t (key_s0_t[92]), .B0_f (key_s0_f[92]), .B1_t (key_s1_t[92]), .B1_f (key_s1_f[92]), .Z0_t (KeyReg_Inst_ff_SDE_92_MUX_inst_X), .Z0_f (new_AGEMA_signal_16442), .Z1_t (new_AGEMA_signal_16443), .Z1_f (new_AGEMA_signal_16444) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_92_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_92_MUX_inst_X), .B0_f (new_AGEMA_signal_16442), .B1_t (new_AGEMA_signal_16443), .B1_f (new_AGEMA_signal_16444), .Z0_t (KeyReg_Inst_ff_SDE_92_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17213), .Z1_t (new_AGEMA_signal_17214), .Z1_f (new_AGEMA_signal_17215) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_92_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_92_MUX_inst_Y), .A0_f (new_AGEMA_signal_17213), .A1_t (new_AGEMA_signal_17214), .A1_f (new_AGEMA_signal_17215), .B0_t (KeyExpansionOutput[92]), .B0_f (new_AGEMA_signal_15749), .B1_t (new_AGEMA_signal_15750), .B1_f (new_AGEMA_signal_15751), .Z0_t (RoundKey[92]), .Z0_f (new_AGEMA_signal_6134), .Z1_t (new_AGEMA_signal_6135), .Z1_f (new_AGEMA_signal_6136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_93_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[93]), .A0_f (new_AGEMA_signal_15746), .A1_t (new_AGEMA_signal_15747), .A1_f (new_AGEMA_signal_15748), .B0_t (key_s0_t[93]), .B0_f (key_s0_f[93]), .B1_t (key_s1_t[93]), .B1_f (key_s1_f[93]), .Z0_t (KeyReg_Inst_ff_SDE_93_MUX_inst_X), .Z0_f (new_AGEMA_signal_16448), .Z1_t (new_AGEMA_signal_16449), .Z1_f (new_AGEMA_signal_16450) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_93_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_93_MUX_inst_X), .B0_f (new_AGEMA_signal_16448), .B1_t (new_AGEMA_signal_16449), .B1_f (new_AGEMA_signal_16450), .Z0_t (KeyReg_Inst_ff_SDE_93_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17216), .Z1_t (new_AGEMA_signal_17217), .Z1_f (new_AGEMA_signal_17218) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_93_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_93_MUX_inst_Y), .A0_f (new_AGEMA_signal_17216), .A1_t (new_AGEMA_signal_17217), .A1_f (new_AGEMA_signal_17218), .B0_t (KeyExpansionOutput[93]), .B0_f (new_AGEMA_signal_15746), .B1_t (new_AGEMA_signal_15747), .B1_f (new_AGEMA_signal_15748), .Z0_t (RoundKey[93]), .Z0_f (new_AGEMA_signal_6143), .Z1_t (new_AGEMA_signal_6144), .Z1_f (new_AGEMA_signal_6145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_94_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[94]), .A0_f (new_AGEMA_signal_15740), .A1_t (new_AGEMA_signal_15741), .A1_f (new_AGEMA_signal_15742), .B0_t (key_s0_t[94]), .B0_f (key_s0_f[94]), .B1_t (key_s1_t[94]), .B1_f (key_s1_f[94]), .Z0_t (KeyReg_Inst_ff_SDE_94_MUX_inst_X), .Z0_f (new_AGEMA_signal_16454), .Z1_t (new_AGEMA_signal_16455), .Z1_f (new_AGEMA_signal_16456) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_94_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_94_MUX_inst_X), .B0_f (new_AGEMA_signal_16454), .B1_t (new_AGEMA_signal_16455), .B1_f (new_AGEMA_signal_16456), .Z0_t (KeyReg_Inst_ff_SDE_94_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17219), .Z1_t (new_AGEMA_signal_17220), .Z1_f (new_AGEMA_signal_17221) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_94_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_94_MUX_inst_Y), .A0_f (new_AGEMA_signal_17219), .A1_t (new_AGEMA_signal_17220), .A1_f (new_AGEMA_signal_17221), .B0_t (KeyExpansionOutput[94]), .B0_f (new_AGEMA_signal_15740), .B1_t (new_AGEMA_signal_15741), .B1_f (new_AGEMA_signal_15742), .Z0_t (RoundKey[94]), .Z0_f (new_AGEMA_signal_6152), .Z1_t (new_AGEMA_signal_6153), .Z1_f (new_AGEMA_signal_6154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_95_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[95]), .A0_f (new_AGEMA_signal_15737), .A1_t (new_AGEMA_signal_15738), .A1_f (new_AGEMA_signal_15739), .B0_t (key_s0_t[95]), .B0_f (key_s0_f[95]), .B1_t (key_s1_t[95]), .B1_f (key_s1_f[95]), .Z0_t (KeyReg_Inst_ff_SDE_95_MUX_inst_X), .Z0_f (new_AGEMA_signal_16460), .Z1_t (new_AGEMA_signal_16461), .Z1_f (new_AGEMA_signal_16462) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_95_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_95_MUX_inst_X), .B0_f (new_AGEMA_signal_16460), .B1_t (new_AGEMA_signal_16461), .B1_f (new_AGEMA_signal_16462), .Z0_t (KeyReg_Inst_ff_SDE_95_MUX_inst_Y), .Z0_f (new_AGEMA_signal_17222), .Z1_t (new_AGEMA_signal_17223), .Z1_f (new_AGEMA_signal_17224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_95_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_95_MUX_inst_Y), .A0_f (new_AGEMA_signal_17222), .A1_t (new_AGEMA_signal_17223), .A1_f (new_AGEMA_signal_17224), .B0_t (KeyExpansionOutput[95]), .B0_f (new_AGEMA_signal_15737), .B1_t (new_AGEMA_signal_15738), .B1_f (new_AGEMA_signal_15739), .Z0_t (RoundKey[95]), .Z0_f (new_AGEMA_signal_6161), .Z1_t (new_AGEMA_signal_6162), .Z1_f (new_AGEMA_signal_6163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_96_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[96]), .A0_f (new_AGEMA_signal_13502), .A1_t (new_AGEMA_signal_13503), .A1_f (new_AGEMA_signal_13504), .B0_t (key_s0_t[96]), .B0_f (key_s0_f[96]), .B1_t (key_s1_t[96]), .B1_f (key_s1_f[96]), .Z0_t (KeyReg_Inst_ff_SDE_96_MUX_inst_X), .Z0_f (new_AGEMA_signal_13979), .Z1_t (new_AGEMA_signal_13980), .Z1_f (new_AGEMA_signal_13981) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_96_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_96_MUX_inst_X), .B0_f (new_AGEMA_signal_13979), .B1_t (new_AGEMA_signal_13980), .B1_f (new_AGEMA_signal_13981), .Z0_t (KeyReg_Inst_ff_SDE_96_MUX_inst_Y), .Z0_f (new_AGEMA_signal_14828), .Z1_t (new_AGEMA_signal_14829), .Z1_f (new_AGEMA_signal_14830) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_96_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_96_MUX_inst_Y), .A0_f (new_AGEMA_signal_14828), .A1_t (new_AGEMA_signal_14829), .A1_f (new_AGEMA_signal_14830), .B0_t (KeyExpansionOutput[96]), .B0_f (new_AGEMA_signal_13502), .B1_t (new_AGEMA_signal_13503), .B1_f (new_AGEMA_signal_13504), .Z0_t (RoundKey[96]), .Z0_f (new_AGEMA_signal_6170), .Z1_t (new_AGEMA_signal_6171), .Z1_f (new_AGEMA_signal_6172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_97_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[97]), .A0_f (new_AGEMA_signal_14003), .A1_t (new_AGEMA_signal_14004), .A1_f (new_AGEMA_signal_14005), .B0_t (key_s0_t[97]), .B0_f (key_s0_f[97]), .B1_t (key_s1_t[97]), .B1_f (key_s1_f[97]), .Z0_t (KeyReg_Inst_ff_SDE_97_MUX_inst_X), .Z0_f (new_AGEMA_signal_14834), .Z1_t (new_AGEMA_signal_14835), .Z1_f (new_AGEMA_signal_14836) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_97_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_97_MUX_inst_X), .B0_f (new_AGEMA_signal_14834), .B1_t (new_AGEMA_signal_14835), .B1_f (new_AGEMA_signal_14836), .Z0_t (KeyReg_Inst_ff_SDE_97_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15608), .Z1_t (new_AGEMA_signal_15609), .Z1_f (new_AGEMA_signal_15610) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_97_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_97_MUX_inst_Y), .A0_f (new_AGEMA_signal_15608), .A1_t (new_AGEMA_signal_15609), .A1_f (new_AGEMA_signal_15610), .B0_t (KeyExpansionOutput[97]), .B0_f (new_AGEMA_signal_14003), .B1_t (new_AGEMA_signal_14004), .B1_f (new_AGEMA_signal_14005), .Z0_t (RoundKey[97]), .Z0_f (new_AGEMA_signal_6179), .Z1_t (new_AGEMA_signal_6180), .Z1_f (new_AGEMA_signal_6181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_98_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[98]), .A0_f (new_AGEMA_signal_14000), .A1_t (new_AGEMA_signal_14001), .A1_f (new_AGEMA_signal_14002), .B0_t (key_s0_t[98]), .B0_f (key_s0_f[98]), .B1_t (key_s1_t[98]), .B1_f (key_s1_f[98]), .Z0_t (KeyReg_Inst_ff_SDE_98_MUX_inst_X), .Z0_f (new_AGEMA_signal_14840), .Z1_t (new_AGEMA_signal_14841), .Z1_f (new_AGEMA_signal_14842) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_98_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_98_MUX_inst_X), .B0_f (new_AGEMA_signal_14840), .B1_t (new_AGEMA_signal_14841), .B1_f (new_AGEMA_signal_14842), .Z0_t (KeyReg_Inst_ff_SDE_98_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15611), .Z1_t (new_AGEMA_signal_15612), .Z1_f (new_AGEMA_signal_15613) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_98_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_98_MUX_inst_Y), .A0_f (new_AGEMA_signal_15611), .A1_t (new_AGEMA_signal_15612), .A1_f (new_AGEMA_signal_15613), .B0_t (KeyExpansionOutput[98]), .B0_f (new_AGEMA_signal_14000), .B1_t (new_AGEMA_signal_14001), .B1_f (new_AGEMA_signal_14002), .Z0_t (RoundKey[98]), .Z0_f (new_AGEMA_signal_6188), .Z1_t (new_AGEMA_signal_6189), .Z1_f (new_AGEMA_signal_6190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_99_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[99]), .A0_f (new_AGEMA_signal_13997), .A1_t (new_AGEMA_signal_13998), .A1_f (new_AGEMA_signal_13999), .B0_t (key_s0_t[99]), .B0_f (key_s0_f[99]), .B1_t (key_s1_t[99]), .B1_f (key_s1_f[99]), .Z0_t (KeyReg_Inst_ff_SDE_99_MUX_inst_X), .Z0_f (new_AGEMA_signal_14846), .Z1_t (new_AGEMA_signal_14847), .Z1_f (new_AGEMA_signal_14848) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_99_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_99_MUX_inst_X), .B0_f (new_AGEMA_signal_14846), .B1_t (new_AGEMA_signal_14847), .B1_f (new_AGEMA_signal_14848), .Z0_t (KeyReg_Inst_ff_SDE_99_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15614), .Z1_t (new_AGEMA_signal_15615), .Z1_f (new_AGEMA_signal_15616) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_99_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_99_MUX_inst_Y), .A0_f (new_AGEMA_signal_15614), .A1_t (new_AGEMA_signal_15615), .A1_f (new_AGEMA_signal_15616), .B0_t (KeyExpansionOutput[99]), .B0_f (new_AGEMA_signal_13997), .B1_t (new_AGEMA_signal_13998), .B1_f (new_AGEMA_signal_13999), .Z0_t (RoundKey[99]), .Z0_f (new_AGEMA_signal_6197), .Z1_t (new_AGEMA_signal_6198), .Z1_f (new_AGEMA_signal_6199) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_100_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[100]), .A0_f (new_AGEMA_signal_14063), .A1_t (new_AGEMA_signal_14064), .A1_f (new_AGEMA_signal_14065), .B0_t (key_s0_t[100]), .B0_f (key_s0_f[100]), .B1_t (key_s1_t[100]), .B1_f (key_s1_f[100]), .Z0_t (KeyReg_Inst_ff_SDE_100_MUX_inst_X), .Z0_f (new_AGEMA_signal_14852), .Z1_t (new_AGEMA_signal_14853), .Z1_f (new_AGEMA_signal_14854) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_100_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_100_MUX_inst_X), .B0_f (new_AGEMA_signal_14852), .B1_t (new_AGEMA_signal_14853), .B1_f (new_AGEMA_signal_14854), .Z0_t (KeyReg_Inst_ff_SDE_100_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15617), .Z1_t (new_AGEMA_signal_15618), .Z1_f (new_AGEMA_signal_15619) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_100_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_100_MUX_inst_Y), .A0_f (new_AGEMA_signal_15617), .A1_t (new_AGEMA_signal_15618), .A1_f (new_AGEMA_signal_15619), .B0_t (KeyExpansionOutput[100]), .B0_f (new_AGEMA_signal_14063), .B1_t (new_AGEMA_signal_14064), .B1_f (new_AGEMA_signal_14065), .Z0_t (RoundKey[100]), .Z0_f (new_AGEMA_signal_5072), .Z1_t (new_AGEMA_signal_5073), .Z1_f (new_AGEMA_signal_5074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_101_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[101]), .A0_f (new_AGEMA_signal_14060), .A1_t (new_AGEMA_signal_14061), .A1_f (new_AGEMA_signal_14062), .B0_t (key_s0_t[101]), .B0_f (key_s0_f[101]), .B1_t (key_s1_t[101]), .B1_f (key_s1_f[101]), .Z0_t (KeyReg_Inst_ff_SDE_101_MUX_inst_X), .Z0_f (new_AGEMA_signal_14858), .Z1_t (new_AGEMA_signal_14859), .Z1_f (new_AGEMA_signal_14860) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_101_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_101_MUX_inst_X), .B0_f (new_AGEMA_signal_14858), .B1_t (new_AGEMA_signal_14859), .B1_f (new_AGEMA_signal_14860), .Z0_t (KeyReg_Inst_ff_SDE_101_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15620), .Z1_t (new_AGEMA_signal_15621), .Z1_f (new_AGEMA_signal_15622) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_101_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_101_MUX_inst_Y), .A0_f (new_AGEMA_signal_15620), .A1_t (new_AGEMA_signal_15621), .A1_f (new_AGEMA_signal_15622), .B0_t (KeyExpansionOutput[101]), .B0_f (new_AGEMA_signal_14060), .B1_t (new_AGEMA_signal_14061), .B1_f (new_AGEMA_signal_14062), .Z0_t (RoundKey[101]), .Z0_f (new_AGEMA_signal_5081), .Z1_t (new_AGEMA_signal_5082), .Z1_f (new_AGEMA_signal_5083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_102_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[102]), .A0_f (new_AGEMA_signal_14057), .A1_t (new_AGEMA_signal_14058), .A1_f (new_AGEMA_signal_14059), .B0_t (key_s0_t[102]), .B0_f (key_s0_f[102]), .B1_t (key_s1_t[102]), .B1_f (key_s1_f[102]), .Z0_t (KeyReg_Inst_ff_SDE_102_MUX_inst_X), .Z0_f (new_AGEMA_signal_14864), .Z1_t (new_AGEMA_signal_14865), .Z1_f (new_AGEMA_signal_14866) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_102_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_102_MUX_inst_X), .B0_f (new_AGEMA_signal_14864), .B1_t (new_AGEMA_signal_14865), .B1_f (new_AGEMA_signal_14866), .Z0_t (KeyReg_Inst_ff_SDE_102_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15623), .Z1_t (new_AGEMA_signal_15624), .Z1_f (new_AGEMA_signal_15625) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_102_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_102_MUX_inst_Y), .A0_f (new_AGEMA_signal_15623), .A1_t (new_AGEMA_signal_15624), .A1_f (new_AGEMA_signal_15625), .B0_t (KeyExpansionOutput[102]), .B0_f (new_AGEMA_signal_14057), .B1_t (new_AGEMA_signal_14058), .B1_f (new_AGEMA_signal_14059), .Z0_t (RoundKey[102]), .Z0_f (new_AGEMA_signal_5090), .Z1_t (new_AGEMA_signal_5091), .Z1_f (new_AGEMA_signal_5092) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_103_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[103]), .A0_f (new_AGEMA_signal_14054), .A1_t (new_AGEMA_signal_14055), .A1_f (new_AGEMA_signal_14056), .B0_t (key_s0_t[103]), .B0_f (key_s0_f[103]), .B1_t (key_s1_t[103]), .B1_f (key_s1_f[103]), .Z0_t (KeyReg_Inst_ff_SDE_103_MUX_inst_X), .Z0_f (new_AGEMA_signal_14870), .Z1_t (new_AGEMA_signal_14871), .Z1_f (new_AGEMA_signal_14872) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_103_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_103_MUX_inst_X), .B0_f (new_AGEMA_signal_14870), .B1_t (new_AGEMA_signal_14871), .B1_f (new_AGEMA_signal_14872), .Z0_t (KeyReg_Inst_ff_SDE_103_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15626), .Z1_t (new_AGEMA_signal_15627), .Z1_f (new_AGEMA_signal_15628) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_103_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_103_MUX_inst_Y), .A0_f (new_AGEMA_signal_15626), .A1_t (new_AGEMA_signal_15627), .A1_f (new_AGEMA_signal_15628), .B0_t (KeyExpansionOutput[103]), .B0_f (new_AGEMA_signal_14054), .B1_t (new_AGEMA_signal_14055), .B1_f (new_AGEMA_signal_14056), .Z0_t (RoundKey[103]), .Z0_f (new_AGEMA_signal_5099), .Z1_t (new_AGEMA_signal_5100), .Z1_f (new_AGEMA_signal_5101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_104_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[104]), .A0_f (new_AGEMA_signal_13499), .A1_t (new_AGEMA_signal_13500), .A1_f (new_AGEMA_signal_13501), .B0_t (key_s0_t[104]), .B0_f (key_s0_f[104]), .B1_t (key_s1_t[104]), .B1_f (key_s1_f[104]), .Z0_t (KeyReg_Inst_ff_SDE_104_MUX_inst_X), .Z0_f (new_AGEMA_signal_13985), .Z1_t (new_AGEMA_signal_13986), .Z1_f (new_AGEMA_signal_13987) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_104_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_104_MUX_inst_X), .B0_f (new_AGEMA_signal_13985), .B1_t (new_AGEMA_signal_13986), .B1_f (new_AGEMA_signal_13987), .Z0_t (KeyReg_Inst_ff_SDE_104_MUX_inst_Y), .Z0_f (new_AGEMA_signal_14873), .Z1_t (new_AGEMA_signal_14874), .Z1_f (new_AGEMA_signal_14875) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_104_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_104_MUX_inst_Y), .A0_f (new_AGEMA_signal_14873), .A1_t (new_AGEMA_signal_14874), .A1_f (new_AGEMA_signal_14875), .B0_t (KeyExpansionOutput[104]), .B0_f (new_AGEMA_signal_13499), .B1_t (new_AGEMA_signal_13500), .B1_f (new_AGEMA_signal_13501), .Z0_t (RoundKey[104]), .Z0_f (new_AGEMA_signal_5108), .Z1_t (new_AGEMA_signal_5109), .Z1_f (new_AGEMA_signal_5110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_105_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[105]), .A0_f (new_AGEMA_signal_14051), .A1_t (new_AGEMA_signal_14052), .A1_f (new_AGEMA_signal_14053), .B0_t (key_s0_t[105]), .B0_f (key_s0_f[105]), .B1_t (key_s1_t[105]), .B1_f (key_s1_f[105]), .Z0_t (KeyReg_Inst_ff_SDE_105_MUX_inst_X), .Z0_f (new_AGEMA_signal_14879), .Z1_t (new_AGEMA_signal_14880), .Z1_f (new_AGEMA_signal_14881) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_105_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_105_MUX_inst_X), .B0_f (new_AGEMA_signal_14879), .B1_t (new_AGEMA_signal_14880), .B1_f (new_AGEMA_signal_14881), .Z0_t (KeyReg_Inst_ff_SDE_105_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15629), .Z1_t (new_AGEMA_signal_15630), .Z1_f (new_AGEMA_signal_15631) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_105_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_105_MUX_inst_Y), .A0_f (new_AGEMA_signal_15629), .A1_t (new_AGEMA_signal_15630), .A1_f (new_AGEMA_signal_15631), .B0_t (KeyExpansionOutput[105]), .B0_f (new_AGEMA_signal_14051), .B1_t (new_AGEMA_signal_14052), .B1_f (new_AGEMA_signal_14053), .Z0_t (RoundKey[105]), .Z0_f (new_AGEMA_signal_5117), .Z1_t (new_AGEMA_signal_5118), .Z1_f (new_AGEMA_signal_5119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_106_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[106]), .A0_f (new_AGEMA_signal_14048), .A1_t (new_AGEMA_signal_14049), .A1_f (new_AGEMA_signal_14050), .B0_t (key_s0_t[106]), .B0_f (key_s0_f[106]), .B1_t (key_s1_t[106]), .B1_f (key_s1_f[106]), .Z0_t (KeyReg_Inst_ff_SDE_106_MUX_inst_X), .Z0_f (new_AGEMA_signal_14885), .Z1_t (new_AGEMA_signal_14886), .Z1_f (new_AGEMA_signal_14887) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_106_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_106_MUX_inst_X), .B0_f (new_AGEMA_signal_14885), .B1_t (new_AGEMA_signal_14886), .B1_f (new_AGEMA_signal_14887), .Z0_t (KeyReg_Inst_ff_SDE_106_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15632), .Z1_t (new_AGEMA_signal_15633), .Z1_f (new_AGEMA_signal_15634) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_106_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_106_MUX_inst_Y), .A0_f (new_AGEMA_signal_15632), .A1_t (new_AGEMA_signal_15633), .A1_f (new_AGEMA_signal_15634), .B0_t (KeyExpansionOutput[106]), .B0_f (new_AGEMA_signal_14048), .B1_t (new_AGEMA_signal_14049), .B1_f (new_AGEMA_signal_14050), .Z0_t (RoundKey[106]), .Z0_f (new_AGEMA_signal_5126), .Z1_t (new_AGEMA_signal_5127), .Z1_f (new_AGEMA_signal_5128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_107_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[107]), .A0_f (new_AGEMA_signal_14045), .A1_t (new_AGEMA_signal_14046), .A1_f (new_AGEMA_signal_14047), .B0_t (key_s0_t[107]), .B0_f (key_s0_f[107]), .B1_t (key_s1_t[107]), .B1_f (key_s1_f[107]), .Z0_t (KeyReg_Inst_ff_SDE_107_MUX_inst_X), .Z0_f (new_AGEMA_signal_14891), .Z1_t (new_AGEMA_signal_14892), .Z1_f (new_AGEMA_signal_14893) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_107_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_107_MUX_inst_X), .B0_f (new_AGEMA_signal_14891), .B1_t (new_AGEMA_signal_14892), .B1_f (new_AGEMA_signal_14893), .Z0_t (KeyReg_Inst_ff_SDE_107_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15635), .Z1_t (new_AGEMA_signal_15636), .Z1_f (new_AGEMA_signal_15637) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_107_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_107_MUX_inst_Y), .A0_f (new_AGEMA_signal_15635), .A1_t (new_AGEMA_signal_15636), .A1_f (new_AGEMA_signal_15637), .B0_t (KeyExpansionOutput[107]), .B0_f (new_AGEMA_signal_14045), .B1_t (new_AGEMA_signal_14046), .B1_f (new_AGEMA_signal_14047), .Z0_t (RoundKey[107]), .Z0_f (new_AGEMA_signal_5135), .Z1_t (new_AGEMA_signal_5136), .Z1_f (new_AGEMA_signal_5137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_108_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[108]), .A0_f (new_AGEMA_signal_14042), .A1_t (new_AGEMA_signal_14043), .A1_f (new_AGEMA_signal_14044), .B0_t (key_s0_t[108]), .B0_f (key_s0_f[108]), .B1_t (key_s1_t[108]), .B1_f (key_s1_f[108]), .Z0_t (KeyReg_Inst_ff_SDE_108_MUX_inst_X), .Z0_f (new_AGEMA_signal_14897), .Z1_t (new_AGEMA_signal_14898), .Z1_f (new_AGEMA_signal_14899) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_108_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_108_MUX_inst_X), .B0_f (new_AGEMA_signal_14897), .B1_t (new_AGEMA_signal_14898), .B1_f (new_AGEMA_signal_14899), .Z0_t (KeyReg_Inst_ff_SDE_108_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15638), .Z1_t (new_AGEMA_signal_15639), .Z1_f (new_AGEMA_signal_15640) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_108_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_108_MUX_inst_Y), .A0_f (new_AGEMA_signal_15638), .A1_t (new_AGEMA_signal_15639), .A1_f (new_AGEMA_signal_15640), .B0_t (KeyExpansionOutput[108]), .B0_f (new_AGEMA_signal_14042), .B1_t (new_AGEMA_signal_14043), .B1_f (new_AGEMA_signal_14044), .Z0_t (RoundKey[108]), .Z0_f (new_AGEMA_signal_5144), .Z1_t (new_AGEMA_signal_5145), .Z1_f (new_AGEMA_signal_5146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_109_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[109]), .A0_f (new_AGEMA_signal_14039), .A1_t (new_AGEMA_signal_14040), .A1_f (new_AGEMA_signal_14041), .B0_t (key_s0_t[109]), .B0_f (key_s0_f[109]), .B1_t (key_s1_t[109]), .B1_f (key_s1_f[109]), .Z0_t (KeyReg_Inst_ff_SDE_109_MUX_inst_X), .Z0_f (new_AGEMA_signal_14903), .Z1_t (new_AGEMA_signal_14904), .Z1_f (new_AGEMA_signal_14905) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_109_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_109_MUX_inst_X), .B0_f (new_AGEMA_signal_14903), .B1_t (new_AGEMA_signal_14904), .B1_f (new_AGEMA_signal_14905), .Z0_t (KeyReg_Inst_ff_SDE_109_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15641), .Z1_t (new_AGEMA_signal_15642), .Z1_f (new_AGEMA_signal_15643) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_109_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_109_MUX_inst_Y), .A0_f (new_AGEMA_signal_15641), .A1_t (new_AGEMA_signal_15642), .A1_f (new_AGEMA_signal_15643), .B0_t (KeyExpansionOutput[109]), .B0_f (new_AGEMA_signal_14039), .B1_t (new_AGEMA_signal_14040), .B1_f (new_AGEMA_signal_14041), .Z0_t (RoundKey[109]), .Z0_f (new_AGEMA_signal_5153), .Z1_t (new_AGEMA_signal_5154), .Z1_f (new_AGEMA_signal_5155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_110_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[110]), .A0_f (new_AGEMA_signal_14036), .A1_t (new_AGEMA_signal_14037), .A1_f (new_AGEMA_signal_14038), .B0_t (key_s0_t[110]), .B0_f (key_s0_f[110]), .B1_t (key_s1_t[110]), .B1_f (key_s1_f[110]), .Z0_t (KeyReg_Inst_ff_SDE_110_MUX_inst_X), .Z0_f (new_AGEMA_signal_14909), .Z1_t (new_AGEMA_signal_14910), .Z1_f (new_AGEMA_signal_14911) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_110_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_110_MUX_inst_X), .B0_f (new_AGEMA_signal_14909), .B1_t (new_AGEMA_signal_14910), .B1_f (new_AGEMA_signal_14911), .Z0_t (KeyReg_Inst_ff_SDE_110_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15644), .Z1_t (new_AGEMA_signal_15645), .Z1_f (new_AGEMA_signal_15646) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_110_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_110_MUX_inst_Y), .A0_f (new_AGEMA_signal_15644), .A1_t (new_AGEMA_signal_15645), .A1_f (new_AGEMA_signal_15646), .B0_t (KeyExpansionOutput[110]), .B0_f (new_AGEMA_signal_14036), .B1_t (new_AGEMA_signal_14037), .B1_f (new_AGEMA_signal_14038), .Z0_t (RoundKey[110]), .Z0_f (new_AGEMA_signal_5171), .Z1_t (new_AGEMA_signal_5172), .Z1_f (new_AGEMA_signal_5173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_111_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[111]), .A0_f (new_AGEMA_signal_14033), .A1_t (new_AGEMA_signal_14034), .A1_f (new_AGEMA_signal_14035), .B0_t (key_s0_t[111]), .B0_f (key_s0_f[111]), .B1_t (key_s1_t[111]), .B1_f (key_s1_f[111]), .Z0_t (KeyReg_Inst_ff_SDE_111_MUX_inst_X), .Z0_f (new_AGEMA_signal_14915), .Z1_t (new_AGEMA_signal_14916), .Z1_f (new_AGEMA_signal_14917) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_111_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_111_MUX_inst_X), .B0_f (new_AGEMA_signal_14915), .B1_t (new_AGEMA_signal_14916), .B1_f (new_AGEMA_signal_14917), .Z0_t (KeyReg_Inst_ff_SDE_111_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15647), .Z1_t (new_AGEMA_signal_15648), .Z1_f (new_AGEMA_signal_15649) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_111_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_111_MUX_inst_Y), .A0_f (new_AGEMA_signal_15647), .A1_t (new_AGEMA_signal_15648), .A1_f (new_AGEMA_signal_15649), .B0_t (KeyExpansionOutput[111]), .B0_f (new_AGEMA_signal_14033), .B1_t (new_AGEMA_signal_14034), .B1_f (new_AGEMA_signal_14035), .Z0_t (RoundKey[111]), .Z0_f (new_AGEMA_signal_5180), .Z1_t (new_AGEMA_signal_5181), .Z1_f (new_AGEMA_signal_5182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_112_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[112]), .A0_f (new_AGEMA_signal_13496), .A1_t (new_AGEMA_signal_13497), .A1_f (new_AGEMA_signal_13498), .B0_t (key_s0_t[112]), .B0_f (key_s0_f[112]), .B1_t (key_s1_t[112]), .B1_f (key_s1_f[112]), .Z0_t (KeyReg_Inst_ff_SDE_112_MUX_inst_X), .Z0_f (new_AGEMA_signal_13991), .Z1_t (new_AGEMA_signal_13992), .Z1_f (new_AGEMA_signal_13993) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_112_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_112_MUX_inst_X), .B0_f (new_AGEMA_signal_13991), .B1_t (new_AGEMA_signal_13992), .B1_f (new_AGEMA_signal_13993), .Z0_t (KeyReg_Inst_ff_SDE_112_MUX_inst_Y), .Z0_f (new_AGEMA_signal_14918), .Z1_t (new_AGEMA_signal_14919), .Z1_f (new_AGEMA_signal_14920) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_112_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_112_MUX_inst_Y), .A0_f (new_AGEMA_signal_14918), .A1_t (new_AGEMA_signal_14919), .A1_f (new_AGEMA_signal_14920), .B0_t (KeyExpansionOutput[112]), .B0_f (new_AGEMA_signal_13496), .B1_t (new_AGEMA_signal_13497), .B1_f (new_AGEMA_signal_13498), .Z0_t (RoundKey[112]), .Z0_f (new_AGEMA_signal_5189), .Z1_t (new_AGEMA_signal_5190), .Z1_f (new_AGEMA_signal_5191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_113_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[113]), .A0_f (new_AGEMA_signal_14030), .A1_t (new_AGEMA_signal_14031), .A1_f (new_AGEMA_signal_14032), .B0_t (key_s0_t[113]), .B0_f (key_s0_f[113]), .B1_t (key_s1_t[113]), .B1_f (key_s1_f[113]), .Z0_t (KeyReg_Inst_ff_SDE_113_MUX_inst_X), .Z0_f (new_AGEMA_signal_14924), .Z1_t (new_AGEMA_signal_14925), .Z1_f (new_AGEMA_signal_14926) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_113_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_113_MUX_inst_X), .B0_f (new_AGEMA_signal_14924), .B1_t (new_AGEMA_signal_14925), .B1_f (new_AGEMA_signal_14926), .Z0_t (KeyReg_Inst_ff_SDE_113_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15650), .Z1_t (new_AGEMA_signal_15651), .Z1_f (new_AGEMA_signal_15652) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_113_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_113_MUX_inst_Y), .A0_f (new_AGEMA_signal_15650), .A1_t (new_AGEMA_signal_15651), .A1_f (new_AGEMA_signal_15652), .B0_t (KeyExpansionOutput[113]), .B0_f (new_AGEMA_signal_14030), .B1_t (new_AGEMA_signal_14031), .B1_f (new_AGEMA_signal_14032), .Z0_t (RoundKey[113]), .Z0_f (new_AGEMA_signal_5198), .Z1_t (new_AGEMA_signal_5199), .Z1_f (new_AGEMA_signal_5200) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_114_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[114]), .A0_f (new_AGEMA_signal_14027), .A1_t (new_AGEMA_signal_14028), .A1_f (new_AGEMA_signal_14029), .B0_t (key_s0_t[114]), .B0_f (key_s0_f[114]), .B1_t (key_s1_t[114]), .B1_f (key_s1_f[114]), .Z0_t (KeyReg_Inst_ff_SDE_114_MUX_inst_X), .Z0_f (new_AGEMA_signal_14930), .Z1_t (new_AGEMA_signal_14931), .Z1_f (new_AGEMA_signal_14932) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_114_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_114_MUX_inst_X), .B0_f (new_AGEMA_signal_14930), .B1_t (new_AGEMA_signal_14931), .B1_f (new_AGEMA_signal_14932), .Z0_t (KeyReg_Inst_ff_SDE_114_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15653), .Z1_t (new_AGEMA_signal_15654), .Z1_f (new_AGEMA_signal_15655) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_114_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_114_MUX_inst_Y), .A0_f (new_AGEMA_signal_15653), .A1_t (new_AGEMA_signal_15654), .A1_f (new_AGEMA_signal_15655), .B0_t (KeyExpansionOutput[114]), .B0_f (new_AGEMA_signal_14027), .B1_t (new_AGEMA_signal_14028), .B1_f (new_AGEMA_signal_14029), .Z0_t (RoundKey[114]), .Z0_f (new_AGEMA_signal_5207), .Z1_t (new_AGEMA_signal_5208), .Z1_f (new_AGEMA_signal_5209) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_115_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[115]), .A0_f (new_AGEMA_signal_14024), .A1_t (new_AGEMA_signal_14025), .A1_f (new_AGEMA_signal_14026), .B0_t (key_s0_t[115]), .B0_f (key_s0_f[115]), .B1_t (key_s1_t[115]), .B1_f (key_s1_f[115]), .Z0_t (KeyReg_Inst_ff_SDE_115_MUX_inst_X), .Z0_f (new_AGEMA_signal_14936), .Z1_t (new_AGEMA_signal_14937), .Z1_f (new_AGEMA_signal_14938) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_115_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_115_MUX_inst_X), .B0_f (new_AGEMA_signal_14936), .B1_t (new_AGEMA_signal_14937), .B1_f (new_AGEMA_signal_14938), .Z0_t (KeyReg_Inst_ff_SDE_115_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15656), .Z1_t (new_AGEMA_signal_15657), .Z1_f (new_AGEMA_signal_15658) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_115_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_115_MUX_inst_Y), .A0_f (new_AGEMA_signal_15656), .A1_t (new_AGEMA_signal_15657), .A1_f (new_AGEMA_signal_15658), .B0_t (KeyExpansionOutput[115]), .B0_f (new_AGEMA_signal_14024), .B1_t (new_AGEMA_signal_14025), .B1_f (new_AGEMA_signal_14026), .Z0_t (RoundKey[115]), .Z0_f (new_AGEMA_signal_5216), .Z1_t (new_AGEMA_signal_5217), .Z1_f (new_AGEMA_signal_5218) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_116_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[116]), .A0_f (new_AGEMA_signal_14021), .A1_t (new_AGEMA_signal_14022), .A1_f (new_AGEMA_signal_14023), .B0_t (key_s0_t[116]), .B0_f (key_s0_f[116]), .B1_t (key_s1_t[116]), .B1_f (key_s1_f[116]), .Z0_t (KeyReg_Inst_ff_SDE_116_MUX_inst_X), .Z0_f (new_AGEMA_signal_14942), .Z1_t (new_AGEMA_signal_14943), .Z1_f (new_AGEMA_signal_14944) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_116_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_116_MUX_inst_X), .B0_f (new_AGEMA_signal_14942), .B1_t (new_AGEMA_signal_14943), .B1_f (new_AGEMA_signal_14944), .Z0_t (KeyReg_Inst_ff_SDE_116_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15659), .Z1_t (new_AGEMA_signal_15660), .Z1_f (new_AGEMA_signal_15661) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_116_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_116_MUX_inst_Y), .A0_f (new_AGEMA_signal_15659), .A1_t (new_AGEMA_signal_15660), .A1_f (new_AGEMA_signal_15661), .B0_t (KeyExpansionOutput[116]), .B0_f (new_AGEMA_signal_14021), .B1_t (new_AGEMA_signal_14022), .B1_f (new_AGEMA_signal_14023), .Z0_t (RoundKey[116]), .Z0_f (new_AGEMA_signal_5225), .Z1_t (new_AGEMA_signal_5226), .Z1_f (new_AGEMA_signal_5227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_117_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[117]), .A0_f (new_AGEMA_signal_14018), .A1_t (new_AGEMA_signal_14019), .A1_f (new_AGEMA_signal_14020), .B0_t (key_s0_t[117]), .B0_f (key_s0_f[117]), .B1_t (key_s1_t[117]), .B1_f (key_s1_f[117]), .Z0_t (KeyReg_Inst_ff_SDE_117_MUX_inst_X), .Z0_f (new_AGEMA_signal_14948), .Z1_t (new_AGEMA_signal_14949), .Z1_f (new_AGEMA_signal_14950) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_117_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_117_MUX_inst_X), .B0_f (new_AGEMA_signal_14948), .B1_t (new_AGEMA_signal_14949), .B1_f (new_AGEMA_signal_14950), .Z0_t (KeyReg_Inst_ff_SDE_117_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15662), .Z1_t (new_AGEMA_signal_15663), .Z1_f (new_AGEMA_signal_15664) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_117_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_117_MUX_inst_Y), .A0_f (new_AGEMA_signal_15662), .A1_t (new_AGEMA_signal_15663), .A1_f (new_AGEMA_signal_15664), .B0_t (KeyExpansionOutput[117]), .B0_f (new_AGEMA_signal_14018), .B1_t (new_AGEMA_signal_14019), .B1_f (new_AGEMA_signal_14020), .Z0_t (RoundKey[117]), .Z0_f (new_AGEMA_signal_5234), .Z1_t (new_AGEMA_signal_5235), .Z1_f (new_AGEMA_signal_5236) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_118_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[118]), .A0_f (new_AGEMA_signal_14015), .A1_t (new_AGEMA_signal_14016), .A1_f (new_AGEMA_signal_14017), .B0_t (key_s0_t[118]), .B0_f (key_s0_f[118]), .B1_t (key_s1_t[118]), .B1_f (key_s1_f[118]), .Z0_t (KeyReg_Inst_ff_SDE_118_MUX_inst_X), .Z0_f (new_AGEMA_signal_14954), .Z1_t (new_AGEMA_signal_14955), .Z1_f (new_AGEMA_signal_14956) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_118_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_118_MUX_inst_X), .B0_f (new_AGEMA_signal_14954), .B1_t (new_AGEMA_signal_14955), .B1_f (new_AGEMA_signal_14956), .Z0_t (KeyReg_Inst_ff_SDE_118_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15665), .Z1_t (new_AGEMA_signal_15666), .Z1_f (new_AGEMA_signal_15667) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_118_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_118_MUX_inst_Y), .A0_f (new_AGEMA_signal_15665), .A1_t (new_AGEMA_signal_15666), .A1_f (new_AGEMA_signal_15667), .B0_t (KeyExpansionOutput[118]), .B0_f (new_AGEMA_signal_14015), .B1_t (new_AGEMA_signal_14016), .B1_f (new_AGEMA_signal_14017), .Z0_t (RoundKey[118]), .Z0_f (new_AGEMA_signal_5243), .Z1_t (new_AGEMA_signal_5244), .Z1_f (new_AGEMA_signal_5245) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_119_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[119]), .A0_f (new_AGEMA_signal_14012), .A1_t (new_AGEMA_signal_14013), .A1_f (new_AGEMA_signal_14014), .B0_t (key_s0_t[119]), .B0_f (key_s0_f[119]), .B1_t (key_s1_t[119]), .B1_f (key_s1_f[119]), .Z0_t (KeyReg_Inst_ff_SDE_119_MUX_inst_X), .Z0_f (new_AGEMA_signal_14960), .Z1_t (new_AGEMA_signal_14961), .Z1_f (new_AGEMA_signal_14962) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_119_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_119_MUX_inst_X), .B0_f (new_AGEMA_signal_14960), .B1_t (new_AGEMA_signal_14961), .B1_f (new_AGEMA_signal_14962), .Z0_t (KeyReg_Inst_ff_SDE_119_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15668), .Z1_t (new_AGEMA_signal_15669), .Z1_f (new_AGEMA_signal_15670) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_119_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_119_MUX_inst_Y), .A0_f (new_AGEMA_signal_15668), .A1_t (new_AGEMA_signal_15669), .A1_f (new_AGEMA_signal_15670), .B0_t (KeyExpansionOutput[119]), .B0_f (new_AGEMA_signal_14012), .B1_t (new_AGEMA_signal_14013), .B1_f (new_AGEMA_signal_14014), .Z0_t (RoundKey[119]), .Z0_f (new_AGEMA_signal_5252), .Z1_t (new_AGEMA_signal_5253), .Z1_f (new_AGEMA_signal_5254) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_120_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[120]), .A0_f (new_AGEMA_signal_14009), .A1_t (new_AGEMA_signal_14010), .A1_f (new_AGEMA_signal_14011), .B0_t (key_s0_t[120]), .B0_f (key_s0_f[120]), .B1_t (key_s1_t[120]), .B1_f (key_s1_f[120]), .Z0_t (KeyReg_Inst_ff_SDE_120_MUX_inst_X), .Z0_f (new_AGEMA_signal_14966), .Z1_t (new_AGEMA_signal_14967), .Z1_f (new_AGEMA_signal_14968) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_120_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_120_MUX_inst_X), .B0_f (new_AGEMA_signal_14966), .B1_t (new_AGEMA_signal_14967), .B1_f (new_AGEMA_signal_14968), .Z0_t (KeyReg_Inst_ff_SDE_120_MUX_inst_Y), .Z0_f (new_AGEMA_signal_15671), .Z1_t (new_AGEMA_signal_15672), .Z1_f (new_AGEMA_signal_15673) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_120_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_120_MUX_inst_Y), .A0_f (new_AGEMA_signal_15671), .A1_t (new_AGEMA_signal_15672), .A1_f (new_AGEMA_signal_15673), .B0_t (KeyExpansionOutput[120]), .B0_f (new_AGEMA_signal_14009), .B1_t (new_AGEMA_signal_14010), .B1_f (new_AGEMA_signal_14011), .Z0_t (RoundKey[120]), .Z0_f (new_AGEMA_signal_5270), .Z1_t (new_AGEMA_signal_5271), .Z1_f (new_AGEMA_signal_5272) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_121_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[121]), .A0_f (new_AGEMA_signal_15053), .A1_t (new_AGEMA_signal_15054), .A1_f (new_AGEMA_signal_15055), .B0_t (key_s0_t[121]), .B0_f (key_s0_f[121]), .B1_t (key_s1_t[121]), .B1_f (key_s1_f[121]), .Z0_t (KeyReg_Inst_ff_SDE_121_MUX_inst_X), .Z0_f (new_AGEMA_signal_15677), .Z1_t (new_AGEMA_signal_15678), .Z1_f (new_AGEMA_signal_15679) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_121_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_121_MUX_inst_X), .B0_f (new_AGEMA_signal_15677), .B1_t (new_AGEMA_signal_15678), .B1_f (new_AGEMA_signal_15679), .Z0_t (KeyReg_Inst_ff_SDE_121_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16463), .Z1_t (new_AGEMA_signal_16464), .Z1_f (new_AGEMA_signal_16465) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_121_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_121_MUX_inst_Y), .A0_f (new_AGEMA_signal_16463), .A1_t (new_AGEMA_signal_16464), .A1_f (new_AGEMA_signal_16465), .B0_t (KeyExpansionOutput[121]), .B0_f (new_AGEMA_signal_15053), .B1_t (new_AGEMA_signal_15054), .B1_f (new_AGEMA_signal_15055), .Z0_t (RoundKey[121]), .Z0_f (new_AGEMA_signal_5279), .Z1_t (new_AGEMA_signal_5280), .Z1_f (new_AGEMA_signal_5281) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_122_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[122]), .A0_f (new_AGEMA_signal_15050), .A1_t (new_AGEMA_signal_15051), .A1_f (new_AGEMA_signal_15052), .B0_t (key_s0_t[122]), .B0_f (key_s0_f[122]), .B1_t (key_s1_t[122]), .B1_f (key_s1_f[122]), .Z0_t (KeyReg_Inst_ff_SDE_122_MUX_inst_X), .Z0_f (new_AGEMA_signal_15683), .Z1_t (new_AGEMA_signal_15684), .Z1_f (new_AGEMA_signal_15685) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_122_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_122_MUX_inst_X), .B0_f (new_AGEMA_signal_15683), .B1_t (new_AGEMA_signal_15684), .B1_f (new_AGEMA_signal_15685), .Z0_t (KeyReg_Inst_ff_SDE_122_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16466), .Z1_t (new_AGEMA_signal_16467), .Z1_f (new_AGEMA_signal_16468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_122_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_122_MUX_inst_Y), .A0_f (new_AGEMA_signal_16466), .A1_t (new_AGEMA_signal_16467), .A1_f (new_AGEMA_signal_16468), .B0_t (KeyExpansionOutput[122]), .B0_f (new_AGEMA_signal_15050), .B1_t (new_AGEMA_signal_15051), .B1_f (new_AGEMA_signal_15052), .Z0_t (RoundKey[122]), .Z0_f (new_AGEMA_signal_5288), .Z1_t (new_AGEMA_signal_5289), .Z1_f (new_AGEMA_signal_5290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_123_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[123]), .A0_f (new_AGEMA_signal_15047), .A1_t (new_AGEMA_signal_15048), .A1_f (new_AGEMA_signal_15049), .B0_t (key_s0_t[123]), .B0_f (key_s0_f[123]), .B1_t (key_s1_t[123]), .B1_f (key_s1_f[123]), .Z0_t (KeyReg_Inst_ff_SDE_123_MUX_inst_X), .Z0_f (new_AGEMA_signal_15689), .Z1_t (new_AGEMA_signal_15690), .Z1_f (new_AGEMA_signal_15691) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_123_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_123_MUX_inst_X), .B0_f (new_AGEMA_signal_15689), .B1_t (new_AGEMA_signal_15690), .B1_f (new_AGEMA_signal_15691), .Z0_t (KeyReg_Inst_ff_SDE_123_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16469), .Z1_t (new_AGEMA_signal_16470), .Z1_f (new_AGEMA_signal_16471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_123_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_123_MUX_inst_Y), .A0_f (new_AGEMA_signal_16469), .A1_t (new_AGEMA_signal_16470), .A1_f (new_AGEMA_signal_16471), .B0_t (KeyExpansionOutput[123]), .B0_f (new_AGEMA_signal_15047), .B1_t (new_AGEMA_signal_15048), .B1_f (new_AGEMA_signal_15049), .Z0_t (RoundKey[123]), .Z0_f (new_AGEMA_signal_5297), .Z1_t (new_AGEMA_signal_5298), .Z1_f (new_AGEMA_signal_5299) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_124_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[124]), .A0_f (new_AGEMA_signal_15044), .A1_t (new_AGEMA_signal_15045), .A1_f (new_AGEMA_signal_15046), .B0_t (key_s0_t[124]), .B0_f (key_s0_f[124]), .B1_t (key_s1_t[124]), .B1_f (key_s1_f[124]), .Z0_t (KeyReg_Inst_ff_SDE_124_MUX_inst_X), .Z0_f (new_AGEMA_signal_15695), .Z1_t (new_AGEMA_signal_15696), .Z1_f (new_AGEMA_signal_15697) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_124_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_124_MUX_inst_X), .B0_f (new_AGEMA_signal_15695), .B1_t (new_AGEMA_signal_15696), .B1_f (new_AGEMA_signal_15697), .Z0_t (KeyReg_Inst_ff_SDE_124_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16472), .Z1_t (new_AGEMA_signal_16473), .Z1_f (new_AGEMA_signal_16474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_124_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_124_MUX_inst_Y), .A0_f (new_AGEMA_signal_16472), .A1_t (new_AGEMA_signal_16473), .A1_f (new_AGEMA_signal_16474), .B0_t (KeyExpansionOutput[124]), .B0_f (new_AGEMA_signal_15044), .B1_t (new_AGEMA_signal_15045), .B1_f (new_AGEMA_signal_15046), .Z0_t (RoundKey[124]), .Z0_f (new_AGEMA_signal_5306), .Z1_t (new_AGEMA_signal_5307), .Z1_f (new_AGEMA_signal_5308) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_125_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[125]), .A0_f (new_AGEMA_signal_15041), .A1_t (new_AGEMA_signal_15042), .A1_f (new_AGEMA_signal_15043), .B0_t (key_s0_t[125]), .B0_f (key_s0_f[125]), .B1_t (key_s1_t[125]), .B1_f (key_s1_f[125]), .Z0_t (KeyReg_Inst_ff_SDE_125_MUX_inst_X), .Z0_f (new_AGEMA_signal_15701), .Z1_t (new_AGEMA_signal_15702), .Z1_f (new_AGEMA_signal_15703) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_125_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_125_MUX_inst_X), .B0_f (new_AGEMA_signal_15701), .B1_t (new_AGEMA_signal_15702), .B1_f (new_AGEMA_signal_15703), .Z0_t (KeyReg_Inst_ff_SDE_125_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16475), .Z1_t (new_AGEMA_signal_16476), .Z1_f (new_AGEMA_signal_16477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_125_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_125_MUX_inst_Y), .A0_f (new_AGEMA_signal_16475), .A1_t (new_AGEMA_signal_16476), .A1_f (new_AGEMA_signal_16477), .B0_t (KeyExpansionOutput[125]), .B0_f (new_AGEMA_signal_15041), .B1_t (new_AGEMA_signal_15042), .B1_f (new_AGEMA_signal_15043), .Z0_t (RoundKey[125]), .Z0_f (new_AGEMA_signal_5315), .Z1_t (new_AGEMA_signal_5316), .Z1_f (new_AGEMA_signal_5317) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_126_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[126]), .A0_f (new_AGEMA_signal_15038), .A1_t (new_AGEMA_signal_15039), .A1_f (new_AGEMA_signal_15040), .B0_t (key_s0_t[126]), .B0_f (key_s0_f[126]), .B1_t (key_s1_t[126]), .B1_f (key_s1_f[126]), .Z0_t (KeyReg_Inst_ff_SDE_126_MUX_inst_X), .Z0_f (new_AGEMA_signal_15707), .Z1_t (new_AGEMA_signal_15708), .Z1_f (new_AGEMA_signal_15709) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_126_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_126_MUX_inst_X), .B0_f (new_AGEMA_signal_15707), .B1_t (new_AGEMA_signal_15708), .B1_f (new_AGEMA_signal_15709), .Z0_t (KeyReg_Inst_ff_SDE_126_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16478), .Z1_t (new_AGEMA_signal_16479), .Z1_f (new_AGEMA_signal_16480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_126_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_126_MUX_inst_Y), .A0_f (new_AGEMA_signal_16478), .A1_t (new_AGEMA_signal_16479), .A1_f (new_AGEMA_signal_16480), .B0_t (KeyExpansionOutput[126]), .B0_f (new_AGEMA_signal_15038), .B1_t (new_AGEMA_signal_15039), .B1_f (new_AGEMA_signal_15040), .Z0_t (RoundKey[126]), .Z0_f (new_AGEMA_signal_5324), .Z1_t (new_AGEMA_signal_5325), .Z1_f (new_AGEMA_signal_5326) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_127_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[127]), .A0_f (new_AGEMA_signal_15035), .A1_t (new_AGEMA_signal_15036), .A1_f (new_AGEMA_signal_15037), .B0_t (key_s0_t[127]), .B0_f (key_s0_f[127]), .B1_t (key_s1_t[127]), .B1_f (key_s1_f[127]), .Z0_t (KeyReg_Inst_ff_SDE_127_MUX_inst_X), .Z0_f (new_AGEMA_signal_15713), .Z1_t (new_AGEMA_signal_15714), .Z1_f (new_AGEMA_signal_15715) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_127_MUX_inst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyReg_Inst_ff_SDE_127_MUX_inst_X), .B0_f (new_AGEMA_signal_15713), .B1_t (new_AGEMA_signal_15714), .B1_f (new_AGEMA_signal_15715), .Z0_t (KeyReg_Inst_ff_SDE_127_MUX_inst_Y), .Z0_f (new_AGEMA_signal_16481), .Z1_t (new_AGEMA_signal_16482), .Z1_f (new_AGEMA_signal_16483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_127_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_127_MUX_inst_Y), .A0_f (new_AGEMA_signal_16481), .A1_t (new_AGEMA_signal_16482), .A1_f (new_AGEMA_signal_16483), .B0_t (KeyExpansionOutput[127]), .B0_f (new_AGEMA_signal_15035), .B1_t (new_AGEMA_signal_15036), .B1_f (new_AGEMA_signal_15037), .Z0_t (RoundKey[127]), .Z0_f (new_AGEMA_signal_5333), .Z1_t (new_AGEMA_signal_5334), .Z1_f (new_AGEMA_signal_5335) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U128 ( .A0_t (RoundKey[9]), .A0_f (new_AGEMA_signal_6206), .A1_t (new_AGEMA_signal_6207), .A1_f (new_AGEMA_signal_6208), .B0_t (KeyExpansionOutput[41]), .B0_f (new_AGEMA_signal_15719), .B1_t (new_AGEMA_signal_15720), .B1_f (new_AGEMA_signal_15721), .Z0_t (KeyExpansionOutput[9]), .Z0_f (new_AGEMA_signal_16484), .Z1_t (new_AGEMA_signal_16485), .Z1_f (new_AGEMA_signal_16486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U127 ( .A0_t (RoundKey[8]), .A0_f (new_AGEMA_signal_6107), .A1_t (new_AGEMA_signal_6108), .A1_f (new_AGEMA_signal_6109), .B0_t (KeyExpansionOutput[40]), .B0_f (new_AGEMA_signal_14972), .B1_t (new_AGEMA_signal_14973), .B1_f (new_AGEMA_signal_14974), .Z0_t (KeyExpansionOutput[8]), .Z0_f (new_AGEMA_signal_15716), .Z1_t (new_AGEMA_signal_15717), .Z1_f (new_AGEMA_signal_15718) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U126 ( .A0_t (RoundKey[7]), .A0_f (new_AGEMA_signal_6008), .A1_t (new_AGEMA_signal_6009), .A1_f (new_AGEMA_signal_6010), .B0_t (KeyExpansionOutput[39]), .B0_f (new_AGEMA_signal_15722), .B1_t (new_AGEMA_signal_15723), .B1_f (new_AGEMA_signal_15724), .Z0_t (KeyExpansionOutput[7]), .Z0_f (new_AGEMA_signal_16487), .Z1_t (new_AGEMA_signal_16488), .Z1_f (new_AGEMA_signal_16489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U125 ( .A0_t (RoundKey[6]), .A0_f (new_AGEMA_signal_5909), .A1_t (new_AGEMA_signal_5910), .A1_f (new_AGEMA_signal_5911), .B0_t (KeyExpansionOutput[38]), .B0_f (new_AGEMA_signal_15725), .B1_t (new_AGEMA_signal_15726), .B1_f (new_AGEMA_signal_15727), .Z0_t (KeyExpansionOutput[6]), .Z0_f (new_AGEMA_signal_16490), .Z1_t (new_AGEMA_signal_16491), .Z1_f (new_AGEMA_signal_16492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U124 ( .A0_t (RoundKey[5]), .A0_f (new_AGEMA_signal_5810), .A1_t (new_AGEMA_signal_5811), .A1_f (new_AGEMA_signal_5812), .B0_t (KeyExpansionOutput[37]), .B0_f (new_AGEMA_signal_15728), .B1_t (new_AGEMA_signal_15729), .B1_f (new_AGEMA_signal_15730), .Z0_t (KeyExpansionOutput[5]), .Z0_f (new_AGEMA_signal_16493), .Z1_t (new_AGEMA_signal_16494), .Z1_f (new_AGEMA_signal_16495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U123 ( .A0_t (RoundKey[4]), .A0_f (new_AGEMA_signal_5711), .A1_t (new_AGEMA_signal_5712), .A1_f (new_AGEMA_signal_5713), .B0_t (KeyExpansionOutput[36]), .B0_f (new_AGEMA_signal_15731), .B1_t (new_AGEMA_signal_15732), .B1_f (new_AGEMA_signal_15733), .Z0_t (KeyExpansionOutput[4]), .Z0_f (new_AGEMA_signal_16496), .Z1_t (new_AGEMA_signal_16497), .Z1_f (new_AGEMA_signal_16498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U122 ( .A0_t (RoundKey[41]), .A0_f (new_AGEMA_signal_5630), .A1_t (new_AGEMA_signal_5631), .A1_f (new_AGEMA_signal_5632), .B0_t (KeyExpansionOutput[73]), .B0_f (new_AGEMA_signal_14969), .B1_t (new_AGEMA_signal_14970), .B1_f (new_AGEMA_signal_14971), .Z0_t (KeyExpansionOutput[41]), .Z0_f (new_AGEMA_signal_15719), .Z1_t (new_AGEMA_signal_15720), .Z1_f (new_AGEMA_signal_15721) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U121 ( .A0_t (RoundKey[73]), .A0_f (new_AGEMA_signal_5945), .A1_t (new_AGEMA_signal_5946), .A1_f (new_AGEMA_signal_5947), .B0_t (KeyExpansionOutput[105]), .B0_f (new_AGEMA_signal_14051), .B1_t (new_AGEMA_signal_14052), .B1_f (new_AGEMA_signal_14053), .Z0_t (KeyExpansionOutput[73]), .Z0_f (new_AGEMA_signal_14969), .Z1_t (new_AGEMA_signal_14970), .Z1_f (new_AGEMA_signal_14971) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U120 ( .A0_t (RoundKey[40]), .A0_f (new_AGEMA_signal_5621), .A1_t (new_AGEMA_signal_5622), .A1_f (new_AGEMA_signal_5623), .B0_t (KeyExpansionOutput[72]), .B0_f (new_AGEMA_signal_13994), .B1_t (new_AGEMA_signal_13995), .B1_f (new_AGEMA_signal_13996), .Z0_t (KeyExpansionOutput[40]), .Z0_f (new_AGEMA_signal_14972), .Z1_t (new_AGEMA_signal_14973), .Z1_f (new_AGEMA_signal_14974) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U119 ( .A0_t (RoundKey[72]), .A0_f (new_AGEMA_signal_5936), .A1_t (new_AGEMA_signal_5937), .A1_f (new_AGEMA_signal_5938), .B0_t (KeyExpansionOutput[104]), .B0_f (new_AGEMA_signal_13499), .B1_t (new_AGEMA_signal_13500), .B1_f (new_AGEMA_signal_13501), .Z0_t (KeyExpansionOutput[72]), .Z0_f (new_AGEMA_signal_13994), .Z1_t (new_AGEMA_signal_13995), .Z1_f (new_AGEMA_signal_13996) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U118 ( .A0_t (RoundKey[3]), .A0_f (new_AGEMA_signal_5612), .A1_t (new_AGEMA_signal_5613), .A1_f (new_AGEMA_signal_5614), .B0_t (KeyExpansionOutput[35]), .B0_f (new_AGEMA_signal_15734), .B1_t (new_AGEMA_signal_15735), .B1_f (new_AGEMA_signal_15736), .Z0_t (KeyExpansionOutput[3]), .Z0_f (new_AGEMA_signal_16499), .Z1_t (new_AGEMA_signal_16500), .Z1_f (new_AGEMA_signal_16501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U117 ( .A0_t (RoundKey[39]), .A0_f (new_AGEMA_signal_5603), .A1_t (new_AGEMA_signal_5604), .A1_f (new_AGEMA_signal_5605), .B0_t (KeyExpansionOutput[71]), .B0_f (new_AGEMA_signal_14975), .B1_t (new_AGEMA_signal_14976), .B1_f (new_AGEMA_signal_14977), .Z0_t (KeyExpansionOutput[39]), .Z0_f (new_AGEMA_signal_15722), .Z1_t (new_AGEMA_signal_15723), .Z1_f (new_AGEMA_signal_15724) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U116 ( .A0_t (RoundKey[71]), .A0_f (new_AGEMA_signal_5927), .A1_t (new_AGEMA_signal_5928), .A1_f (new_AGEMA_signal_5929), .B0_t (KeyExpansionOutput[103]), .B0_f (new_AGEMA_signal_14054), .B1_t (new_AGEMA_signal_14055), .B1_f (new_AGEMA_signal_14056), .Z0_t (KeyExpansionOutput[71]), .Z0_f (new_AGEMA_signal_14975), .Z1_t (new_AGEMA_signal_14976), .Z1_f (new_AGEMA_signal_14977) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U115 ( .A0_t (RoundKey[38]), .A0_f (new_AGEMA_signal_5594), .A1_t (new_AGEMA_signal_5595), .A1_f (new_AGEMA_signal_5596), .B0_t (KeyExpansionOutput[70]), .B0_f (new_AGEMA_signal_14978), .B1_t (new_AGEMA_signal_14979), .B1_f (new_AGEMA_signal_14980), .Z0_t (KeyExpansionOutput[38]), .Z0_f (new_AGEMA_signal_15725), .Z1_t (new_AGEMA_signal_15726), .Z1_f (new_AGEMA_signal_15727) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U114 ( .A0_t (RoundKey[70]), .A0_f (new_AGEMA_signal_5918), .A1_t (new_AGEMA_signal_5919), .A1_f (new_AGEMA_signal_5920), .B0_t (KeyExpansionOutput[102]), .B0_f (new_AGEMA_signal_14057), .B1_t (new_AGEMA_signal_14058), .B1_f (new_AGEMA_signal_14059), .Z0_t (KeyExpansionOutput[70]), .Z0_f (new_AGEMA_signal_14978), .Z1_t (new_AGEMA_signal_14979), .Z1_f (new_AGEMA_signal_14980) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U113 ( .A0_t (RoundKey[37]), .A0_f (new_AGEMA_signal_5585), .A1_t (new_AGEMA_signal_5586), .A1_f (new_AGEMA_signal_5587), .B0_t (KeyExpansionOutput[69]), .B0_f (new_AGEMA_signal_14981), .B1_t (new_AGEMA_signal_14982), .B1_f (new_AGEMA_signal_14983), .Z0_t (KeyExpansionOutput[37]), .Z0_f (new_AGEMA_signal_15728), .Z1_t (new_AGEMA_signal_15729), .Z1_f (new_AGEMA_signal_15730) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U112 ( .A0_t (RoundKey[69]), .A0_f (new_AGEMA_signal_5900), .A1_t (new_AGEMA_signal_5901), .A1_f (new_AGEMA_signal_5902), .B0_t (KeyExpansionOutput[101]), .B0_f (new_AGEMA_signal_14060), .B1_t (new_AGEMA_signal_14061), .B1_f (new_AGEMA_signal_14062), .Z0_t (KeyExpansionOutput[69]), .Z0_f (new_AGEMA_signal_14981), .Z1_t (new_AGEMA_signal_14982), .Z1_f (new_AGEMA_signal_14983) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U111 ( .A0_t (RoundKey[36]), .A0_f (new_AGEMA_signal_5576), .A1_t (new_AGEMA_signal_5577), .A1_f (new_AGEMA_signal_5578), .B0_t (KeyExpansionOutput[68]), .B0_f (new_AGEMA_signal_14984), .B1_t (new_AGEMA_signal_14985), .B1_f (new_AGEMA_signal_14986), .Z0_t (KeyExpansionOutput[36]), .Z0_f (new_AGEMA_signal_15731), .Z1_t (new_AGEMA_signal_15732), .Z1_f (new_AGEMA_signal_15733) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U110 ( .A0_t (RoundKey[68]), .A0_f (new_AGEMA_signal_5891), .A1_t (new_AGEMA_signal_5892), .A1_f (new_AGEMA_signal_5893), .B0_t (KeyExpansionOutput[100]), .B0_f (new_AGEMA_signal_14063), .B1_t (new_AGEMA_signal_14064), .B1_f (new_AGEMA_signal_14065), .Z0_t (KeyExpansionOutput[68]), .Z0_f (new_AGEMA_signal_14984), .Z1_t (new_AGEMA_signal_14985), .Z1_f (new_AGEMA_signal_14986) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U109 ( .A0_t (RoundKey[35]), .A0_f (new_AGEMA_signal_5567), .A1_t (new_AGEMA_signal_5568), .A1_f (new_AGEMA_signal_5569), .B0_t (KeyExpansionOutput[67]), .B0_f (new_AGEMA_signal_14987), .B1_t (new_AGEMA_signal_14988), .B1_f (new_AGEMA_signal_14989), .Z0_t (KeyExpansionOutput[35]), .Z0_f (new_AGEMA_signal_15734), .Z1_t (new_AGEMA_signal_15735), .Z1_f (new_AGEMA_signal_15736) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U108 ( .A0_t (RoundKey[67]), .A0_f (new_AGEMA_signal_5882), .A1_t (new_AGEMA_signal_5883), .A1_f (new_AGEMA_signal_5884), .B0_t (KeyExpansionOutput[99]), .B0_f (new_AGEMA_signal_13997), .B1_t (new_AGEMA_signal_13998), .B1_f (new_AGEMA_signal_13999), .Z0_t (KeyExpansionOutput[67]), .Z0_f (new_AGEMA_signal_14987), .Z1_t (new_AGEMA_signal_14988), .Z1_f (new_AGEMA_signal_14989) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U107 ( .A0_t (RoundKey[99]), .A0_f (new_AGEMA_signal_6197), .A1_t (new_AGEMA_signal_6198), .A1_f (new_AGEMA_signal_6199), .B0_t (KeyExpansionIns_tmp[3]), .B0_f (new_AGEMA_signal_13583), .B1_t (new_AGEMA_signal_13584), .B1_f (new_AGEMA_signal_13585), .Z0_t (KeyExpansionOutput[99]), .Z0_f (new_AGEMA_signal_13997), .Z1_t (new_AGEMA_signal_13998), .Z1_f (new_AGEMA_signal_13999) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U106 ( .A0_t (RoundKey[31]), .A0_f (new_AGEMA_signal_5531), .A1_t (new_AGEMA_signal_5532), .A1_f (new_AGEMA_signal_5533), .B0_t (KeyExpansionOutput[63]), .B0_f (new_AGEMA_signal_16502), .B1_t (new_AGEMA_signal_16503), .B1_f (new_AGEMA_signal_16504), .Z0_t (KeyExpansionOutput[31]), .Z0_f (new_AGEMA_signal_17225), .Z1_t (new_AGEMA_signal_17226), .Z1_f (new_AGEMA_signal_17227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U105 ( .A0_t (RoundKey[63]), .A0_f (new_AGEMA_signal_5846), .A1_t (new_AGEMA_signal_5847), .A1_f (new_AGEMA_signal_5848), .B0_t (KeyExpansionOutput[95]), .B0_f (new_AGEMA_signal_15737), .B1_t (new_AGEMA_signal_15738), .B1_f (new_AGEMA_signal_15739), .Z0_t (KeyExpansionOutput[63]), .Z0_f (new_AGEMA_signal_16502), .Z1_t (new_AGEMA_signal_16503), .Z1_f (new_AGEMA_signal_16504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U104 ( .A0_t (RoundKey[95]), .A0_f (new_AGEMA_signal_6161), .A1_t (new_AGEMA_signal_6162), .A1_f (new_AGEMA_signal_6163), .B0_t (KeyExpansionOutput[127]), .B0_f (new_AGEMA_signal_15035), .B1_t (new_AGEMA_signal_15036), .B1_f (new_AGEMA_signal_15037), .Z0_t (KeyExpansionOutput[95]), .Z0_f (new_AGEMA_signal_15737), .Z1_t (new_AGEMA_signal_15738), .Z1_f (new_AGEMA_signal_15739) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U103 ( .A0_t (RoundKey[30]), .A0_f (new_AGEMA_signal_5522), .A1_t (new_AGEMA_signal_5523), .A1_f (new_AGEMA_signal_5524), .B0_t (KeyExpansionOutput[62]), .B0_f (new_AGEMA_signal_16505), .B1_t (new_AGEMA_signal_16506), .B1_f (new_AGEMA_signal_16507), .Z0_t (KeyExpansionOutput[30]), .Z0_f (new_AGEMA_signal_17228), .Z1_t (new_AGEMA_signal_17229), .Z1_f (new_AGEMA_signal_17230) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U102 ( .A0_t (RoundKey[62]), .A0_f (new_AGEMA_signal_5837), .A1_t (new_AGEMA_signal_5838), .A1_f (new_AGEMA_signal_5839), .B0_t (KeyExpansionOutput[94]), .B0_f (new_AGEMA_signal_15740), .B1_t (new_AGEMA_signal_15741), .B1_f (new_AGEMA_signal_15742), .Z0_t (KeyExpansionOutput[62]), .Z0_f (new_AGEMA_signal_16505), .Z1_t (new_AGEMA_signal_16506), .Z1_f (new_AGEMA_signal_16507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U101 ( .A0_t (RoundKey[94]), .A0_f (new_AGEMA_signal_6152), .A1_t (new_AGEMA_signal_6153), .A1_f (new_AGEMA_signal_6154), .B0_t (KeyExpansionOutput[126]), .B0_f (new_AGEMA_signal_15038), .B1_t (new_AGEMA_signal_15039), .B1_f (new_AGEMA_signal_15040), .Z0_t (KeyExpansionOutput[94]), .Z0_f (new_AGEMA_signal_15740), .Z1_t (new_AGEMA_signal_15741), .Z1_f (new_AGEMA_signal_15742) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U100 ( .A0_t (RoundKey[2]), .A0_f (new_AGEMA_signal_5513), .A1_t (new_AGEMA_signal_5514), .A1_f (new_AGEMA_signal_5515), .B0_t (KeyExpansionOutput[34]), .B0_f (new_AGEMA_signal_15743), .B1_t (new_AGEMA_signal_15744), .B1_f (new_AGEMA_signal_15745), .Z0_t (KeyExpansionOutput[2]), .Z0_f (new_AGEMA_signal_16508), .Z1_t (new_AGEMA_signal_16509), .Z1_f (new_AGEMA_signal_16510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U99 ( .A0_t (RoundKey[34]), .A0_f (new_AGEMA_signal_5558), .A1_t (new_AGEMA_signal_5559), .A1_f (new_AGEMA_signal_5560), .B0_t (KeyExpansionOutput[66]), .B0_f (new_AGEMA_signal_14990), .B1_t (new_AGEMA_signal_14991), .B1_f (new_AGEMA_signal_14992), .Z0_t (KeyExpansionOutput[34]), .Z0_f (new_AGEMA_signal_15743), .Z1_t (new_AGEMA_signal_15744), .Z1_f (new_AGEMA_signal_15745) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U98 ( .A0_t (RoundKey[66]), .A0_f (new_AGEMA_signal_5873), .A1_t (new_AGEMA_signal_5874), .A1_f (new_AGEMA_signal_5875), .B0_t (KeyExpansionOutput[98]), .B0_f (new_AGEMA_signal_14000), .B1_t (new_AGEMA_signal_14001), .B1_f (new_AGEMA_signal_14002), .Z0_t (KeyExpansionOutput[66]), .Z0_f (new_AGEMA_signal_14990), .Z1_t (new_AGEMA_signal_14991), .Z1_f (new_AGEMA_signal_14992) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U97 ( .A0_t (RoundKey[98]), .A0_f (new_AGEMA_signal_6188), .A1_t (new_AGEMA_signal_6189), .A1_f (new_AGEMA_signal_6190), .B0_t (KeyExpansionIns_tmp[2]), .B0_f (new_AGEMA_signal_13586), .B1_t (new_AGEMA_signal_13587), .B1_f (new_AGEMA_signal_13588), .Z0_t (KeyExpansionOutput[98]), .Z0_f (new_AGEMA_signal_14000), .Z1_t (new_AGEMA_signal_14001), .Z1_f (new_AGEMA_signal_14002) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U96 ( .A0_t (RoundKey[29]), .A0_f (new_AGEMA_signal_5504), .A1_t (new_AGEMA_signal_5505), .A1_f (new_AGEMA_signal_5506), .B0_t (KeyExpansionOutput[61]), .B0_f (new_AGEMA_signal_16511), .B1_t (new_AGEMA_signal_16512), .B1_f (new_AGEMA_signal_16513), .Z0_t (KeyExpansionOutput[29]), .Z0_f (new_AGEMA_signal_17231), .Z1_t (new_AGEMA_signal_17232), .Z1_f (new_AGEMA_signal_17233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U95 ( .A0_t (RoundKey[61]), .A0_f (new_AGEMA_signal_5828), .A1_t (new_AGEMA_signal_5829), .A1_f (new_AGEMA_signal_5830), .B0_t (KeyExpansionOutput[93]), .B0_f (new_AGEMA_signal_15746), .B1_t (new_AGEMA_signal_15747), .B1_f (new_AGEMA_signal_15748), .Z0_t (KeyExpansionOutput[61]), .Z0_f (new_AGEMA_signal_16511), .Z1_t (new_AGEMA_signal_16512), .Z1_f (new_AGEMA_signal_16513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U94 ( .A0_t (RoundKey[93]), .A0_f (new_AGEMA_signal_6143), .A1_t (new_AGEMA_signal_6144), .A1_f (new_AGEMA_signal_6145), .B0_t (KeyExpansionOutput[125]), .B0_f (new_AGEMA_signal_15041), .B1_t (new_AGEMA_signal_15042), .B1_f (new_AGEMA_signal_15043), .Z0_t (KeyExpansionOutput[93]), .Z0_f (new_AGEMA_signal_15746), .Z1_t (new_AGEMA_signal_15747), .Z1_f (new_AGEMA_signal_15748) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U93 ( .A0_t (RoundKey[28]), .A0_f (new_AGEMA_signal_5495), .A1_t (new_AGEMA_signal_5496), .A1_f (new_AGEMA_signal_5497), .B0_t (KeyExpansionOutput[60]), .B0_f (new_AGEMA_signal_16514), .B1_t (new_AGEMA_signal_16515), .B1_f (new_AGEMA_signal_16516), .Z0_t (KeyExpansionOutput[28]), .Z0_f (new_AGEMA_signal_17234), .Z1_t (new_AGEMA_signal_17235), .Z1_f (new_AGEMA_signal_17236) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U92 ( .A0_t (RoundKey[60]), .A0_f (new_AGEMA_signal_5819), .A1_t (new_AGEMA_signal_5820), .A1_f (new_AGEMA_signal_5821), .B0_t (KeyExpansionOutput[92]), .B0_f (new_AGEMA_signal_15749), .B1_t (new_AGEMA_signal_15750), .B1_f (new_AGEMA_signal_15751), .Z0_t (KeyExpansionOutput[60]), .Z0_f (new_AGEMA_signal_16514), .Z1_t (new_AGEMA_signal_16515), .Z1_f (new_AGEMA_signal_16516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U91 ( .A0_t (RoundKey[92]), .A0_f (new_AGEMA_signal_6134), .A1_t (new_AGEMA_signal_6135), .A1_f (new_AGEMA_signal_6136), .B0_t (KeyExpansionOutput[124]), .B0_f (new_AGEMA_signal_15044), .B1_t (new_AGEMA_signal_15045), .B1_f (new_AGEMA_signal_15046), .Z0_t (KeyExpansionOutput[92]), .Z0_f (new_AGEMA_signal_15749), .Z1_t (new_AGEMA_signal_15750), .Z1_f (new_AGEMA_signal_15751) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U90 ( .A0_t (RoundKey[27]), .A0_f (new_AGEMA_signal_5486), .A1_t (new_AGEMA_signal_5487), .A1_f (new_AGEMA_signal_5488), .B0_t (KeyExpansionOutput[59]), .B0_f (new_AGEMA_signal_16517), .B1_t (new_AGEMA_signal_16518), .B1_f (new_AGEMA_signal_16519), .Z0_t (KeyExpansionOutput[27]), .Z0_f (new_AGEMA_signal_17237), .Z1_t (new_AGEMA_signal_17238), .Z1_f (new_AGEMA_signal_17239) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U89 ( .A0_t (RoundKey[59]), .A0_f (new_AGEMA_signal_5801), .A1_t (new_AGEMA_signal_5802), .A1_f (new_AGEMA_signal_5803), .B0_t (KeyExpansionOutput[91]), .B0_f (new_AGEMA_signal_15752), .B1_t (new_AGEMA_signal_15753), .B1_f (new_AGEMA_signal_15754), .Z0_t (KeyExpansionOutput[59]), .Z0_f (new_AGEMA_signal_16517), .Z1_t (new_AGEMA_signal_16518), .Z1_f (new_AGEMA_signal_16519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U88 ( .A0_t (RoundKey[91]), .A0_f (new_AGEMA_signal_6125), .A1_t (new_AGEMA_signal_6126), .A1_f (new_AGEMA_signal_6127), .B0_t (KeyExpansionOutput[123]), .B0_f (new_AGEMA_signal_15047), .B1_t (new_AGEMA_signal_15048), .B1_f (new_AGEMA_signal_15049), .Z0_t (KeyExpansionOutput[91]), .Z0_f (new_AGEMA_signal_15752), .Z1_t (new_AGEMA_signal_15753), .Z1_f (new_AGEMA_signal_15754) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U87 ( .A0_t (RoundKey[26]), .A0_f (new_AGEMA_signal_5477), .A1_t (new_AGEMA_signal_5478), .A1_f (new_AGEMA_signal_5479), .B0_t (KeyExpansionOutput[58]), .B0_f (new_AGEMA_signal_16520), .B1_t (new_AGEMA_signal_16521), .B1_f (new_AGEMA_signal_16522), .Z0_t (KeyExpansionOutput[26]), .Z0_f (new_AGEMA_signal_17240), .Z1_t (new_AGEMA_signal_17241), .Z1_f (new_AGEMA_signal_17242) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U86 ( .A0_t (RoundKey[58]), .A0_f (new_AGEMA_signal_5792), .A1_t (new_AGEMA_signal_5793), .A1_f (new_AGEMA_signal_5794), .B0_t (KeyExpansionOutput[90]), .B0_f (new_AGEMA_signal_15755), .B1_t (new_AGEMA_signal_15756), .B1_f (new_AGEMA_signal_15757), .Z0_t (KeyExpansionOutput[58]), .Z0_f (new_AGEMA_signal_16520), .Z1_t (new_AGEMA_signal_16521), .Z1_f (new_AGEMA_signal_16522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U85 ( .A0_t (RoundKey[90]), .A0_f (new_AGEMA_signal_6116), .A1_t (new_AGEMA_signal_6117), .A1_f (new_AGEMA_signal_6118), .B0_t (KeyExpansionOutput[122]), .B0_f (new_AGEMA_signal_15050), .B1_t (new_AGEMA_signal_15051), .B1_f (new_AGEMA_signal_15052), .Z0_t (KeyExpansionOutput[90]), .Z0_f (new_AGEMA_signal_15755), .Z1_t (new_AGEMA_signal_15756), .Z1_f (new_AGEMA_signal_15757) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U84 ( .A0_t (RoundKey[25]), .A0_f (new_AGEMA_signal_5468), .A1_t (new_AGEMA_signal_5469), .A1_f (new_AGEMA_signal_5470), .B0_t (KeyExpansionOutput[57]), .B0_f (new_AGEMA_signal_16523), .B1_t (new_AGEMA_signal_16524), .B1_f (new_AGEMA_signal_16525), .Z0_t (KeyExpansionOutput[25]), .Z0_f (new_AGEMA_signal_17243), .Z1_t (new_AGEMA_signal_17244), .Z1_f (new_AGEMA_signal_17245) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U83 ( .A0_t (RoundKey[57]), .A0_f (new_AGEMA_signal_5783), .A1_t (new_AGEMA_signal_5784), .A1_f (new_AGEMA_signal_5785), .B0_t (KeyExpansionOutput[89]), .B0_f (new_AGEMA_signal_15758), .B1_t (new_AGEMA_signal_15759), .B1_f (new_AGEMA_signal_15760), .Z0_t (KeyExpansionOutput[57]), .Z0_f (new_AGEMA_signal_16523), .Z1_t (new_AGEMA_signal_16524), .Z1_f (new_AGEMA_signal_16525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U82 ( .A0_t (RoundKey[89]), .A0_f (new_AGEMA_signal_6098), .A1_t (new_AGEMA_signal_6099), .A1_f (new_AGEMA_signal_6100), .B0_t (KeyExpansionOutput[121]), .B0_f (new_AGEMA_signal_15053), .B1_t (new_AGEMA_signal_15054), .B1_f (new_AGEMA_signal_15055), .Z0_t (KeyExpansionOutput[89]), .Z0_f (new_AGEMA_signal_15758), .Z1_t (new_AGEMA_signal_15759), .Z1_f (new_AGEMA_signal_15760) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U81 ( .A0_t (RoundKey[24]), .A0_f (new_AGEMA_signal_5459), .A1_t (new_AGEMA_signal_5460), .A1_f (new_AGEMA_signal_5461), .B0_t (KeyExpansionOutput[56]), .B0_f (new_AGEMA_signal_15761), .B1_t (new_AGEMA_signal_15762), .B1_f (new_AGEMA_signal_15763), .Z0_t (KeyExpansionOutput[24]), .Z0_f (new_AGEMA_signal_16526), .Z1_t (new_AGEMA_signal_16527), .Z1_f (new_AGEMA_signal_16528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U80 ( .A0_t (RoundKey[56]), .A0_f (new_AGEMA_signal_5774), .A1_t (new_AGEMA_signal_5775), .A1_f (new_AGEMA_signal_5776), .B0_t (KeyExpansionOutput[88]), .B0_f (new_AGEMA_signal_14993), .B1_t (new_AGEMA_signal_14994), .B1_f (new_AGEMA_signal_14995), .Z0_t (KeyExpansionOutput[56]), .Z0_f (new_AGEMA_signal_15761), .Z1_t (new_AGEMA_signal_15762), .Z1_f (new_AGEMA_signal_15763) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U79 ( .A0_t (RoundKey[88]), .A0_f (new_AGEMA_signal_6089), .A1_t (new_AGEMA_signal_6090), .A1_f (new_AGEMA_signal_6091), .B0_t (KeyExpansionOutput[120]), .B0_f (new_AGEMA_signal_14009), .B1_t (new_AGEMA_signal_14010), .B1_f (new_AGEMA_signal_14011), .Z0_t (KeyExpansionOutput[88]), .Z0_f (new_AGEMA_signal_14993), .Z1_t (new_AGEMA_signal_14994), .Z1_f (new_AGEMA_signal_14995) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U78 ( .A0_t (RoundKey[23]), .A0_f (new_AGEMA_signal_5450), .A1_t (new_AGEMA_signal_5451), .A1_f (new_AGEMA_signal_5452), .B0_t (KeyExpansionOutput[55]), .B0_f (new_AGEMA_signal_15764), .B1_t (new_AGEMA_signal_15765), .B1_f (new_AGEMA_signal_15766), .Z0_t (KeyExpansionOutput[23]), .Z0_f (new_AGEMA_signal_16529), .Z1_t (new_AGEMA_signal_16530), .Z1_f (new_AGEMA_signal_16531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U77 ( .A0_t (RoundKey[55]), .A0_f (new_AGEMA_signal_5765), .A1_t (new_AGEMA_signal_5766), .A1_f (new_AGEMA_signal_5767), .B0_t (KeyExpansionOutput[87]), .B0_f (new_AGEMA_signal_14996), .B1_t (new_AGEMA_signal_14997), .B1_f (new_AGEMA_signal_14998), .Z0_t (KeyExpansionOutput[55]), .Z0_f (new_AGEMA_signal_15764), .Z1_t (new_AGEMA_signal_15765), .Z1_f (new_AGEMA_signal_15766) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U76 ( .A0_t (RoundKey[87]), .A0_f (new_AGEMA_signal_6080), .A1_t (new_AGEMA_signal_6081), .A1_f (new_AGEMA_signal_6082), .B0_t (KeyExpansionOutput[119]), .B0_f (new_AGEMA_signal_14012), .B1_t (new_AGEMA_signal_14013), .B1_f (new_AGEMA_signal_14014), .Z0_t (KeyExpansionOutput[87]), .Z0_f (new_AGEMA_signal_14996), .Z1_t (new_AGEMA_signal_14997), .Z1_f (new_AGEMA_signal_14998) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U75 ( .A0_t (RoundKey[22]), .A0_f (new_AGEMA_signal_5441), .A1_t (new_AGEMA_signal_5442), .A1_f (new_AGEMA_signal_5443), .B0_t (KeyExpansionOutput[54]), .B0_f (new_AGEMA_signal_15767), .B1_t (new_AGEMA_signal_15768), .B1_f (new_AGEMA_signal_15769), .Z0_t (KeyExpansionOutput[22]), .Z0_f (new_AGEMA_signal_16532), .Z1_t (new_AGEMA_signal_16533), .Z1_f (new_AGEMA_signal_16534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U74 ( .A0_t (RoundKey[54]), .A0_f (new_AGEMA_signal_5756), .A1_t (new_AGEMA_signal_5757), .A1_f (new_AGEMA_signal_5758), .B0_t (KeyExpansionOutput[86]), .B0_f (new_AGEMA_signal_14999), .B1_t (new_AGEMA_signal_15000), .B1_f (new_AGEMA_signal_15001), .Z0_t (KeyExpansionOutput[54]), .Z0_f (new_AGEMA_signal_15767), .Z1_t (new_AGEMA_signal_15768), .Z1_f (new_AGEMA_signal_15769) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U73 ( .A0_t (RoundKey[86]), .A0_f (new_AGEMA_signal_6071), .A1_t (new_AGEMA_signal_6072), .A1_f (new_AGEMA_signal_6073), .B0_t (KeyExpansionOutput[118]), .B0_f (new_AGEMA_signal_14015), .B1_t (new_AGEMA_signal_14016), .B1_f (new_AGEMA_signal_14017), .Z0_t (KeyExpansionOutput[86]), .Z0_f (new_AGEMA_signal_14999), .Z1_t (new_AGEMA_signal_15000), .Z1_f (new_AGEMA_signal_15001) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U72 ( .A0_t (RoundKey[21]), .A0_f (new_AGEMA_signal_5432), .A1_t (new_AGEMA_signal_5433), .A1_f (new_AGEMA_signal_5434), .B0_t (KeyExpansionOutput[53]), .B0_f (new_AGEMA_signal_15770), .B1_t (new_AGEMA_signal_15771), .B1_f (new_AGEMA_signal_15772), .Z0_t (KeyExpansionOutput[21]), .Z0_f (new_AGEMA_signal_16535), .Z1_t (new_AGEMA_signal_16536), .Z1_f (new_AGEMA_signal_16537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U71 ( .A0_t (RoundKey[53]), .A0_f (new_AGEMA_signal_5747), .A1_t (new_AGEMA_signal_5748), .A1_f (new_AGEMA_signal_5749), .B0_t (KeyExpansionOutput[85]), .B0_f (new_AGEMA_signal_15002), .B1_t (new_AGEMA_signal_15003), .B1_f (new_AGEMA_signal_15004), .Z0_t (KeyExpansionOutput[53]), .Z0_f (new_AGEMA_signal_15770), .Z1_t (new_AGEMA_signal_15771), .Z1_f (new_AGEMA_signal_15772) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U70 ( .A0_t (RoundKey[85]), .A0_f (new_AGEMA_signal_6062), .A1_t (new_AGEMA_signal_6063), .A1_f (new_AGEMA_signal_6064), .B0_t (KeyExpansionOutput[117]), .B0_f (new_AGEMA_signal_14018), .B1_t (new_AGEMA_signal_14019), .B1_f (new_AGEMA_signal_14020), .Z0_t (KeyExpansionOutput[85]), .Z0_f (new_AGEMA_signal_15002), .Z1_t (new_AGEMA_signal_15003), .Z1_f (new_AGEMA_signal_15004) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U69 ( .A0_t (RoundKey[20]), .A0_f (new_AGEMA_signal_5423), .A1_t (new_AGEMA_signal_5424), .A1_f (new_AGEMA_signal_5425), .B0_t (KeyExpansionOutput[52]), .B0_f (new_AGEMA_signal_15773), .B1_t (new_AGEMA_signal_15774), .B1_f (new_AGEMA_signal_15775), .Z0_t (KeyExpansionOutput[20]), .Z0_f (new_AGEMA_signal_16538), .Z1_t (new_AGEMA_signal_16539), .Z1_f (new_AGEMA_signal_16540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U68 ( .A0_t (RoundKey[52]), .A0_f (new_AGEMA_signal_5738), .A1_t (new_AGEMA_signal_5739), .A1_f (new_AGEMA_signal_5740), .B0_t (KeyExpansionOutput[84]), .B0_f (new_AGEMA_signal_15005), .B1_t (new_AGEMA_signal_15006), .B1_f (new_AGEMA_signal_15007), .Z0_t (KeyExpansionOutput[52]), .Z0_f (new_AGEMA_signal_15773), .Z1_t (new_AGEMA_signal_15774), .Z1_f (new_AGEMA_signal_15775) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U67 ( .A0_t (RoundKey[84]), .A0_f (new_AGEMA_signal_6053), .A1_t (new_AGEMA_signal_6054), .A1_f (new_AGEMA_signal_6055), .B0_t (KeyExpansionOutput[116]), .B0_f (new_AGEMA_signal_14021), .B1_t (new_AGEMA_signal_14022), .B1_f (new_AGEMA_signal_14023), .Z0_t (KeyExpansionOutput[84]), .Z0_f (new_AGEMA_signal_15005), .Z1_t (new_AGEMA_signal_15006), .Z1_f (new_AGEMA_signal_15007) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U66 ( .A0_t (RoundKey[1]), .A0_f (new_AGEMA_signal_5414), .A1_t (new_AGEMA_signal_5415), .A1_f (new_AGEMA_signal_5416), .B0_t (KeyExpansionOutput[33]), .B0_f (new_AGEMA_signal_15776), .B1_t (new_AGEMA_signal_15777), .B1_f (new_AGEMA_signal_15778), .Z0_t (KeyExpansionOutput[1]), .Z0_f (new_AGEMA_signal_16541), .Z1_t (new_AGEMA_signal_16542), .Z1_f (new_AGEMA_signal_16543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U65 ( .A0_t (RoundKey[33]), .A0_f (new_AGEMA_signal_5549), .A1_t (new_AGEMA_signal_5550), .A1_f (new_AGEMA_signal_5551), .B0_t (KeyExpansionOutput[65]), .B0_f (new_AGEMA_signal_15008), .B1_t (new_AGEMA_signal_15009), .B1_f (new_AGEMA_signal_15010), .Z0_t (KeyExpansionOutput[33]), .Z0_f (new_AGEMA_signal_15776), .Z1_t (new_AGEMA_signal_15777), .Z1_f (new_AGEMA_signal_15778) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U64 ( .A0_t (RoundKey[65]), .A0_f (new_AGEMA_signal_5864), .A1_t (new_AGEMA_signal_5865), .A1_f (new_AGEMA_signal_5866), .B0_t (KeyExpansionOutput[97]), .B0_f (new_AGEMA_signal_14003), .B1_t (new_AGEMA_signal_14004), .B1_f (new_AGEMA_signal_14005), .Z0_t (KeyExpansionOutput[65]), .Z0_f (new_AGEMA_signal_15008), .Z1_t (new_AGEMA_signal_15009), .Z1_f (new_AGEMA_signal_15010) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U63 ( .A0_t (RoundKey[97]), .A0_f (new_AGEMA_signal_6179), .A1_t (new_AGEMA_signal_6180), .A1_f (new_AGEMA_signal_6181), .B0_t (KeyExpansionIns_tmp[1]), .B0_f (new_AGEMA_signal_13589), .B1_t (new_AGEMA_signal_13590), .B1_f (new_AGEMA_signal_13591), .Z0_t (KeyExpansionOutput[97]), .Z0_f (new_AGEMA_signal_14003), .Z1_t (new_AGEMA_signal_14004), .Z1_f (new_AGEMA_signal_14005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U62 ( .A0_t (RoundKey[19]), .A0_f (new_AGEMA_signal_5405), .A1_t (new_AGEMA_signal_5406), .A1_f (new_AGEMA_signal_5407), .B0_t (KeyExpansionOutput[51]), .B0_f (new_AGEMA_signal_15779), .B1_t (new_AGEMA_signal_15780), .B1_f (new_AGEMA_signal_15781), .Z0_t (KeyExpansionOutput[19]), .Z0_f (new_AGEMA_signal_16544), .Z1_t (new_AGEMA_signal_16545), .Z1_f (new_AGEMA_signal_16546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U61 ( .A0_t (RoundKey[51]), .A0_f (new_AGEMA_signal_5729), .A1_t (new_AGEMA_signal_5730), .A1_f (new_AGEMA_signal_5731), .B0_t (KeyExpansionOutput[83]), .B0_f (new_AGEMA_signal_15011), .B1_t (new_AGEMA_signal_15012), .B1_f (new_AGEMA_signal_15013), .Z0_t (KeyExpansionOutput[51]), .Z0_f (new_AGEMA_signal_15779), .Z1_t (new_AGEMA_signal_15780), .Z1_f (new_AGEMA_signal_15781) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U60 ( .A0_t (RoundKey[83]), .A0_f (new_AGEMA_signal_6044), .A1_t (new_AGEMA_signal_6045), .A1_f (new_AGEMA_signal_6046), .B0_t (KeyExpansionOutput[115]), .B0_f (new_AGEMA_signal_14024), .B1_t (new_AGEMA_signal_14025), .B1_f (new_AGEMA_signal_14026), .Z0_t (KeyExpansionOutput[83]), .Z0_f (new_AGEMA_signal_15011), .Z1_t (new_AGEMA_signal_15012), .Z1_f (new_AGEMA_signal_15013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U59 ( .A0_t (RoundKey[18]), .A0_f (new_AGEMA_signal_5396), .A1_t (new_AGEMA_signal_5397), .A1_f (new_AGEMA_signal_5398), .B0_t (KeyExpansionOutput[50]), .B0_f (new_AGEMA_signal_15782), .B1_t (new_AGEMA_signal_15783), .B1_f (new_AGEMA_signal_15784), .Z0_t (KeyExpansionOutput[18]), .Z0_f (new_AGEMA_signal_16547), .Z1_t (new_AGEMA_signal_16548), .Z1_f (new_AGEMA_signal_16549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U58 ( .A0_t (RoundKey[50]), .A0_f (new_AGEMA_signal_5720), .A1_t (new_AGEMA_signal_5721), .A1_f (new_AGEMA_signal_5722), .B0_t (KeyExpansionOutput[82]), .B0_f (new_AGEMA_signal_15014), .B1_t (new_AGEMA_signal_15015), .B1_f (new_AGEMA_signal_15016), .Z0_t (KeyExpansionOutput[50]), .Z0_f (new_AGEMA_signal_15782), .Z1_t (new_AGEMA_signal_15783), .Z1_f (new_AGEMA_signal_15784) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U57 ( .A0_t (RoundKey[82]), .A0_f (new_AGEMA_signal_6035), .A1_t (new_AGEMA_signal_6036), .A1_f (new_AGEMA_signal_6037), .B0_t (KeyExpansionOutput[114]), .B0_f (new_AGEMA_signal_14027), .B1_t (new_AGEMA_signal_14028), .B1_f (new_AGEMA_signal_14029), .Z0_t (KeyExpansionOutput[82]), .Z0_f (new_AGEMA_signal_15014), .Z1_t (new_AGEMA_signal_15015), .Z1_f (new_AGEMA_signal_15016) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U56 ( .A0_t (RoundKey[17]), .A0_f (new_AGEMA_signal_5387), .A1_t (new_AGEMA_signal_5388), .A1_f (new_AGEMA_signal_5389), .B0_t (KeyExpansionOutput[49]), .B0_f (new_AGEMA_signal_15785), .B1_t (new_AGEMA_signal_15786), .B1_f (new_AGEMA_signal_15787), .Z0_t (KeyExpansionOutput[17]), .Z0_f (new_AGEMA_signal_16550), .Z1_t (new_AGEMA_signal_16551), .Z1_f (new_AGEMA_signal_16552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U55 ( .A0_t (RoundKey[49]), .A0_f (new_AGEMA_signal_5702), .A1_t (new_AGEMA_signal_5703), .A1_f (new_AGEMA_signal_5704), .B0_t (KeyExpansionOutput[81]), .B0_f (new_AGEMA_signal_15017), .B1_t (new_AGEMA_signal_15018), .B1_f (new_AGEMA_signal_15019), .Z0_t (KeyExpansionOutput[49]), .Z0_f (new_AGEMA_signal_15785), .Z1_t (new_AGEMA_signal_15786), .Z1_f (new_AGEMA_signal_15787) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U54 ( .A0_t (RoundKey[81]), .A0_f (new_AGEMA_signal_6026), .A1_t (new_AGEMA_signal_6027), .A1_f (new_AGEMA_signal_6028), .B0_t (KeyExpansionOutput[113]), .B0_f (new_AGEMA_signal_14030), .B1_t (new_AGEMA_signal_14031), .B1_f (new_AGEMA_signal_14032), .Z0_t (KeyExpansionOutput[81]), .Z0_f (new_AGEMA_signal_15017), .Z1_t (new_AGEMA_signal_15018), .Z1_f (new_AGEMA_signal_15019) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U53 ( .A0_t (RoundKey[16]), .A0_f (new_AGEMA_signal_5378), .A1_t (new_AGEMA_signal_5379), .A1_f (new_AGEMA_signal_5380), .B0_t (KeyExpansionOutput[48]), .B0_f (new_AGEMA_signal_15020), .B1_t (new_AGEMA_signal_15021), .B1_f (new_AGEMA_signal_15022), .Z0_t (KeyExpansionOutput[16]), .Z0_f (new_AGEMA_signal_15788), .Z1_t (new_AGEMA_signal_15789), .Z1_f (new_AGEMA_signal_15790) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U52 ( .A0_t (RoundKey[48]), .A0_f (new_AGEMA_signal_5693), .A1_t (new_AGEMA_signal_5694), .A1_f (new_AGEMA_signal_5695), .B0_t (KeyExpansionOutput[80]), .B0_f (new_AGEMA_signal_14006), .B1_t (new_AGEMA_signal_14007), .B1_f (new_AGEMA_signal_14008), .Z0_t (KeyExpansionOutput[48]), .Z0_f (new_AGEMA_signal_15020), .Z1_t (new_AGEMA_signal_15021), .Z1_f (new_AGEMA_signal_15022) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U51 ( .A0_t (RoundKey[80]), .A0_f (new_AGEMA_signal_6017), .A1_t (new_AGEMA_signal_6018), .A1_f (new_AGEMA_signal_6019), .B0_t (KeyExpansionOutput[112]), .B0_f (new_AGEMA_signal_13496), .B1_t (new_AGEMA_signal_13497), .B1_f (new_AGEMA_signal_13498), .Z0_t (KeyExpansionOutput[80]), .Z0_f (new_AGEMA_signal_14006), .Z1_t (new_AGEMA_signal_14007), .Z1_f (new_AGEMA_signal_14008) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U50 ( .A0_t (RoundKey[15]), .A0_f (new_AGEMA_signal_5369), .A1_t (new_AGEMA_signal_5370), .A1_f (new_AGEMA_signal_5371), .B0_t (KeyExpansionOutput[47]), .B0_f (new_AGEMA_signal_15791), .B1_t (new_AGEMA_signal_15792), .B1_f (new_AGEMA_signal_15793), .Z0_t (KeyExpansionOutput[15]), .Z0_f (new_AGEMA_signal_16553), .Z1_t (new_AGEMA_signal_16554), .Z1_f (new_AGEMA_signal_16555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U49 ( .A0_t (RoundKey[47]), .A0_f (new_AGEMA_signal_5684), .A1_t (new_AGEMA_signal_5685), .A1_f (new_AGEMA_signal_5686), .B0_t (KeyExpansionOutput[79]), .B0_f (new_AGEMA_signal_15023), .B1_t (new_AGEMA_signal_15024), .B1_f (new_AGEMA_signal_15025), .Z0_t (KeyExpansionOutput[47]), .Z0_f (new_AGEMA_signal_15791), .Z1_t (new_AGEMA_signal_15792), .Z1_f (new_AGEMA_signal_15793) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U48 ( .A0_t (RoundKey[79]), .A0_f (new_AGEMA_signal_5999), .A1_t (new_AGEMA_signal_6000), .A1_f (new_AGEMA_signal_6001), .B0_t (KeyExpansionOutput[111]), .B0_f (new_AGEMA_signal_14033), .B1_t (new_AGEMA_signal_14034), .B1_f (new_AGEMA_signal_14035), .Z0_t (KeyExpansionOutput[79]), .Z0_f (new_AGEMA_signal_15023), .Z1_t (new_AGEMA_signal_15024), .Z1_f (new_AGEMA_signal_15025) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U47 ( .A0_t (RoundKey[14]), .A0_f (new_AGEMA_signal_5360), .A1_t (new_AGEMA_signal_5361), .A1_f (new_AGEMA_signal_5362), .B0_t (KeyExpansionOutput[46]), .B0_f (new_AGEMA_signal_15794), .B1_t (new_AGEMA_signal_15795), .B1_f (new_AGEMA_signal_15796), .Z0_t (KeyExpansionOutput[14]), .Z0_f (new_AGEMA_signal_16556), .Z1_t (new_AGEMA_signal_16557), .Z1_f (new_AGEMA_signal_16558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U46 ( .A0_t (RoundKey[46]), .A0_f (new_AGEMA_signal_5675), .A1_t (new_AGEMA_signal_5676), .A1_f (new_AGEMA_signal_5677), .B0_t (KeyExpansionOutput[78]), .B0_f (new_AGEMA_signal_15026), .B1_t (new_AGEMA_signal_15027), .B1_f (new_AGEMA_signal_15028), .Z0_t (KeyExpansionOutput[46]), .Z0_f (new_AGEMA_signal_15794), .Z1_t (new_AGEMA_signal_15795), .Z1_f (new_AGEMA_signal_15796) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U45 ( .A0_t (RoundKey[78]), .A0_f (new_AGEMA_signal_5990), .A1_t (new_AGEMA_signal_5991), .A1_f (new_AGEMA_signal_5992), .B0_t (KeyExpansionOutput[110]), .B0_f (new_AGEMA_signal_14036), .B1_t (new_AGEMA_signal_14037), .B1_f (new_AGEMA_signal_14038), .Z0_t (KeyExpansionOutput[78]), .Z0_f (new_AGEMA_signal_15026), .Z1_t (new_AGEMA_signal_15027), .Z1_f (new_AGEMA_signal_15028) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U44 ( .A0_t (RoundKey[13]), .A0_f (new_AGEMA_signal_5351), .A1_t (new_AGEMA_signal_5352), .A1_f (new_AGEMA_signal_5353), .B0_t (KeyExpansionOutput[45]), .B0_f (new_AGEMA_signal_15797), .B1_t (new_AGEMA_signal_15798), .B1_f (new_AGEMA_signal_15799), .Z0_t (KeyExpansionOutput[13]), .Z0_f (new_AGEMA_signal_16559), .Z1_t (new_AGEMA_signal_16560), .Z1_f (new_AGEMA_signal_16561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U43 ( .A0_t (RoundKey[45]), .A0_f (new_AGEMA_signal_5666), .A1_t (new_AGEMA_signal_5667), .A1_f (new_AGEMA_signal_5668), .B0_t (KeyExpansionOutput[77]), .B0_f (new_AGEMA_signal_15029), .B1_t (new_AGEMA_signal_15030), .B1_f (new_AGEMA_signal_15031), .Z0_t (KeyExpansionOutput[45]), .Z0_f (new_AGEMA_signal_15797), .Z1_t (new_AGEMA_signal_15798), .Z1_f (new_AGEMA_signal_15799) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U42 ( .A0_t (RoundKey[77]), .A0_f (new_AGEMA_signal_5981), .A1_t (new_AGEMA_signal_5982), .A1_f (new_AGEMA_signal_5983), .B0_t (KeyExpansionOutput[109]), .B0_f (new_AGEMA_signal_14039), .B1_t (new_AGEMA_signal_14040), .B1_f (new_AGEMA_signal_14041), .Z0_t (KeyExpansionOutput[77]), .Z0_f (new_AGEMA_signal_15029), .Z1_t (new_AGEMA_signal_15030), .Z1_f (new_AGEMA_signal_15031) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U41 ( .A0_t (RoundKey[12]), .A0_f (new_AGEMA_signal_5342), .A1_t (new_AGEMA_signal_5343), .A1_f (new_AGEMA_signal_5344), .B0_t (KeyExpansionOutput[44]), .B0_f (new_AGEMA_signal_15800), .B1_t (new_AGEMA_signal_15801), .B1_f (new_AGEMA_signal_15802), .Z0_t (KeyExpansionOutput[12]), .Z0_f (new_AGEMA_signal_16562), .Z1_t (new_AGEMA_signal_16563), .Z1_f (new_AGEMA_signal_16564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U40 ( .A0_t (RoundKey[44]), .A0_f (new_AGEMA_signal_5657), .A1_t (new_AGEMA_signal_5658), .A1_f (new_AGEMA_signal_5659), .B0_t (KeyExpansionOutput[76]), .B0_f (new_AGEMA_signal_15032), .B1_t (new_AGEMA_signal_15033), .B1_f (new_AGEMA_signal_15034), .Z0_t (KeyExpansionOutput[44]), .Z0_f (new_AGEMA_signal_15800), .Z1_t (new_AGEMA_signal_15801), .Z1_f (new_AGEMA_signal_15802) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U39 ( .A0_t (RoundKey[76]), .A0_f (new_AGEMA_signal_5972), .A1_t (new_AGEMA_signal_5973), .A1_f (new_AGEMA_signal_5974), .B0_t (KeyExpansionOutput[108]), .B0_f (new_AGEMA_signal_14042), .B1_t (new_AGEMA_signal_14043), .B1_f (new_AGEMA_signal_14044), .Z0_t (KeyExpansionOutput[76]), .Z0_f (new_AGEMA_signal_15032), .Z1_t (new_AGEMA_signal_15033), .Z1_f (new_AGEMA_signal_15034) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U38 ( .A0_t (RoundKey[127]), .A0_f (new_AGEMA_signal_5333), .A1_t (new_AGEMA_signal_5334), .A1_f (new_AGEMA_signal_5335), .B0_t (KeyExpansionIns_tmp[31]), .B0_f (new_AGEMA_signal_14069), .B1_t (new_AGEMA_signal_14070), .B1_f (new_AGEMA_signal_14071), .Z0_t (KeyExpansionOutput[127]), .Z0_f (new_AGEMA_signal_15035), .Z1_t (new_AGEMA_signal_15036), .Z1_f (new_AGEMA_signal_15037) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U37 ( .A0_t (RoundKey[126]), .A0_f (new_AGEMA_signal_5324), .A1_t (new_AGEMA_signal_5325), .A1_f (new_AGEMA_signal_5326), .B0_t (KeyExpansionIns_tmp[30]), .B0_f (new_AGEMA_signal_14072), .B1_t (new_AGEMA_signal_14073), .B1_f (new_AGEMA_signal_14074), .Z0_t (KeyExpansionOutput[126]), .Z0_f (new_AGEMA_signal_15038), .Z1_t (new_AGEMA_signal_15039), .Z1_f (new_AGEMA_signal_15040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U36 ( .A0_t (RoundKey[125]), .A0_f (new_AGEMA_signal_5315), .A1_t (new_AGEMA_signal_5316), .A1_f (new_AGEMA_signal_5317), .B0_t (KeyExpansionIns_tmp[29]), .B0_f (new_AGEMA_signal_14075), .B1_t (new_AGEMA_signal_14076), .B1_f (new_AGEMA_signal_14077), .Z0_t (KeyExpansionOutput[125]), .Z0_f (new_AGEMA_signal_15041), .Z1_t (new_AGEMA_signal_15042), .Z1_f (new_AGEMA_signal_15043) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U35 ( .A0_t (RoundKey[124]), .A0_f (new_AGEMA_signal_5306), .A1_t (new_AGEMA_signal_5307), .A1_f (new_AGEMA_signal_5308), .B0_t (KeyExpansionIns_tmp[28]), .B0_f (new_AGEMA_signal_14078), .B1_t (new_AGEMA_signal_14079), .B1_f (new_AGEMA_signal_14080), .Z0_t (KeyExpansionOutput[124]), .Z0_f (new_AGEMA_signal_15044), .Z1_t (new_AGEMA_signal_15045), .Z1_f (new_AGEMA_signal_15046) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U34 ( .A0_t (RoundKey[123]), .A0_f (new_AGEMA_signal_5297), .A1_t (new_AGEMA_signal_5298), .A1_f (new_AGEMA_signal_5299), .B0_t (KeyExpansionIns_tmp[27]), .B0_f (new_AGEMA_signal_14081), .B1_t (new_AGEMA_signal_14082), .B1_f (new_AGEMA_signal_14083), .Z0_t (KeyExpansionOutput[123]), .Z0_f (new_AGEMA_signal_15047), .Z1_t (new_AGEMA_signal_15048), .Z1_f (new_AGEMA_signal_15049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U33 ( .A0_t (RoundKey[122]), .A0_f (new_AGEMA_signal_5288), .A1_t (new_AGEMA_signal_5289), .A1_f (new_AGEMA_signal_5290), .B0_t (KeyExpansionIns_tmp[26]), .B0_f (new_AGEMA_signal_14084), .B1_t (new_AGEMA_signal_14085), .B1_f (new_AGEMA_signal_14086), .Z0_t (KeyExpansionOutput[122]), .Z0_f (new_AGEMA_signal_15050), .Z1_t (new_AGEMA_signal_15051), .Z1_f (new_AGEMA_signal_15052) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U32 ( .A0_t (RoundKey[121]), .A0_f (new_AGEMA_signal_5279), .A1_t (new_AGEMA_signal_5280), .A1_f (new_AGEMA_signal_5281), .B0_t (KeyExpansionIns_tmp[25]), .B0_f (new_AGEMA_signal_14087), .B1_t (new_AGEMA_signal_14088), .B1_f (new_AGEMA_signal_14089), .Z0_t (KeyExpansionOutput[121]), .Z0_f (new_AGEMA_signal_15053), .Z1_t (new_AGEMA_signal_15054), .Z1_f (new_AGEMA_signal_15055) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U31 ( .A0_t (RoundKey[120]), .A0_f (new_AGEMA_signal_5270), .A1_t (new_AGEMA_signal_5271), .A1_f (new_AGEMA_signal_5272), .B0_t (KeyExpansionIns_tmp[24]), .B0_f (new_AGEMA_signal_13505), .B1_t (new_AGEMA_signal_13506), .B1_f (new_AGEMA_signal_13507), .Z0_t (KeyExpansionOutput[120]), .Z0_f (new_AGEMA_signal_14009), .Z1_t (new_AGEMA_signal_14010), .Z1_f (new_AGEMA_signal_14011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U30 ( .A0_t (RoundKey[11]), .A0_f (new_AGEMA_signal_5261), .A1_t (new_AGEMA_signal_5262), .A1_f (new_AGEMA_signal_5263), .B0_t (KeyExpansionOutput[43]), .B0_f (new_AGEMA_signal_15803), .B1_t (new_AGEMA_signal_15804), .B1_f (new_AGEMA_signal_15805), .Z0_t (KeyExpansionOutput[11]), .Z0_f (new_AGEMA_signal_16565), .Z1_t (new_AGEMA_signal_16566), .Z1_f (new_AGEMA_signal_16567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U29 ( .A0_t (RoundKey[43]), .A0_f (new_AGEMA_signal_5648), .A1_t (new_AGEMA_signal_5649), .A1_f (new_AGEMA_signal_5650), .B0_t (KeyExpansionOutput[75]), .B0_f (new_AGEMA_signal_15056), .B1_t (new_AGEMA_signal_15057), .B1_f (new_AGEMA_signal_15058), .Z0_t (KeyExpansionOutput[43]), .Z0_f (new_AGEMA_signal_15803), .Z1_t (new_AGEMA_signal_15804), .Z1_f (new_AGEMA_signal_15805) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U28 ( .A0_t (RoundKey[75]), .A0_f (new_AGEMA_signal_5963), .A1_t (new_AGEMA_signal_5964), .A1_f (new_AGEMA_signal_5965), .B0_t (KeyExpansionOutput[107]), .B0_f (new_AGEMA_signal_14045), .B1_t (new_AGEMA_signal_14046), .B1_f (new_AGEMA_signal_14047), .Z0_t (KeyExpansionOutput[75]), .Z0_f (new_AGEMA_signal_15056), .Z1_t (new_AGEMA_signal_15057), .Z1_f (new_AGEMA_signal_15058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U27 ( .A0_t (RoundKey[119]), .A0_f (new_AGEMA_signal_5252), .A1_t (new_AGEMA_signal_5253), .A1_f (new_AGEMA_signal_5254), .B0_t (KeyExpansionIns_tmp[23]), .B0_f (new_AGEMA_signal_13529), .B1_t (new_AGEMA_signal_13530), .B1_f (new_AGEMA_signal_13531), .Z0_t (KeyExpansionOutput[119]), .Z0_f (new_AGEMA_signal_14012), .Z1_t (new_AGEMA_signal_14013), .Z1_f (new_AGEMA_signal_14014) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U26 ( .A0_t (RoundKey[118]), .A0_f (new_AGEMA_signal_5243), .A1_t (new_AGEMA_signal_5244), .A1_f (new_AGEMA_signal_5245), .B0_t (KeyExpansionIns_tmp[22]), .B0_f (new_AGEMA_signal_13532), .B1_t (new_AGEMA_signal_13533), .B1_f (new_AGEMA_signal_13534), .Z0_t (KeyExpansionOutput[118]), .Z0_f (new_AGEMA_signal_14015), .Z1_t (new_AGEMA_signal_14016), .Z1_f (new_AGEMA_signal_14017) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U25 ( .A0_t (RoundKey[117]), .A0_f (new_AGEMA_signal_5234), .A1_t (new_AGEMA_signal_5235), .A1_f (new_AGEMA_signal_5236), .B0_t (KeyExpansionIns_tmp[21]), .B0_f (new_AGEMA_signal_13535), .B1_t (new_AGEMA_signal_13536), .B1_f (new_AGEMA_signal_13537), .Z0_t (KeyExpansionOutput[117]), .Z0_f (new_AGEMA_signal_14018), .Z1_t (new_AGEMA_signal_14019), .Z1_f (new_AGEMA_signal_14020) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U24 ( .A0_t (RoundKey[116]), .A0_f (new_AGEMA_signal_5225), .A1_t (new_AGEMA_signal_5226), .A1_f (new_AGEMA_signal_5227), .B0_t (KeyExpansionIns_tmp[20]), .B0_f (new_AGEMA_signal_13538), .B1_t (new_AGEMA_signal_13539), .B1_f (new_AGEMA_signal_13540), .Z0_t (KeyExpansionOutput[116]), .Z0_f (new_AGEMA_signal_14021), .Z1_t (new_AGEMA_signal_14022), .Z1_f (new_AGEMA_signal_14023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U23 ( .A0_t (RoundKey[115]), .A0_f (new_AGEMA_signal_5216), .A1_t (new_AGEMA_signal_5217), .A1_f (new_AGEMA_signal_5218), .B0_t (KeyExpansionIns_tmp[19]), .B0_f (new_AGEMA_signal_13541), .B1_t (new_AGEMA_signal_13542), .B1_f (new_AGEMA_signal_13543), .Z0_t (KeyExpansionOutput[115]), .Z0_f (new_AGEMA_signal_14024), .Z1_t (new_AGEMA_signal_14025), .Z1_f (new_AGEMA_signal_14026) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U22 ( .A0_t (RoundKey[114]), .A0_f (new_AGEMA_signal_5207), .A1_t (new_AGEMA_signal_5208), .A1_f (new_AGEMA_signal_5209), .B0_t (KeyExpansionIns_tmp[18]), .B0_f (new_AGEMA_signal_13544), .B1_t (new_AGEMA_signal_13545), .B1_f (new_AGEMA_signal_13546), .Z0_t (KeyExpansionOutput[114]), .Z0_f (new_AGEMA_signal_14027), .Z1_t (new_AGEMA_signal_14028), .Z1_f (new_AGEMA_signal_14029) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U21 ( .A0_t (RoundKey[113]), .A0_f (new_AGEMA_signal_5198), .A1_t (new_AGEMA_signal_5199), .A1_f (new_AGEMA_signal_5200), .B0_t (KeyExpansionIns_tmp[17]), .B0_f (new_AGEMA_signal_13547), .B1_t (new_AGEMA_signal_13548), .B1_f (new_AGEMA_signal_13549), .Z0_t (KeyExpansionOutput[113]), .Z0_f (new_AGEMA_signal_14030), .Z1_t (new_AGEMA_signal_14031), .Z1_f (new_AGEMA_signal_14032) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U20 ( .A0_t (RoundKey[112]), .A0_f (new_AGEMA_signal_5189), .A1_t (new_AGEMA_signal_5190), .A1_f (new_AGEMA_signal_5191), .B0_t (KeyExpansionIns_tmp[16]), .B0_f (new_AGEMA_signal_12899), .B1_t (new_AGEMA_signal_12900), .B1_f (new_AGEMA_signal_12901), .Z0_t (KeyExpansionOutput[112]), .Z0_f (new_AGEMA_signal_13496), .Z1_t (new_AGEMA_signal_13497), .Z1_f (new_AGEMA_signal_13498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U19 ( .A0_t (RoundKey[111]), .A0_f (new_AGEMA_signal_5180), .A1_t (new_AGEMA_signal_5181), .A1_f (new_AGEMA_signal_5182), .B0_t (KeyExpansionIns_tmp[15]), .B0_f (new_AGEMA_signal_13550), .B1_t (new_AGEMA_signal_13551), .B1_f (new_AGEMA_signal_13552), .Z0_t (KeyExpansionOutput[111]), .Z0_f (new_AGEMA_signal_14033), .Z1_t (new_AGEMA_signal_14034), .Z1_f (new_AGEMA_signal_14035) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U18 ( .A0_t (RoundKey[110]), .A0_f (new_AGEMA_signal_5171), .A1_t (new_AGEMA_signal_5172), .A1_f (new_AGEMA_signal_5173), .B0_t (KeyExpansionIns_tmp[14]), .B0_f (new_AGEMA_signal_13553), .B1_t (new_AGEMA_signal_13554), .B1_f (new_AGEMA_signal_13555), .Z0_t (KeyExpansionOutput[110]), .Z0_f (new_AGEMA_signal_14036), .Z1_t (new_AGEMA_signal_14037), .Z1_f (new_AGEMA_signal_14038) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U17 ( .A0_t (RoundKey[10]), .A0_f (new_AGEMA_signal_5162), .A1_t (new_AGEMA_signal_5163), .A1_f (new_AGEMA_signal_5164), .B0_t (KeyExpansionOutput[42]), .B0_f (new_AGEMA_signal_15806), .B1_t (new_AGEMA_signal_15807), .B1_f (new_AGEMA_signal_15808), .Z0_t (KeyExpansionOutput[10]), .Z0_f (new_AGEMA_signal_16568), .Z1_t (new_AGEMA_signal_16569), .Z1_f (new_AGEMA_signal_16570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U16 ( .A0_t (RoundKey[42]), .A0_f (new_AGEMA_signal_5639), .A1_t (new_AGEMA_signal_5640), .A1_f (new_AGEMA_signal_5641), .B0_t (KeyExpansionOutput[74]), .B0_f (new_AGEMA_signal_15059), .B1_t (new_AGEMA_signal_15060), .B1_f (new_AGEMA_signal_15061), .Z0_t (KeyExpansionOutput[42]), .Z0_f (new_AGEMA_signal_15806), .Z1_t (new_AGEMA_signal_15807), .Z1_f (new_AGEMA_signal_15808) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U15 ( .A0_t (RoundKey[74]), .A0_f (new_AGEMA_signal_5954), .A1_t (new_AGEMA_signal_5955), .A1_f (new_AGEMA_signal_5956), .B0_t (KeyExpansionOutput[106]), .B0_f (new_AGEMA_signal_14048), .B1_t (new_AGEMA_signal_14049), .B1_f (new_AGEMA_signal_14050), .Z0_t (KeyExpansionOutput[74]), .Z0_f (new_AGEMA_signal_15059), .Z1_t (new_AGEMA_signal_15060), .Z1_f (new_AGEMA_signal_15061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U14 ( .A0_t (RoundKey[109]), .A0_f (new_AGEMA_signal_5153), .A1_t (new_AGEMA_signal_5154), .A1_f (new_AGEMA_signal_5155), .B0_t (KeyExpansionIns_tmp[13]), .B0_f (new_AGEMA_signal_13556), .B1_t (new_AGEMA_signal_13557), .B1_f (new_AGEMA_signal_13558), .Z0_t (KeyExpansionOutput[109]), .Z0_f (new_AGEMA_signal_14039), .Z1_t (new_AGEMA_signal_14040), .Z1_f (new_AGEMA_signal_14041) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U13 ( .A0_t (RoundKey[108]), .A0_f (new_AGEMA_signal_5144), .A1_t (new_AGEMA_signal_5145), .A1_f (new_AGEMA_signal_5146), .B0_t (KeyExpansionIns_tmp[12]), .B0_f (new_AGEMA_signal_13559), .B1_t (new_AGEMA_signal_13560), .B1_f (new_AGEMA_signal_13561), .Z0_t (KeyExpansionOutput[108]), .Z0_f (new_AGEMA_signal_14042), .Z1_t (new_AGEMA_signal_14043), .Z1_f (new_AGEMA_signal_14044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U12 ( .A0_t (RoundKey[107]), .A0_f (new_AGEMA_signal_5135), .A1_t (new_AGEMA_signal_5136), .A1_f (new_AGEMA_signal_5137), .B0_t (KeyExpansionIns_tmp[11]), .B0_f (new_AGEMA_signal_13562), .B1_t (new_AGEMA_signal_13563), .B1_f (new_AGEMA_signal_13564), .Z0_t (KeyExpansionOutput[107]), .Z0_f (new_AGEMA_signal_14045), .Z1_t (new_AGEMA_signal_14046), .Z1_f (new_AGEMA_signal_14047) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U11 ( .A0_t (RoundKey[106]), .A0_f (new_AGEMA_signal_5126), .A1_t (new_AGEMA_signal_5127), .A1_f (new_AGEMA_signal_5128), .B0_t (KeyExpansionIns_tmp[10]), .B0_f (new_AGEMA_signal_13565), .B1_t (new_AGEMA_signal_13566), .B1_f (new_AGEMA_signal_13567), .Z0_t (KeyExpansionOutput[106]), .Z0_f (new_AGEMA_signal_14048), .Z1_t (new_AGEMA_signal_14049), .Z1_f (new_AGEMA_signal_14050) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U10 ( .A0_t (RoundKey[105]), .A0_f (new_AGEMA_signal_5117), .A1_t (new_AGEMA_signal_5118), .A1_f (new_AGEMA_signal_5119), .B0_t (KeyExpansionIns_tmp[9]), .B0_f (new_AGEMA_signal_13568), .B1_t (new_AGEMA_signal_13569), .B1_f (new_AGEMA_signal_13570), .Z0_t (KeyExpansionOutput[105]), .Z0_f (new_AGEMA_signal_14051), .Z1_t (new_AGEMA_signal_14052), .Z1_f (new_AGEMA_signal_14053) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U9 ( .A0_t (RoundKey[104]), .A0_f (new_AGEMA_signal_5108), .A1_t (new_AGEMA_signal_5109), .A1_f (new_AGEMA_signal_5110), .B0_t (KeyExpansionIns_tmp[8]), .B0_f (new_AGEMA_signal_12932), .B1_t (new_AGEMA_signal_12933), .B1_f (new_AGEMA_signal_12934), .Z0_t (KeyExpansionOutput[104]), .Z0_f (new_AGEMA_signal_13499), .Z1_t (new_AGEMA_signal_13500), .Z1_f (new_AGEMA_signal_13501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U8 ( .A0_t (RoundKey[103]), .A0_f (new_AGEMA_signal_5099), .A1_t (new_AGEMA_signal_5100), .A1_f (new_AGEMA_signal_5101), .B0_t (KeyExpansionIns_tmp[7]), .B0_f (new_AGEMA_signal_13571), .B1_t (new_AGEMA_signal_13572), .B1_f (new_AGEMA_signal_13573), .Z0_t (KeyExpansionOutput[103]), .Z0_f (new_AGEMA_signal_14054), .Z1_t (new_AGEMA_signal_14055), .Z1_f (new_AGEMA_signal_14056) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U7 ( .A0_t (RoundKey[102]), .A0_f (new_AGEMA_signal_5090), .A1_t (new_AGEMA_signal_5091), .A1_f (new_AGEMA_signal_5092), .B0_t (KeyExpansionIns_tmp[6]), .B0_f (new_AGEMA_signal_13574), .B1_t (new_AGEMA_signal_13575), .B1_f (new_AGEMA_signal_13576), .Z0_t (KeyExpansionOutput[102]), .Z0_f (new_AGEMA_signal_14057), .Z1_t (new_AGEMA_signal_14058), .Z1_f (new_AGEMA_signal_14059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U6 ( .A0_t (RoundKey[101]), .A0_f (new_AGEMA_signal_5081), .A1_t (new_AGEMA_signal_5082), .A1_f (new_AGEMA_signal_5083), .B0_t (KeyExpansionIns_tmp[5]), .B0_f (new_AGEMA_signal_13577), .B1_t (new_AGEMA_signal_13578), .B1_f (new_AGEMA_signal_13579), .Z0_t (KeyExpansionOutput[101]), .Z0_f (new_AGEMA_signal_14060), .Z1_t (new_AGEMA_signal_14061), .Z1_f (new_AGEMA_signal_14062) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U5 ( .A0_t (RoundKey[100]), .A0_f (new_AGEMA_signal_5072), .A1_t (new_AGEMA_signal_5073), .A1_f (new_AGEMA_signal_5074), .B0_t (KeyExpansionIns_tmp[4]), .B0_f (new_AGEMA_signal_13580), .B1_t (new_AGEMA_signal_13581), .B1_f (new_AGEMA_signal_13582), .Z0_t (KeyExpansionOutput[100]), .Z0_f (new_AGEMA_signal_14063), .Z1_t (new_AGEMA_signal_14064), .Z1_f (new_AGEMA_signal_14065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U4 ( .A0_t (RoundKey[0]), .A0_f (new_AGEMA_signal_5063), .A1_t (new_AGEMA_signal_5064), .A1_f (new_AGEMA_signal_5065), .B0_t (KeyExpansionOutput[32]), .B0_f (new_AGEMA_signal_15062), .B1_t (new_AGEMA_signal_15063), .B1_f (new_AGEMA_signal_15064), .Z0_t (KeyExpansionOutput[0]), .Z0_f (new_AGEMA_signal_15809), .Z1_t (new_AGEMA_signal_15810), .Z1_f (new_AGEMA_signal_15811) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U3 ( .A0_t (RoundKey[32]), .A0_f (new_AGEMA_signal_5540), .A1_t (new_AGEMA_signal_5541), .A1_f (new_AGEMA_signal_5542), .B0_t (KeyExpansionOutput[64]), .B0_f (new_AGEMA_signal_14066), .B1_t (new_AGEMA_signal_14067), .B1_f (new_AGEMA_signal_14068), .Z0_t (KeyExpansionOutput[32]), .Z0_f (new_AGEMA_signal_15062), .Z1_t (new_AGEMA_signal_15063), .Z1_f (new_AGEMA_signal_15064) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U2 ( .A0_t (RoundKey[64]), .A0_f (new_AGEMA_signal_5855), .A1_t (new_AGEMA_signal_5856), .A1_f (new_AGEMA_signal_5857), .B0_t (KeyExpansionOutput[96]), .B0_f (new_AGEMA_signal_13502), .B1_t (new_AGEMA_signal_13503), .B1_f (new_AGEMA_signal_13504), .Z0_t (KeyExpansionOutput[64]), .Z0_f (new_AGEMA_signal_14066), .Z1_t (new_AGEMA_signal_14067), .Z1_f (new_AGEMA_signal_14068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U1 ( .A0_t (RoundKey[96]), .A0_f (new_AGEMA_signal_6170), .A1_t (new_AGEMA_signal_6171), .A1_f (new_AGEMA_signal_6172), .B0_t (KeyExpansionIns_tmp[0]), .B0_f (new_AGEMA_signal_12965), .B1_t (new_AGEMA_signal_12966), .B1_f (new_AGEMA_signal_12967), .Z0_t (KeyExpansionOutput[96]), .Z0_f (new_AGEMA_signal_13502), .Z1_t (new_AGEMA_signal_13503), .Z1_f (new_AGEMA_signal_13504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U8 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_), .A0_f (new_AGEMA_signal_13508), .A1_t (new_AGEMA_signal_13509), .A1_f (new_AGEMA_signal_13510), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n283), .B1_f (new_AGEMA_signal_6344), .Z0_t (KeyExpansionIns_tmp[31]), .Z0_f (new_AGEMA_signal_14069), .Z1_t (new_AGEMA_signal_14070), .Z1_f (new_AGEMA_signal_14071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U7 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_), .A0_f (new_AGEMA_signal_13511), .A1_t (new_AGEMA_signal_13512), .A1_f (new_AGEMA_signal_13513), .B0_t (1'b0), .B0_f (1'b1), .B1_t (n285), .B1_f (new_AGEMA_signal_6345), .Z0_t (KeyExpansionIns_tmp[30]), .Z0_f (new_AGEMA_signal_14072), .Z1_t (new_AGEMA_signal_14073), .Z1_f (new_AGEMA_signal_14074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U6 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_), .A0_f (new_AGEMA_signal_13514), .A1_t (new_AGEMA_signal_13515), .A1_f (new_AGEMA_signal_13516), .B0_t (1'b0), .B0_f (1'b1), .B1_t (Rcon[5]), .B1_f (new_AGEMA_signal_7471), .Z0_t (KeyExpansionIns_tmp[29]), .Z0_f (new_AGEMA_signal_14075), .Z1_t (new_AGEMA_signal_14076), .Z1_f (new_AGEMA_signal_14077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U5 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_), .A0_f (new_AGEMA_signal_13517), .A1_t (new_AGEMA_signal_13518), .A1_f (new_AGEMA_signal_13519), .B0_t (1'b0), .B0_f (1'b1), .B1_t (Rcon[4]), .B1_f (new_AGEMA_signal_6926), .Z0_t (KeyExpansionIns_tmp[28]), .Z0_f (new_AGEMA_signal_14078), .Z1_t (new_AGEMA_signal_14079), .Z1_f (new_AGEMA_signal_14080) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U4 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_), .A0_f (new_AGEMA_signal_13520), .A1_t (new_AGEMA_signal_13521), .A1_f (new_AGEMA_signal_13522), .B0_t (1'b0), .B0_f (1'b1), .B1_t (Rcon[3]), .B1_f (new_AGEMA_signal_7470), .Z0_t (KeyExpansionIns_tmp[27]), .Z0_f (new_AGEMA_signal_14081), .Z1_t (new_AGEMA_signal_14082), .Z1_f (new_AGEMA_signal_14083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U3 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_), .A0_f (new_AGEMA_signal_13523), .A1_t (new_AGEMA_signal_13524), .A1_f (new_AGEMA_signal_13525), .B0_t (1'b0), .B0_f (1'b1), .B1_t (Rcon[2]), .B1_f (new_AGEMA_signal_7469), .Z0_t (KeyExpansionIns_tmp[26]), .Z0_f (new_AGEMA_signal_14084), .Z1_t (new_AGEMA_signal_14085), .Z1_f (new_AGEMA_signal_14086) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U2 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_), .A0_f (new_AGEMA_signal_13526), .A1_t (new_AGEMA_signal_13527), .A1_f (new_AGEMA_signal_13528), .B0_t (1'b0), .B0_f (1'b1), .B1_t (Rcon[1]), .B1_f (new_AGEMA_signal_6338), .Z0_t (KeyExpansionIns_tmp[25]), .Z0_f (new_AGEMA_signal_14087), .Z1_t (new_AGEMA_signal_14088), .Z1_f (new_AGEMA_signal_14089) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_), .A0_f (new_AGEMA_signal_12866), .A1_t (new_AGEMA_signal_12867), .A1_f (new_AGEMA_signal_12868), .B0_t (1'b0), .B0_f (1'b1), .B1_t (Rcon[0]), .B1_f (new_AGEMA_signal_6337), .Z0_t (KeyExpansionIns_tmp[24]), .Z0_f (new_AGEMA_signal_13505), .Z1_t (new_AGEMA_signal_13506), .Z1_f (new_AGEMA_signal_13507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T1_U1 ( .A0_t (RoundKey[23]), .A0_f (new_AGEMA_signal_5450), .A1_t (new_AGEMA_signal_5451), .A1_f (new_AGEMA_signal_5452), .B0_t (RoundKey[20]), .B0_f (new_AGEMA_signal_5423), .B1_t (new_AGEMA_signal_5424), .B1_f (new_AGEMA_signal_5425), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .Z0_f (new_AGEMA_signal_6213), .Z1_t (new_AGEMA_signal_6214), .Z1_f (new_AGEMA_signal_6215) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T2_U1 ( .A0_t (RoundKey[23]), .A0_f (new_AGEMA_signal_5450), .A1_t (new_AGEMA_signal_5451), .A1_f (new_AGEMA_signal_5452), .B0_t (RoundKey[18]), .B0_f (new_AGEMA_signal_5396), .B1_t (new_AGEMA_signal_5397), .B1_f (new_AGEMA_signal_5398), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .Z0_f (new_AGEMA_signal_6216), .Z1_t (new_AGEMA_signal_6217), .Z1_f (new_AGEMA_signal_6218) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T3_U1 ( .A0_t (RoundKey[23]), .A0_f (new_AGEMA_signal_5450), .A1_t (new_AGEMA_signal_5451), .A1_f (new_AGEMA_signal_5452), .B0_t (RoundKey[17]), .B0_f (new_AGEMA_signal_5387), .B1_t (new_AGEMA_signal_5388), .B1_f (new_AGEMA_signal_5389), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .Z0_f (new_AGEMA_signal_6219), .Z1_t (new_AGEMA_signal_6220), .Z1_f (new_AGEMA_signal_6221) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T4_U1 ( .A0_t (RoundKey[20]), .A0_f (new_AGEMA_signal_5423), .A1_t (new_AGEMA_signal_5424), .A1_f (new_AGEMA_signal_5425), .B0_t (RoundKey[18]), .B0_f (new_AGEMA_signal_5396), .B1_t (new_AGEMA_signal_5397), .B1_f (new_AGEMA_signal_5398), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .Z0_f (new_AGEMA_signal_6222), .Z1_t (new_AGEMA_signal_6223), .Z1_f (new_AGEMA_signal_6224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T5_U1 ( .A0_t (RoundKey[19]), .A0_f (new_AGEMA_signal_5405), .A1_t (new_AGEMA_signal_5406), .A1_f (new_AGEMA_signal_5407), .B0_t (RoundKey[17]), .B0_f (new_AGEMA_signal_5387), .B1_t (new_AGEMA_signal_5388), .B1_f (new_AGEMA_signal_5389), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .Z0_f (new_AGEMA_signal_6225), .Z1_t (new_AGEMA_signal_6226), .Z1_f (new_AGEMA_signal_6227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .A0_f (new_AGEMA_signal_6213), .A1_t (new_AGEMA_signal_6214), .A1_f (new_AGEMA_signal_6215), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .B0_f (new_AGEMA_signal_6225), .B1_t (new_AGEMA_signal_6226), .B1_f (new_AGEMA_signal_6227), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .Z0_f (new_AGEMA_signal_6826), .Z1_t (new_AGEMA_signal_6827), .Z1_f (new_AGEMA_signal_6828) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T7_U1 ( .A0_t (RoundKey[22]), .A0_f (new_AGEMA_signal_5441), .A1_t (new_AGEMA_signal_5442), .A1_f (new_AGEMA_signal_5443), .B0_t (RoundKey[21]), .B0_f (new_AGEMA_signal_5432), .B1_t (new_AGEMA_signal_5433), .B1_f (new_AGEMA_signal_5434), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .Z0_f (new_AGEMA_signal_6228), .Z1_t (new_AGEMA_signal_6229), .Z1_f (new_AGEMA_signal_6230) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T8_U1 ( .A0_t (RoundKey[16]), .A0_f (new_AGEMA_signal_5378), .A1_t (new_AGEMA_signal_5379), .A1_f (new_AGEMA_signal_5380), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .B0_f (new_AGEMA_signal_6826), .B1_t (new_AGEMA_signal_6827), .B1_f (new_AGEMA_signal_6828), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .Z0_f (new_AGEMA_signal_7312), .Z1_t (new_AGEMA_signal_7313), .Z1_f (new_AGEMA_signal_7314) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T9_U1 ( .A0_t (RoundKey[16]), .A0_f (new_AGEMA_signal_5378), .A1_t (new_AGEMA_signal_5379), .A1_f (new_AGEMA_signal_5380), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .B0_f (new_AGEMA_signal_6228), .B1_t (new_AGEMA_signal_6229), .B1_f (new_AGEMA_signal_6230), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .Z0_f (new_AGEMA_signal_6829), .Z1_t (new_AGEMA_signal_6830), .Z1_f (new_AGEMA_signal_6831) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .A0_f (new_AGEMA_signal_6826), .A1_t (new_AGEMA_signal_6827), .A1_f (new_AGEMA_signal_6828), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .B0_f (new_AGEMA_signal_6228), .B1_t (new_AGEMA_signal_6229), .B1_f (new_AGEMA_signal_6230), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .Z0_f (new_AGEMA_signal_7315), .Z1_t (new_AGEMA_signal_7316), .Z1_f (new_AGEMA_signal_7317) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T11_U1 ( .A0_t (RoundKey[22]), .A0_f (new_AGEMA_signal_5441), .A1_t (new_AGEMA_signal_5442), .A1_f (new_AGEMA_signal_5443), .B0_t (RoundKey[18]), .B0_f (new_AGEMA_signal_5396), .B1_t (new_AGEMA_signal_5397), .B1_f (new_AGEMA_signal_5398), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11), .Z0_f (new_AGEMA_signal_6231), .Z1_t (new_AGEMA_signal_6232), .Z1_f (new_AGEMA_signal_6233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T12_U1 ( .A0_t (RoundKey[21]), .A0_f (new_AGEMA_signal_5432), .A1_t (new_AGEMA_signal_5433), .A1_f (new_AGEMA_signal_5434), .B0_t (RoundKey[18]), .B0_f (new_AGEMA_signal_5396), .B1_t (new_AGEMA_signal_5397), .B1_f (new_AGEMA_signal_5398), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12), .Z0_f (new_AGEMA_signal_6234), .Z1_t (new_AGEMA_signal_6235), .Z1_f (new_AGEMA_signal_6236) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .A0_f (new_AGEMA_signal_6219), .A1_t (new_AGEMA_signal_6220), .A1_f (new_AGEMA_signal_6221), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .B0_f (new_AGEMA_signal_6222), .B1_t (new_AGEMA_signal_6223), .B1_f (new_AGEMA_signal_6224), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .Z0_f (new_AGEMA_signal_6832), .Z1_t (new_AGEMA_signal_6833), .Z1_f (new_AGEMA_signal_6834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .A0_f (new_AGEMA_signal_6826), .A1_t (new_AGEMA_signal_6827), .A1_f (new_AGEMA_signal_6828), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11), .B0_f (new_AGEMA_signal_6231), .B1_t (new_AGEMA_signal_6232), .B1_f (new_AGEMA_signal_6233), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14), .Z0_f (new_AGEMA_signal_7318), .Z1_t (new_AGEMA_signal_7319), .Z1_f (new_AGEMA_signal_7320) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .A0_f (new_AGEMA_signal_6225), .A1_t (new_AGEMA_signal_6226), .A1_f (new_AGEMA_signal_6227), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11), .B0_f (new_AGEMA_signal_6231), .B1_t (new_AGEMA_signal_6232), .B1_f (new_AGEMA_signal_6233), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .Z0_f (new_AGEMA_signal_6835), .Z1_t (new_AGEMA_signal_6836), .Z1_f (new_AGEMA_signal_6837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .A0_f (new_AGEMA_signal_6225), .A1_t (new_AGEMA_signal_6226), .A1_f (new_AGEMA_signal_6227), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12), .B0_f (new_AGEMA_signal_6234), .B1_t (new_AGEMA_signal_6235), .B1_f (new_AGEMA_signal_6236), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Z0_f (new_AGEMA_signal_6838), .Z1_t (new_AGEMA_signal_6839), .Z1_f (new_AGEMA_signal_6840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .A0_f (new_AGEMA_signal_6829), .A1_t (new_AGEMA_signal_6830), .A1_f (new_AGEMA_signal_6831), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .B0_f (new_AGEMA_signal_6838), .B1_t (new_AGEMA_signal_6839), .B1_f (new_AGEMA_signal_6840), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .Z0_f (new_AGEMA_signal_7321), .Z1_t (new_AGEMA_signal_7322), .Z1_f (new_AGEMA_signal_7323) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T18_U1 ( .A0_t (RoundKey[20]), .A0_f (new_AGEMA_signal_5423), .A1_t (new_AGEMA_signal_5424), .A1_f (new_AGEMA_signal_5425), .B0_t (RoundKey[16]), .B0_f (new_AGEMA_signal_5378), .B1_t (new_AGEMA_signal_5379), .B1_f (new_AGEMA_signal_5380), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18), .Z0_f (new_AGEMA_signal_6237), .Z1_t (new_AGEMA_signal_6238), .Z1_f (new_AGEMA_signal_6239) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .A0_f (new_AGEMA_signal_6228), .A1_t (new_AGEMA_signal_6229), .A1_f (new_AGEMA_signal_6230), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18), .B0_f (new_AGEMA_signal_6237), .B1_t (new_AGEMA_signal_6238), .B1_f (new_AGEMA_signal_6239), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .Z0_f (new_AGEMA_signal_6841), .Z1_t (new_AGEMA_signal_6842), .Z1_f (new_AGEMA_signal_6843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .A0_f (new_AGEMA_signal_6213), .A1_t (new_AGEMA_signal_6214), .A1_f (new_AGEMA_signal_6215), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .B0_f (new_AGEMA_signal_6841), .B1_t (new_AGEMA_signal_6842), .B1_f (new_AGEMA_signal_6843), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .Z0_f (new_AGEMA_signal_7324), .Z1_t (new_AGEMA_signal_7325), .Z1_f (new_AGEMA_signal_7326) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T21_U1 ( .A0_t (RoundKey[17]), .A0_f (new_AGEMA_signal_5387), .A1_t (new_AGEMA_signal_5388), .A1_f (new_AGEMA_signal_5389), .B0_t (RoundKey[16]), .B0_f (new_AGEMA_signal_5378), .B1_t (new_AGEMA_signal_5379), .B1_f (new_AGEMA_signal_5380), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21), .Z0_f (new_AGEMA_signal_6240), .Z1_t (new_AGEMA_signal_6241), .Z1_f (new_AGEMA_signal_6242) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .A0_f (new_AGEMA_signal_6228), .A1_t (new_AGEMA_signal_6229), .A1_f (new_AGEMA_signal_6230), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21), .B0_f (new_AGEMA_signal_6240), .B1_t (new_AGEMA_signal_6241), .B1_f (new_AGEMA_signal_6242), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .Z0_f (new_AGEMA_signal_6844), .Z1_t (new_AGEMA_signal_6845), .Z1_f (new_AGEMA_signal_6846) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .A0_f (new_AGEMA_signal_6216), .A1_t (new_AGEMA_signal_6217), .A1_f (new_AGEMA_signal_6218), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .B0_f (new_AGEMA_signal_6844), .B1_t (new_AGEMA_signal_6845), .B1_f (new_AGEMA_signal_6846), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .Z0_f (new_AGEMA_signal_7327), .Z1_t (new_AGEMA_signal_7328), .Z1_f (new_AGEMA_signal_7329) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .A0_f (new_AGEMA_signal_6216), .A1_t (new_AGEMA_signal_6217), .A1_f (new_AGEMA_signal_6218), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .B0_f (new_AGEMA_signal_7315), .B1_t (new_AGEMA_signal_7316), .B1_f (new_AGEMA_signal_7317), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24), .Z0_f (new_AGEMA_signal_8096), .Z1_t (new_AGEMA_signal_8097), .Z1_f (new_AGEMA_signal_8098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .A0_f (new_AGEMA_signal_7324), .A1_t (new_AGEMA_signal_7325), .A1_f (new_AGEMA_signal_7326), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .B0_f (new_AGEMA_signal_7321), .B1_t (new_AGEMA_signal_7322), .B1_f (new_AGEMA_signal_7323), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25), .Z0_f (new_AGEMA_signal_8099), .Z1_t (new_AGEMA_signal_8100), .Z1_f (new_AGEMA_signal_8101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .A0_f (new_AGEMA_signal_6219), .A1_t (new_AGEMA_signal_6220), .A1_f (new_AGEMA_signal_6221), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .B0_f (new_AGEMA_signal_6838), .B1_t (new_AGEMA_signal_6839), .B1_f (new_AGEMA_signal_6840), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26), .Z0_f (new_AGEMA_signal_7330), .Z1_t (new_AGEMA_signal_7331), .Z1_f (new_AGEMA_signal_7332) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .A0_f (new_AGEMA_signal_6213), .A1_t (new_AGEMA_signal_6214), .A1_f (new_AGEMA_signal_6215), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12), .B0_f (new_AGEMA_signal_6234), .B1_t (new_AGEMA_signal_6235), .B1_f (new_AGEMA_signal_6236), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .Z0_f (new_AGEMA_signal_6847), .Z1_t (new_AGEMA_signal_6848), .Z1_f (new_AGEMA_signal_6849) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .A0_f (new_AGEMA_signal_6832), .A1_t (new_AGEMA_signal_6833), .A1_f (new_AGEMA_signal_6834), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .B0_f (new_AGEMA_signal_6826), .B1_t (new_AGEMA_signal_6827), .B1_f (new_AGEMA_signal_6828), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1), .Z0_f (new_AGEMA_signal_7333), .Z1_t (new_AGEMA_signal_7334), .Z1_f (new_AGEMA_signal_7335) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .A0_f (new_AGEMA_signal_7327), .A1_t (new_AGEMA_signal_7328), .A1_f (new_AGEMA_signal_7329), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .B0_f (new_AGEMA_signal_7312), .B1_t (new_AGEMA_signal_7313), .B1_f (new_AGEMA_signal_7314), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2), .Z0_f (new_AGEMA_signal_8102), .Z1_t (new_AGEMA_signal_8103), .Z1_f (new_AGEMA_signal_8104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14), .A0_f (new_AGEMA_signal_7318), .A1_t (new_AGEMA_signal_7319), .A1_f (new_AGEMA_signal_7320), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1), .B0_f (new_AGEMA_signal_7333), .B1_t (new_AGEMA_signal_7334), .B1_f (new_AGEMA_signal_7335), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3), .Z0_f (new_AGEMA_signal_8105), .Z1_t (new_AGEMA_signal_8106), .Z1_f (new_AGEMA_signal_8107) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .A0_f (new_AGEMA_signal_6841), .A1_t (new_AGEMA_signal_6842), .A1_f (new_AGEMA_signal_6843), .B0_t (RoundKey[16]), .B0_f (new_AGEMA_signal_5378), .B1_t (new_AGEMA_signal_5379), .B1_f (new_AGEMA_signal_5380), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4), .Z0_f (new_AGEMA_signal_7336), .Z1_t (new_AGEMA_signal_7337), .Z1_f (new_AGEMA_signal_7338) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4), .A0_f (new_AGEMA_signal_7336), .A1_t (new_AGEMA_signal_7337), .A1_f (new_AGEMA_signal_7338), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1), .B0_f (new_AGEMA_signal_7333), .B1_t (new_AGEMA_signal_7334), .B1_f (new_AGEMA_signal_7335), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5), .Z0_f (new_AGEMA_signal_8108), .Z1_t (new_AGEMA_signal_8109), .Z1_f (new_AGEMA_signal_8110) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .A0_f (new_AGEMA_signal_6219), .A1_t (new_AGEMA_signal_6220), .A1_f (new_AGEMA_signal_6221), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .B0_f (new_AGEMA_signal_6838), .B1_t (new_AGEMA_signal_6839), .B1_f (new_AGEMA_signal_6840), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6), .Z0_f (new_AGEMA_signal_7339), .Z1_t (new_AGEMA_signal_7340), .Z1_f (new_AGEMA_signal_7341) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .A0_f (new_AGEMA_signal_6844), .A1_t (new_AGEMA_signal_6845), .A1_f (new_AGEMA_signal_6846), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .B0_f (new_AGEMA_signal_6829), .B1_t (new_AGEMA_signal_6830), .B1_f (new_AGEMA_signal_6831), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7), .Z0_f (new_AGEMA_signal_7342), .Z1_t (new_AGEMA_signal_7343), .Z1_f (new_AGEMA_signal_7344) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26), .A0_f (new_AGEMA_signal_7330), .A1_t (new_AGEMA_signal_7331), .A1_f (new_AGEMA_signal_7332), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6), .B0_f (new_AGEMA_signal_7339), .B1_t (new_AGEMA_signal_7340), .B1_f (new_AGEMA_signal_7341), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8), .Z0_f (new_AGEMA_signal_8111), .Z1_t (new_AGEMA_signal_8112), .Z1_f (new_AGEMA_signal_8113) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .A0_f (new_AGEMA_signal_7324), .A1_t (new_AGEMA_signal_7325), .A1_f (new_AGEMA_signal_7326), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .B0_f (new_AGEMA_signal_7321), .B1_t (new_AGEMA_signal_7322), .B1_f (new_AGEMA_signal_7323), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9), .Z0_f (new_AGEMA_signal_8114), .Z1_t (new_AGEMA_signal_8115), .Z1_f (new_AGEMA_signal_8116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9), .A0_f (new_AGEMA_signal_8114), .A1_t (new_AGEMA_signal_8115), .A1_f (new_AGEMA_signal_8116), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6), .B0_f (new_AGEMA_signal_7339), .B1_t (new_AGEMA_signal_7340), .B1_f (new_AGEMA_signal_7341), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10), .Z0_f (new_AGEMA_signal_8636), .Z1_t (new_AGEMA_signal_8637), .Z1_f (new_AGEMA_signal_8638) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .A0_f (new_AGEMA_signal_6213), .A1_t (new_AGEMA_signal_6214), .A1_f (new_AGEMA_signal_6215), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .B0_f (new_AGEMA_signal_6835), .B1_t (new_AGEMA_signal_6836), .B1_f (new_AGEMA_signal_6837), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11), .Z0_f (new_AGEMA_signal_7345), .Z1_t (new_AGEMA_signal_7346), .Z1_f (new_AGEMA_signal_7347) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .A0_f (new_AGEMA_signal_6222), .A1_t (new_AGEMA_signal_6223), .A1_f (new_AGEMA_signal_6224), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .B0_f (new_AGEMA_signal_6847), .B1_t (new_AGEMA_signal_6848), .B1_f (new_AGEMA_signal_6849), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12), .Z0_f (new_AGEMA_signal_7348), .Z1_t (new_AGEMA_signal_7349), .Z1_f (new_AGEMA_signal_7350) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12), .A0_f (new_AGEMA_signal_7348), .A1_t (new_AGEMA_signal_7349), .A1_f (new_AGEMA_signal_7350), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11), .B0_f (new_AGEMA_signal_7345), .B1_t (new_AGEMA_signal_7346), .B1_f (new_AGEMA_signal_7347), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13), .Z0_f (new_AGEMA_signal_8117), .Z1_t (new_AGEMA_signal_8118), .Z1_f (new_AGEMA_signal_8119) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .A0_f (new_AGEMA_signal_6216), .A1_t (new_AGEMA_signal_6217), .A1_f (new_AGEMA_signal_6218), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .B0_f (new_AGEMA_signal_7315), .B1_t (new_AGEMA_signal_7316), .B1_f (new_AGEMA_signal_7317), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14), .Z0_f (new_AGEMA_signal_8120), .Z1_t (new_AGEMA_signal_8121), .Z1_f (new_AGEMA_signal_8122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14), .A0_f (new_AGEMA_signal_8120), .A1_t (new_AGEMA_signal_8121), .A1_f (new_AGEMA_signal_8122), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11), .B0_f (new_AGEMA_signal_7345), .B1_t (new_AGEMA_signal_7346), .B1_f (new_AGEMA_signal_7347), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15), .Z0_f (new_AGEMA_signal_8639), .Z1_t (new_AGEMA_signal_8640), .Z1_f (new_AGEMA_signal_8641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3), .A0_f (new_AGEMA_signal_8105), .A1_t (new_AGEMA_signal_8106), .A1_f (new_AGEMA_signal_8107), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2), .B0_f (new_AGEMA_signal_8102), .B1_t (new_AGEMA_signal_8103), .B1_f (new_AGEMA_signal_8104), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16), .Z0_f (new_AGEMA_signal_8642), .Z1_t (new_AGEMA_signal_8643), .Z1_f (new_AGEMA_signal_8644) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5), .A0_f (new_AGEMA_signal_8108), .A1_t (new_AGEMA_signal_8109), .A1_f (new_AGEMA_signal_8110), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24), .B0_f (new_AGEMA_signal_8096), .B1_t (new_AGEMA_signal_8097), .B1_f (new_AGEMA_signal_8098), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17), .Z0_f (new_AGEMA_signal_8645), .Z1_t (new_AGEMA_signal_8646), .Z1_f (new_AGEMA_signal_8647) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8), .A0_f (new_AGEMA_signal_8111), .A1_t (new_AGEMA_signal_8112), .A1_f (new_AGEMA_signal_8113), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7), .B0_f (new_AGEMA_signal_7342), .B1_t (new_AGEMA_signal_7343), .B1_f (new_AGEMA_signal_7344), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18), .Z0_f (new_AGEMA_signal_8648), .Z1_t (new_AGEMA_signal_8649), .Z1_f (new_AGEMA_signal_8650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10), .A0_f (new_AGEMA_signal_8636), .A1_t (new_AGEMA_signal_8637), .A1_f (new_AGEMA_signal_8638), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15), .B0_f (new_AGEMA_signal_8639), .B1_t (new_AGEMA_signal_8640), .B1_f (new_AGEMA_signal_8641), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19), .Z0_f (new_AGEMA_signal_8936), .Z1_t (new_AGEMA_signal_8937), .Z1_f (new_AGEMA_signal_8938) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16), .A0_f (new_AGEMA_signal_8642), .A1_t (new_AGEMA_signal_8643), .A1_f (new_AGEMA_signal_8644), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13), .B0_f (new_AGEMA_signal_8117), .B1_t (new_AGEMA_signal_8118), .B1_f (new_AGEMA_signal_8119), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .Z0_f (new_AGEMA_signal_8939), .Z1_t (new_AGEMA_signal_8940), .Z1_f (new_AGEMA_signal_8941) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17), .A0_f (new_AGEMA_signal_8645), .A1_t (new_AGEMA_signal_8646), .A1_f (new_AGEMA_signal_8647), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15), .B0_f (new_AGEMA_signal_8639), .B1_t (new_AGEMA_signal_8640), .B1_f (new_AGEMA_signal_8641), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .Z0_f (new_AGEMA_signal_8942), .Z1_t (new_AGEMA_signal_8943), .Z1_f (new_AGEMA_signal_8944) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18), .A0_f (new_AGEMA_signal_8648), .A1_t (new_AGEMA_signal_8649), .A1_f (new_AGEMA_signal_8650), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13), .B0_f (new_AGEMA_signal_8117), .B1_t (new_AGEMA_signal_8118), .B1_f (new_AGEMA_signal_8119), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .Z0_f (new_AGEMA_signal_8945), .Z1_t (new_AGEMA_signal_8946), .Z1_f (new_AGEMA_signal_8947) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19), .A0_f (new_AGEMA_signal_8936), .A1_t (new_AGEMA_signal_8937), .A1_f (new_AGEMA_signal_8938), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25), .B0_f (new_AGEMA_signal_8099), .B1_t (new_AGEMA_signal_8100), .B1_f (new_AGEMA_signal_8101), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .Z0_f (new_AGEMA_signal_9176), .Z1_t (new_AGEMA_signal_9177), .Z1_f (new_AGEMA_signal_9178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .A0_f (new_AGEMA_signal_8945), .A1_t (new_AGEMA_signal_8946), .A1_f (new_AGEMA_signal_8947), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .B0_f (new_AGEMA_signal_9176), .B1_t (new_AGEMA_signal_9177), .B1_f (new_AGEMA_signal_9178), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .Z0_f (new_AGEMA_signal_9416), .Z1_t (new_AGEMA_signal_9417), .Z1_f (new_AGEMA_signal_9418) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .A0_f (new_AGEMA_signal_8945), .A1_t (new_AGEMA_signal_8946), .A1_f (new_AGEMA_signal_8947), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .B0_f (new_AGEMA_signal_8939), .B1_t (new_AGEMA_signal_8940), .B1_f (new_AGEMA_signal_8941), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z0_f (new_AGEMA_signal_9179), .Z1_t (new_AGEMA_signal_9180), .Z1_f (new_AGEMA_signal_9181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .A0_f (new_AGEMA_signal_8942), .A1_t (new_AGEMA_signal_8943), .A1_f (new_AGEMA_signal_8944), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .B0_f (new_AGEMA_signal_9179), .B1_t (new_AGEMA_signal_9180), .B1_f (new_AGEMA_signal_9181), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26), .Z0_f (new_AGEMA_signal_9419), .Z1_t (new_AGEMA_signal_9420), .Z1_f (new_AGEMA_signal_9421) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .A0_f (new_AGEMA_signal_8939), .A1_t (new_AGEMA_signal_8940), .A1_f (new_AGEMA_signal_8941), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .B0_f (new_AGEMA_signal_8942), .B1_t (new_AGEMA_signal_8943), .B1_f (new_AGEMA_signal_8944), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .Z0_f (new_AGEMA_signal_9182), .Z1_t (new_AGEMA_signal_9183), .Z1_f (new_AGEMA_signal_9184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .A0_f (new_AGEMA_signal_9176), .A1_t (new_AGEMA_signal_9177), .A1_f (new_AGEMA_signal_9178), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .B0_f (new_AGEMA_signal_9179), .B1_t (new_AGEMA_signal_9180), .B1_f (new_AGEMA_signal_9181), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28), .Z0_f (new_AGEMA_signal_9422), .Z1_t (new_AGEMA_signal_9423), .Z1_f (new_AGEMA_signal_9424) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28), .A0_f (new_AGEMA_signal_9422), .A1_t (new_AGEMA_signal_9423), .A1_f (new_AGEMA_signal_9424), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .B0_f (new_AGEMA_signal_9182), .B1_t (new_AGEMA_signal_9183), .B1_f (new_AGEMA_signal_9184), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29), .Z0_f (new_AGEMA_signal_9716), .Z1_t (new_AGEMA_signal_9717), .Z1_f (new_AGEMA_signal_9718) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M30_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26), .A0_f (new_AGEMA_signal_9419), .A1_t (new_AGEMA_signal_9420), .A1_f (new_AGEMA_signal_9421), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .B0_f (new_AGEMA_signal_9416), .B1_t (new_AGEMA_signal_9417), .B1_f (new_AGEMA_signal_9418), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30), .Z0_f (new_AGEMA_signal_9719), .Z1_t (new_AGEMA_signal_9720), .Z1_f (new_AGEMA_signal_9721) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M31_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .A0_f (new_AGEMA_signal_8939), .A1_t (new_AGEMA_signal_8940), .A1_f (new_AGEMA_signal_8941), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .B0_f (new_AGEMA_signal_9176), .B1_t (new_AGEMA_signal_9177), .B1_f (new_AGEMA_signal_9178), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31), .Z0_f (new_AGEMA_signal_9425), .Z1_t (new_AGEMA_signal_9426), .Z1_f (new_AGEMA_signal_9427) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M32_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .A0_f (new_AGEMA_signal_9182), .A1_t (new_AGEMA_signal_9183), .A1_f (new_AGEMA_signal_9184), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31), .B0_f (new_AGEMA_signal_9425), .B1_t (new_AGEMA_signal_9426), .B1_f (new_AGEMA_signal_9427), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32), .Z0_f (new_AGEMA_signal_9722), .Z1_t (new_AGEMA_signal_9723), .Z1_f (new_AGEMA_signal_9724) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M33_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .A0_f (new_AGEMA_signal_9182), .A1_t (new_AGEMA_signal_9183), .A1_f (new_AGEMA_signal_9184), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .B0_f (new_AGEMA_signal_9179), .B1_t (new_AGEMA_signal_9180), .B1_f (new_AGEMA_signal_9181), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33), .Z0_f (new_AGEMA_signal_9428), .Z1_t (new_AGEMA_signal_9429), .Z1_f (new_AGEMA_signal_9430) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M34_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .A0_f (new_AGEMA_signal_8942), .A1_t (new_AGEMA_signal_8943), .A1_f (new_AGEMA_signal_8944), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .B0_f (new_AGEMA_signal_8945), .B1_t (new_AGEMA_signal_8946), .B1_f (new_AGEMA_signal_8947), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34), .Z0_f (new_AGEMA_signal_9185), .Z1_t (new_AGEMA_signal_9186), .Z1_f (new_AGEMA_signal_9187) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M35_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .A0_f (new_AGEMA_signal_9416), .A1_t (new_AGEMA_signal_9417), .A1_f (new_AGEMA_signal_9418), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34), .B0_f (new_AGEMA_signal_9185), .B1_t (new_AGEMA_signal_9186), .B1_f (new_AGEMA_signal_9187), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35), .Z0_f (new_AGEMA_signal_9725), .Z1_t (new_AGEMA_signal_9726), .Z1_f (new_AGEMA_signal_9727) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M36_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .A0_f (new_AGEMA_signal_9416), .A1_t (new_AGEMA_signal_9417), .A1_f (new_AGEMA_signal_9418), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .B0_f (new_AGEMA_signal_9179), .B1_t (new_AGEMA_signal_9180), .B1_f (new_AGEMA_signal_9181), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36), .Z0_f (new_AGEMA_signal_9728), .Z1_t (new_AGEMA_signal_9729), .Z1_f (new_AGEMA_signal_9730) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M37_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .A0_f (new_AGEMA_signal_8942), .A1_t (new_AGEMA_signal_8943), .A1_f (new_AGEMA_signal_8944), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29), .B0_f (new_AGEMA_signal_9716), .B1_t (new_AGEMA_signal_9717), .B1_f (new_AGEMA_signal_9718), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .Z0_f (new_AGEMA_signal_10016), .Z1_t (new_AGEMA_signal_10017), .Z1_f (new_AGEMA_signal_10018) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M38_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32), .A0_f (new_AGEMA_signal_9722), .A1_t (new_AGEMA_signal_9723), .A1_f (new_AGEMA_signal_9724), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33), .B0_f (new_AGEMA_signal_9428), .B1_t (new_AGEMA_signal_9429), .B1_f (new_AGEMA_signal_9430), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .Z0_f (new_AGEMA_signal_10019), .Z1_t (new_AGEMA_signal_10020), .Z1_f (new_AGEMA_signal_10021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M39_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .A0_f (new_AGEMA_signal_9176), .A1_t (new_AGEMA_signal_9177), .A1_f (new_AGEMA_signal_9178), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30), .B0_f (new_AGEMA_signal_9719), .B1_t (new_AGEMA_signal_9720), .B1_f (new_AGEMA_signal_9721), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .Z0_f (new_AGEMA_signal_10022), .Z1_t (new_AGEMA_signal_10023), .Z1_f (new_AGEMA_signal_10024) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M40_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35), .A0_f (new_AGEMA_signal_9725), .A1_t (new_AGEMA_signal_9726), .A1_f (new_AGEMA_signal_9727), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36), .B0_f (new_AGEMA_signal_9728), .B1_t (new_AGEMA_signal_9729), .B1_f (new_AGEMA_signal_9730), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .Z0_f (new_AGEMA_signal_10025), .Z1_t (new_AGEMA_signal_10026), .Z1_f (new_AGEMA_signal_10027) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M41_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .A0_f (new_AGEMA_signal_10019), .A1_t (new_AGEMA_signal_10020), .A1_f (new_AGEMA_signal_10021), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .B0_f (new_AGEMA_signal_10025), .B1_t (new_AGEMA_signal_10026), .B1_f (new_AGEMA_signal_10027), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .Z0_f (new_AGEMA_signal_10256), .Z1_t (new_AGEMA_signal_10257), .Z1_f (new_AGEMA_signal_10258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M42_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .A0_f (new_AGEMA_signal_10016), .A1_t (new_AGEMA_signal_10017), .A1_f (new_AGEMA_signal_10018), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .B0_f (new_AGEMA_signal_10022), .B1_t (new_AGEMA_signal_10023), .B1_f (new_AGEMA_signal_10024), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .Z0_f (new_AGEMA_signal_10259), .Z1_t (new_AGEMA_signal_10260), .Z1_f (new_AGEMA_signal_10261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M43_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .A0_f (new_AGEMA_signal_10016), .A1_t (new_AGEMA_signal_10017), .A1_f (new_AGEMA_signal_10018), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .B0_f (new_AGEMA_signal_10019), .B1_t (new_AGEMA_signal_10020), .B1_f (new_AGEMA_signal_10021), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43), .Z0_f (new_AGEMA_signal_10262), .Z1_t (new_AGEMA_signal_10263), .Z1_f (new_AGEMA_signal_10264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M44_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .A0_f (new_AGEMA_signal_10022), .A1_t (new_AGEMA_signal_10023), .A1_f (new_AGEMA_signal_10024), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .B0_f (new_AGEMA_signal_10025), .B1_t (new_AGEMA_signal_10026), .B1_f (new_AGEMA_signal_10027), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44), .Z0_f (new_AGEMA_signal_10265), .Z1_t (new_AGEMA_signal_10266), .Z1_f (new_AGEMA_signal_10267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M45_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .A0_f (new_AGEMA_signal_10259), .A1_t (new_AGEMA_signal_10260), .A1_f (new_AGEMA_signal_10261), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .B0_f (new_AGEMA_signal_10256), .B1_t (new_AGEMA_signal_10257), .B1_f (new_AGEMA_signal_10258), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45), .Z0_f (new_AGEMA_signal_10976), .Z1_t (new_AGEMA_signal_10977), .Z1_f (new_AGEMA_signal_10978) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M46_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44), .A0_f (new_AGEMA_signal_10265), .A1_t (new_AGEMA_signal_10266), .A1_f (new_AGEMA_signal_10267), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .B0_f (new_AGEMA_signal_6826), .B1_t (new_AGEMA_signal_6827), .B1_f (new_AGEMA_signal_6828), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46), .Z0_f (new_AGEMA_signal_10979), .Z1_t (new_AGEMA_signal_10980), .Z1_f (new_AGEMA_signal_10981) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M47_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .A0_f (new_AGEMA_signal_10025), .A1_t (new_AGEMA_signal_10026), .A1_f (new_AGEMA_signal_10027), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .B0_f (new_AGEMA_signal_7312), .B1_t (new_AGEMA_signal_7313), .B1_f (new_AGEMA_signal_7314), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47), .Z0_f (new_AGEMA_signal_10268), .Z1_t (new_AGEMA_signal_10269), .Z1_f (new_AGEMA_signal_10270) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M48_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .A0_f (new_AGEMA_signal_10022), .A1_t (new_AGEMA_signal_10023), .A1_f (new_AGEMA_signal_10024), .B0_t (RoundKey[16]), .B0_f (new_AGEMA_signal_5378), .B1_t (new_AGEMA_signal_5379), .B1_f (new_AGEMA_signal_5380), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48), .Z0_f (new_AGEMA_signal_10271), .Z1_t (new_AGEMA_signal_10272), .Z1_f (new_AGEMA_signal_10273) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M49_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43), .A0_f (new_AGEMA_signal_10262), .A1_t (new_AGEMA_signal_10263), .A1_f (new_AGEMA_signal_10264), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .B0_f (new_AGEMA_signal_6838), .B1_t (new_AGEMA_signal_6839), .B1_f (new_AGEMA_signal_6840), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49), .Z0_f (new_AGEMA_signal_10982), .Z1_t (new_AGEMA_signal_10983), .Z1_f (new_AGEMA_signal_10984) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M50_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .A0_f (new_AGEMA_signal_10019), .A1_t (new_AGEMA_signal_10020), .A1_f (new_AGEMA_signal_10021), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .B0_f (new_AGEMA_signal_6829), .B1_t (new_AGEMA_signal_6830), .B1_f (new_AGEMA_signal_6831), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50), .Z0_f (new_AGEMA_signal_10274), .Z1_t (new_AGEMA_signal_10275), .Z1_f (new_AGEMA_signal_10276) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M51_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .A0_f (new_AGEMA_signal_10016), .A1_t (new_AGEMA_signal_10017), .A1_f (new_AGEMA_signal_10018), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .B0_f (new_AGEMA_signal_7321), .B1_t (new_AGEMA_signal_7322), .B1_f (new_AGEMA_signal_7323), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51), .Z0_f (new_AGEMA_signal_10277), .Z1_t (new_AGEMA_signal_10278), .Z1_f (new_AGEMA_signal_10279) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M52_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .A0_f (new_AGEMA_signal_10259), .A1_t (new_AGEMA_signal_10260), .A1_f (new_AGEMA_signal_10261), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .B0_f (new_AGEMA_signal_6835), .B1_t (new_AGEMA_signal_6836), .B1_f (new_AGEMA_signal_6837), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52), .Z0_f (new_AGEMA_signal_10985), .Z1_t (new_AGEMA_signal_10986), .Z1_f (new_AGEMA_signal_10987) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M53_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45), .A0_f (new_AGEMA_signal_10976), .A1_t (new_AGEMA_signal_10977), .A1_f (new_AGEMA_signal_10978), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .B0_f (new_AGEMA_signal_6847), .B1_t (new_AGEMA_signal_6848), .B1_f (new_AGEMA_signal_6849), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53), .Z0_f (new_AGEMA_signal_11696), .Z1_t (new_AGEMA_signal_11697), .Z1_f (new_AGEMA_signal_11698) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M54_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .A0_f (new_AGEMA_signal_10256), .A1_t (new_AGEMA_signal_10257), .A1_f (new_AGEMA_signal_10258), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .B0_f (new_AGEMA_signal_7315), .B1_t (new_AGEMA_signal_7316), .B1_f (new_AGEMA_signal_7317), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54), .Z0_f (new_AGEMA_signal_10988), .Z1_t (new_AGEMA_signal_10989), .Z1_f (new_AGEMA_signal_10990) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M55_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44), .A0_f (new_AGEMA_signal_10265), .A1_t (new_AGEMA_signal_10266), .A1_f (new_AGEMA_signal_10267), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .B0_f (new_AGEMA_signal_6832), .B1_t (new_AGEMA_signal_6833), .B1_f (new_AGEMA_signal_6834), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55), .Z0_f (new_AGEMA_signal_10991), .Z1_t (new_AGEMA_signal_10992), .Z1_f (new_AGEMA_signal_10993) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M56_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .A0_f (new_AGEMA_signal_10025), .A1_t (new_AGEMA_signal_10026), .A1_f (new_AGEMA_signal_10027), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .B0_f (new_AGEMA_signal_7327), .B1_t (new_AGEMA_signal_7328), .B1_f (new_AGEMA_signal_7329), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56), .Z0_f (new_AGEMA_signal_10280), .Z1_t (new_AGEMA_signal_10281), .Z1_f (new_AGEMA_signal_10282) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M57_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .A0_f (new_AGEMA_signal_10022), .A1_t (new_AGEMA_signal_10023), .A1_f (new_AGEMA_signal_10024), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .B0_f (new_AGEMA_signal_6841), .B1_t (new_AGEMA_signal_6842), .B1_f (new_AGEMA_signal_6843), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57), .Z0_f (new_AGEMA_signal_10283), .Z1_t (new_AGEMA_signal_10284), .Z1_f (new_AGEMA_signal_10285) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M58_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43), .A0_f (new_AGEMA_signal_10262), .A1_t (new_AGEMA_signal_10263), .A1_f (new_AGEMA_signal_10264), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .B0_f (new_AGEMA_signal_6219), .B1_t (new_AGEMA_signal_6220), .B1_f (new_AGEMA_signal_6221), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58), .Z0_f (new_AGEMA_signal_10994), .Z1_t (new_AGEMA_signal_10995), .Z1_f (new_AGEMA_signal_10996) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M59_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .A0_f (new_AGEMA_signal_10019), .A1_t (new_AGEMA_signal_10020), .A1_f (new_AGEMA_signal_10021), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .B0_f (new_AGEMA_signal_6844), .B1_t (new_AGEMA_signal_6845), .B1_f (new_AGEMA_signal_6846), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59), .Z0_f (new_AGEMA_signal_10286), .Z1_t (new_AGEMA_signal_10287), .Z1_f (new_AGEMA_signal_10288) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M60_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .A0_f (new_AGEMA_signal_10016), .A1_t (new_AGEMA_signal_10017), .A1_f (new_AGEMA_signal_10018), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .B0_f (new_AGEMA_signal_7324), .B1_t (new_AGEMA_signal_7325), .B1_f (new_AGEMA_signal_7326), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60), .Z0_f (new_AGEMA_signal_10289), .Z1_t (new_AGEMA_signal_10290), .Z1_f (new_AGEMA_signal_10291) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M61_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .A0_f (new_AGEMA_signal_10259), .A1_t (new_AGEMA_signal_10260), .A1_f (new_AGEMA_signal_10261), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .B0_f (new_AGEMA_signal_6213), .B1_t (new_AGEMA_signal_6214), .B1_f (new_AGEMA_signal_6215), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .Z0_f (new_AGEMA_signal_10997), .Z1_t (new_AGEMA_signal_10998), .Z1_f (new_AGEMA_signal_10999) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M62_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45), .A0_f (new_AGEMA_signal_10976), .A1_t (new_AGEMA_signal_10977), .A1_f (new_AGEMA_signal_10978), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .B0_f (new_AGEMA_signal_6222), .B1_t (new_AGEMA_signal_6223), .B1_f (new_AGEMA_signal_6224), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62), .Z0_f (new_AGEMA_signal_11699), .Z1_t (new_AGEMA_signal_11700), .Z1_f (new_AGEMA_signal_11701) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M63_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .A0_f (new_AGEMA_signal_10256), .A1_t (new_AGEMA_signal_10257), .A1_f (new_AGEMA_signal_10258), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .B0_f (new_AGEMA_signal_6216), .B1_t (new_AGEMA_signal_6217), .B1_f (new_AGEMA_signal_6218), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63), .Z0_f (new_AGEMA_signal_11000), .Z1_t (new_AGEMA_signal_11001), .Z1_f (new_AGEMA_signal_11002) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .A0_f (new_AGEMA_signal_10997), .A1_t (new_AGEMA_signal_10998), .A1_f (new_AGEMA_signal_10999), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62), .B0_f (new_AGEMA_signal_11699), .B1_t (new_AGEMA_signal_11700), .B1_f (new_AGEMA_signal_11701), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .Z0_f (new_AGEMA_signal_12296), .Z1_t (new_AGEMA_signal_12297), .Z1_f (new_AGEMA_signal_12298) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50), .A0_f (new_AGEMA_signal_10274), .A1_t (new_AGEMA_signal_10275), .A1_f (new_AGEMA_signal_10276), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56), .B0_f (new_AGEMA_signal_10280), .B1_t (new_AGEMA_signal_10281), .B1_f (new_AGEMA_signal_10282), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .Z0_f (new_AGEMA_signal_11003), .Z1_t (new_AGEMA_signal_11004), .Z1_f (new_AGEMA_signal_11005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46), .A0_f (new_AGEMA_signal_10979), .A1_t (new_AGEMA_signal_10980), .A1_f (new_AGEMA_signal_10981), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48), .B0_f (new_AGEMA_signal_10271), .B1_t (new_AGEMA_signal_10272), .B1_f (new_AGEMA_signal_10273), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2), .Z0_f (new_AGEMA_signal_11702), .Z1_t (new_AGEMA_signal_11703), .Z1_f (new_AGEMA_signal_11704) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47), .A0_f (new_AGEMA_signal_10268), .A1_t (new_AGEMA_signal_10269), .A1_f (new_AGEMA_signal_10270), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55), .B0_f (new_AGEMA_signal_10991), .B1_t (new_AGEMA_signal_10992), .B1_f (new_AGEMA_signal_10993), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3), .Z0_f (new_AGEMA_signal_11705), .Z1_t (new_AGEMA_signal_11706), .Z1_f (new_AGEMA_signal_11707) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54), .A0_f (new_AGEMA_signal_10988), .A1_t (new_AGEMA_signal_10989), .A1_f (new_AGEMA_signal_10990), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58), .B0_f (new_AGEMA_signal_10994), .B1_t (new_AGEMA_signal_10995), .B1_f (new_AGEMA_signal_10996), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4), .Z0_f (new_AGEMA_signal_11708), .Z1_t (new_AGEMA_signal_11709), .Z1_f (new_AGEMA_signal_11710) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49), .A0_f (new_AGEMA_signal_10982), .A1_t (new_AGEMA_signal_10983), .A1_f (new_AGEMA_signal_10984), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .B0_f (new_AGEMA_signal_10997), .B1_t (new_AGEMA_signal_10998), .B1_f (new_AGEMA_signal_10999), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5), .Z0_f (new_AGEMA_signal_11711), .Z1_t (new_AGEMA_signal_11712), .Z1_f (new_AGEMA_signal_11713) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62), .A0_f (new_AGEMA_signal_11699), .A1_t (new_AGEMA_signal_11700), .A1_f (new_AGEMA_signal_11701), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5), .B0_f (new_AGEMA_signal_11711), .B1_t (new_AGEMA_signal_11712), .B1_f (new_AGEMA_signal_11713), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .Z0_f (new_AGEMA_signal_12299), .Z1_t (new_AGEMA_signal_12300), .Z1_f (new_AGEMA_signal_12301) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46), .A0_f (new_AGEMA_signal_10979), .A1_t (new_AGEMA_signal_10980), .A1_f (new_AGEMA_signal_10981), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3), .B0_f (new_AGEMA_signal_11705), .B1_t (new_AGEMA_signal_11706), .B1_f (new_AGEMA_signal_11707), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7), .Z0_f (new_AGEMA_signal_12302), .Z1_t (new_AGEMA_signal_12303), .Z1_f (new_AGEMA_signal_12304) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51), .A0_f (new_AGEMA_signal_10277), .A1_t (new_AGEMA_signal_10278), .A1_f (new_AGEMA_signal_10279), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59), .B0_f (new_AGEMA_signal_10286), .B1_t (new_AGEMA_signal_10287), .B1_f (new_AGEMA_signal_10288), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8), .Z0_f (new_AGEMA_signal_11006), .Z1_t (new_AGEMA_signal_11007), .Z1_f (new_AGEMA_signal_11008) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52), .A0_f (new_AGEMA_signal_10985), .A1_t (new_AGEMA_signal_10986), .A1_f (new_AGEMA_signal_10987), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53), .B0_f (new_AGEMA_signal_11696), .B1_t (new_AGEMA_signal_11697), .B1_f (new_AGEMA_signal_11698), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9), .Z0_f (new_AGEMA_signal_12305), .Z1_t (new_AGEMA_signal_12306), .Z1_f (new_AGEMA_signal_12307) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53), .A0_f (new_AGEMA_signal_11696), .A1_t (new_AGEMA_signal_11697), .A1_f (new_AGEMA_signal_11698), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4), .B0_f (new_AGEMA_signal_11708), .B1_t (new_AGEMA_signal_11709), .B1_f (new_AGEMA_signal_11710), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10), .Z0_f (new_AGEMA_signal_12308), .Z1_t (new_AGEMA_signal_12309), .Z1_f (new_AGEMA_signal_12310) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60), .A0_f (new_AGEMA_signal_10289), .A1_t (new_AGEMA_signal_10290), .A1_f (new_AGEMA_signal_10291), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2), .B0_f (new_AGEMA_signal_11702), .B1_t (new_AGEMA_signal_11703), .B1_f (new_AGEMA_signal_11704), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11), .Z0_f (new_AGEMA_signal_12311), .Z1_t (new_AGEMA_signal_12312), .Z1_f (new_AGEMA_signal_12313) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48), .A0_f (new_AGEMA_signal_10271), .A1_t (new_AGEMA_signal_10272), .A1_f (new_AGEMA_signal_10273), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51), .B0_f (new_AGEMA_signal_10277), .B1_t (new_AGEMA_signal_10278), .B1_f (new_AGEMA_signal_10279), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12), .Z0_f (new_AGEMA_signal_11009), .Z1_t (new_AGEMA_signal_11010), .Z1_f (new_AGEMA_signal_11011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50), .A0_f (new_AGEMA_signal_10274), .A1_t (new_AGEMA_signal_10275), .A1_f (new_AGEMA_signal_10276), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .B0_f (new_AGEMA_signal_12296), .B1_t (new_AGEMA_signal_12297), .B1_f (new_AGEMA_signal_12298), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13), .Z0_f (new_AGEMA_signal_12836), .Z1_t (new_AGEMA_signal_12837), .Z1_f (new_AGEMA_signal_12838) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52), .A0_f (new_AGEMA_signal_10985), .A1_t (new_AGEMA_signal_10986), .A1_f (new_AGEMA_signal_10987), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .B0_f (new_AGEMA_signal_10997), .B1_t (new_AGEMA_signal_10998), .B1_f (new_AGEMA_signal_10999), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14), .Z0_f (new_AGEMA_signal_11714), .Z1_t (new_AGEMA_signal_11715), .Z1_f (new_AGEMA_signal_11716) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55), .A0_f (new_AGEMA_signal_10991), .A1_t (new_AGEMA_signal_10992), .A1_f (new_AGEMA_signal_10993), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .B0_f (new_AGEMA_signal_11003), .B1_t (new_AGEMA_signal_11004), .B1_f (new_AGEMA_signal_11005), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15), .Z0_f (new_AGEMA_signal_11717), .Z1_t (new_AGEMA_signal_11718), .Z1_f (new_AGEMA_signal_11719) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56), .A0_f (new_AGEMA_signal_10280), .A1_t (new_AGEMA_signal_10281), .A1_f (new_AGEMA_signal_10282), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .B0_f (new_AGEMA_signal_12296), .B1_t (new_AGEMA_signal_12297), .B1_f (new_AGEMA_signal_12298), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16), .Z0_f (new_AGEMA_signal_12839), .Z1_t (new_AGEMA_signal_12840), .Z1_f (new_AGEMA_signal_12841) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57), .A0_f (new_AGEMA_signal_10283), .A1_t (new_AGEMA_signal_10284), .A1_f (new_AGEMA_signal_10285), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .B0_f (new_AGEMA_signal_11003), .B1_t (new_AGEMA_signal_11004), .B1_f (new_AGEMA_signal_11005), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17), .Z0_f (new_AGEMA_signal_11720), .Z1_t (new_AGEMA_signal_11721), .Z1_f (new_AGEMA_signal_11722) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58), .A0_f (new_AGEMA_signal_10994), .A1_t (new_AGEMA_signal_10995), .A1_f (new_AGEMA_signal_10996), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8), .B0_f (new_AGEMA_signal_11006), .B1_t (new_AGEMA_signal_11007), .B1_f (new_AGEMA_signal_11008), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18), .Z0_f (new_AGEMA_signal_11723), .Z1_t (new_AGEMA_signal_11724), .Z1_f (new_AGEMA_signal_11725) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63), .A0_f (new_AGEMA_signal_11000), .A1_t (new_AGEMA_signal_11001), .A1_f (new_AGEMA_signal_11002), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4), .B0_f (new_AGEMA_signal_11708), .B1_t (new_AGEMA_signal_11709), .B1_f (new_AGEMA_signal_11710), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19), .Z0_f (new_AGEMA_signal_12314), .Z1_t (new_AGEMA_signal_12315), .Z1_f (new_AGEMA_signal_12316) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .A0_f (new_AGEMA_signal_12296), .A1_t (new_AGEMA_signal_12297), .A1_f (new_AGEMA_signal_12298), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .B0_f (new_AGEMA_signal_11003), .B1_t (new_AGEMA_signal_11004), .B1_f (new_AGEMA_signal_11005), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20), .Z0_f (new_AGEMA_signal_12842), .Z1_t (new_AGEMA_signal_12843), .Z1_f (new_AGEMA_signal_12844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .A0_f (new_AGEMA_signal_11003), .A1_t (new_AGEMA_signal_11004), .A1_f (new_AGEMA_signal_11005), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7), .B0_f (new_AGEMA_signal_12302), .B1_t (new_AGEMA_signal_12303), .B1_f (new_AGEMA_signal_12304), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21), .Z0_f (new_AGEMA_signal_12845), .Z1_t (new_AGEMA_signal_12846), .Z1_f (new_AGEMA_signal_12847) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3), .A0_f (new_AGEMA_signal_11705), .A1_t (new_AGEMA_signal_11706), .A1_f (new_AGEMA_signal_11707), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12), .B0_f (new_AGEMA_signal_11009), .B1_t (new_AGEMA_signal_11010), .B1_f (new_AGEMA_signal_11011), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22), .Z0_f (new_AGEMA_signal_12317), .Z1_t (new_AGEMA_signal_12318), .Z1_f (new_AGEMA_signal_12319) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18), .A0_f (new_AGEMA_signal_11723), .A1_t (new_AGEMA_signal_11724), .A1_f (new_AGEMA_signal_11725), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2), .B0_f (new_AGEMA_signal_11702), .B1_t (new_AGEMA_signal_11703), .B1_f (new_AGEMA_signal_11704), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23), .Z0_f (new_AGEMA_signal_12320), .Z1_t (new_AGEMA_signal_12321), .Z1_f (new_AGEMA_signal_12322) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15), .A0_f (new_AGEMA_signal_11717), .A1_t (new_AGEMA_signal_11718), .A1_f (new_AGEMA_signal_11719), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9), .B0_f (new_AGEMA_signal_12305), .B1_t (new_AGEMA_signal_12306), .B1_f (new_AGEMA_signal_12307), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24), .Z0_f (new_AGEMA_signal_12848), .Z1_t (new_AGEMA_signal_12849), .Z1_f (new_AGEMA_signal_12850) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .A0_f (new_AGEMA_signal_12299), .A1_t (new_AGEMA_signal_12300), .A1_f (new_AGEMA_signal_12301), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10), .B0_f (new_AGEMA_signal_12308), .B1_t (new_AGEMA_signal_12309), .B1_f (new_AGEMA_signal_12310), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25), .Z0_f (new_AGEMA_signal_12851), .Z1_t (new_AGEMA_signal_12852), .Z1_f (new_AGEMA_signal_12853) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7), .A0_f (new_AGEMA_signal_12302), .A1_t (new_AGEMA_signal_12303), .A1_f (new_AGEMA_signal_12304), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9), .B0_f (new_AGEMA_signal_12305), .B1_t (new_AGEMA_signal_12306), .B1_f (new_AGEMA_signal_12307), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26), .Z0_f (new_AGEMA_signal_12854), .Z1_t (new_AGEMA_signal_12855), .Z1_f (new_AGEMA_signal_12856) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8), .A0_f (new_AGEMA_signal_11006), .A1_t (new_AGEMA_signal_11007), .A1_f (new_AGEMA_signal_11008), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10), .B0_f (new_AGEMA_signal_12308), .B1_t (new_AGEMA_signal_12309), .B1_f (new_AGEMA_signal_12310), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27), .Z0_f (new_AGEMA_signal_12857), .Z1_t (new_AGEMA_signal_12858), .Z1_f (new_AGEMA_signal_12859) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11), .A0_f (new_AGEMA_signal_12311), .A1_t (new_AGEMA_signal_12312), .A1_f (new_AGEMA_signal_12313), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14), .B0_f (new_AGEMA_signal_11714), .B1_t (new_AGEMA_signal_11715), .B1_f (new_AGEMA_signal_11716), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28), .Z0_f (new_AGEMA_signal_12860), .Z1_t (new_AGEMA_signal_12861), .Z1_f (new_AGEMA_signal_12862) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11), .A0_f (new_AGEMA_signal_12311), .A1_t (new_AGEMA_signal_12312), .A1_f (new_AGEMA_signal_12313), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17), .B0_f (new_AGEMA_signal_11720), .B1_t (new_AGEMA_signal_11721), .B1_f (new_AGEMA_signal_11722), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29), .Z0_f (new_AGEMA_signal_12863), .Z1_t (new_AGEMA_signal_12864), .Z1_f (new_AGEMA_signal_12865) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .A0_f (new_AGEMA_signal_12299), .A1_t (new_AGEMA_signal_12300), .A1_f (new_AGEMA_signal_12301), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24), .B0_f (new_AGEMA_signal_12848), .B1_t (new_AGEMA_signal_12849), .B1_f (new_AGEMA_signal_12850), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_), .Z0_f (new_AGEMA_signal_13508), .Z1_t (new_AGEMA_signal_13509), .Z1_f (new_AGEMA_signal_13510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16), .A0_f (new_AGEMA_signal_12839), .A1_t (new_AGEMA_signal_12840), .A1_f (new_AGEMA_signal_12841), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26), .B0_f (new_AGEMA_signal_12854), .B1_t (new_AGEMA_signal_12855), .B1_f (new_AGEMA_signal_12856), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_), .Z0_f (new_AGEMA_signal_13511), .Z1_t (new_AGEMA_signal_13512), .Z1_f (new_AGEMA_signal_13513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19), .A0_f (new_AGEMA_signal_12314), .A1_t (new_AGEMA_signal_12315), .A1_f (new_AGEMA_signal_12316), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28), .B0_f (new_AGEMA_signal_12860), .B1_t (new_AGEMA_signal_12861), .B1_f (new_AGEMA_signal_12862), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_), .Z0_f (new_AGEMA_signal_13514), .Z1_t (new_AGEMA_signal_13515), .Z1_f (new_AGEMA_signal_13516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .A0_f (new_AGEMA_signal_12299), .A1_t (new_AGEMA_signal_12300), .A1_f (new_AGEMA_signal_12301), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21), .B0_f (new_AGEMA_signal_12845), .B1_t (new_AGEMA_signal_12846), .B1_f (new_AGEMA_signal_12847), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_), .Z0_f (new_AGEMA_signal_13517), .Z1_t (new_AGEMA_signal_13518), .Z1_f (new_AGEMA_signal_13519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20), .A0_f (new_AGEMA_signal_12842), .A1_t (new_AGEMA_signal_12843), .A1_f (new_AGEMA_signal_12844), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22), .B0_f (new_AGEMA_signal_12317), .B1_t (new_AGEMA_signal_12318), .B1_f (new_AGEMA_signal_12319), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_), .Z0_f (new_AGEMA_signal_13520), .Z1_t (new_AGEMA_signal_13521), .Z1_f (new_AGEMA_signal_13522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25), .A0_f (new_AGEMA_signal_12851), .A1_t (new_AGEMA_signal_12852), .A1_f (new_AGEMA_signal_12853), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29), .B0_f (new_AGEMA_signal_12863), .B1_t (new_AGEMA_signal_12864), .B1_f (new_AGEMA_signal_12865), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_), .Z0_f (new_AGEMA_signal_13523), .Z1_t (new_AGEMA_signal_13524), .Z1_f (new_AGEMA_signal_13525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13), .A0_f (new_AGEMA_signal_12836), .A1_t (new_AGEMA_signal_12837), .A1_f (new_AGEMA_signal_12838), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27), .B0_f (new_AGEMA_signal_12857), .B1_t (new_AGEMA_signal_12858), .B1_f (new_AGEMA_signal_12859), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_), .Z0_f (new_AGEMA_signal_13526), .Z1_t (new_AGEMA_signal_13527), .Z1_f (new_AGEMA_signal_13528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .A0_f (new_AGEMA_signal_12299), .A1_t (new_AGEMA_signal_12300), .A1_f (new_AGEMA_signal_12301), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23), .B0_f (new_AGEMA_signal_12320), .B1_t (new_AGEMA_signal_12321), .B1_f (new_AGEMA_signal_12322), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_), .Z0_f (new_AGEMA_signal_12866), .Z1_t (new_AGEMA_signal_12867), .Z1_f (new_AGEMA_signal_12868) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T1_U1 ( .A0_t (RoundKey[15]), .A0_f (new_AGEMA_signal_5369), .A1_t (new_AGEMA_signal_5370), .A1_f (new_AGEMA_signal_5371), .B0_t (RoundKey[12]), .B0_f (new_AGEMA_signal_5342), .B1_t (new_AGEMA_signal_5343), .B1_f (new_AGEMA_signal_5344), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .Z0_f (new_AGEMA_signal_6243), .Z1_t (new_AGEMA_signal_6244), .Z1_f (new_AGEMA_signal_6245) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T2_U1 ( .A0_t (RoundKey[15]), .A0_f (new_AGEMA_signal_5369), .A1_t (new_AGEMA_signal_5370), .A1_f (new_AGEMA_signal_5371), .B0_t (RoundKey[10]), .B0_f (new_AGEMA_signal_5162), .B1_t (new_AGEMA_signal_5163), .B1_f (new_AGEMA_signal_5164), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .Z0_f (new_AGEMA_signal_6246), .Z1_t (new_AGEMA_signal_6247), .Z1_f (new_AGEMA_signal_6248) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T3_U1 ( .A0_t (RoundKey[15]), .A0_f (new_AGEMA_signal_5369), .A1_t (new_AGEMA_signal_5370), .A1_f (new_AGEMA_signal_5371), .B0_t (RoundKey[9]), .B0_f (new_AGEMA_signal_6206), .B1_t (new_AGEMA_signal_6207), .B1_f (new_AGEMA_signal_6208), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .Z0_f (new_AGEMA_signal_6249), .Z1_t (new_AGEMA_signal_6250), .Z1_f (new_AGEMA_signal_6251) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T4_U1 ( .A0_t (RoundKey[12]), .A0_f (new_AGEMA_signal_5342), .A1_t (new_AGEMA_signal_5343), .A1_f (new_AGEMA_signal_5344), .B0_t (RoundKey[10]), .B0_f (new_AGEMA_signal_5162), .B1_t (new_AGEMA_signal_5163), .B1_f (new_AGEMA_signal_5164), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .Z0_f (new_AGEMA_signal_6252), .Z1_t (new_AGEMA_signal_6253), .Z1_f (new_AGEMA_signal_6254) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T5_U1 ( .A0_t (RoundKey[11]), .A0_f (new_AGEMA_signal_5261), .A1_t (new_AGEMA_signal_5262), .A1_f (new_AGEMA_signal_5263), .B0_t (RoundKey[9]), .B0_f (new_AGEMA_signal_6206), .B1_t (new_AGEMA_signal_6207), .B1_f (new_AGEMA_signal_6208), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .Z0_f (new_AGEMA_signal_6255), .Z1_t (new_AGEMA_signal_6256), .Z1_f (new_AGEMA_signal_6257) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .A0_f (new_AGEMA_signal_6243), .A1_t (new_AGEMA_signal_6244), .A1_f (new_AGEMA_signal_6245), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .B0_f (new_AGEMA_signal_6255), .B1_t (new_AGEMA_signal_6256), .B1_f (new_AGEMA_signal_6257), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .Z0_f (new_AGEMA_signal_6850), .Z1_t (new_AGEMA_signal_6851), .Z1_f (new_AGEMA_signal_6852) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T7_U1 ( .A0_t (RoundKey[14]), .A0_f (new_AGEMA_signal_5360), .A1_t (new_AGEMA_signal_5361), .A1_f (new_AGEMA_signal_5362), .B0_t (RoundKey[13]), .B0_f (new_AGEMA_signal_5351), .B1_t (new_AGEMA_signal_5352), .B1_f (new_AGEMA_signal_5353), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .Z0_f (new_AGEMA_signal_6258), .Z1_t (new_AGEMA_signal_6259), .Z1_f (new_AGEMA_signal_6260) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T8_U1 ( .A0_t (RoundKey[8]), .A0_f (new_AGEMA_signal_6107), .A1_t (new_AGEMA_signal_6108), .A1_f (new_AGEMA_signal_6109), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .B0_f (new_AGEMA_signal_6850), .B1_t (new_AGEMA_signal_6851), .B1_f (new_AGEMA_signal_6852), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .Z0_f (new_AGEMA_signal_7351), .Z1_t (new_AGEMA_signal_7352), .Z1_f (new_AGEMA_signal_7353) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T9_U1 ( .A0_t (RoundKey[8]), .A0_f (new_AGEMA_signal_6107), .A1_t (new_AGEMA_signal_6108), .A1_f (new_AGEMA_signal_6109), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .B0_f (new_AGEMA_signal_6258), .B1_t (new_AGEMA_signal_6259), .B1_f (new_AGEMA_signal_6260), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .Z0_f (new_AGEMA_signal_6853), .Z1_t (new_AGEMA_signal_6854), .Z1_f (new_AGEMA_signal_6855) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .A0_f (new_AGEMA_signal_6850), .A1_t (new_AGEMA_signal_6851), .A1_f (new_AGEMA_signal_6852), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .B0_f (new_AGEMA_signal_6258), .B1_t (new_AGEMA_signal_6259), .B1_f (new_AGEMA_signal_6260), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .Z0_f (new_AGEMA_signal_7354), .Z1_t (new_AGEMA_signal_7355), .Z1_f (new_AGEMA_signal_7356) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T11_U1 ( .A0_t (RoundKey[14]), .A0_f (new_AGEMA_signal_5360), .A1_t (new_AGEMA_signal_5361), .A1_f (new_AGEMA_signal_5362), .B0_t (RoundKey[10]), .B0_f (new_AGEMA_signal_5162), .B1_t (new_AGEMA_signal_5163), .B1_f (new_AGEMA_signal_5164), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11), .Z0_f (new_AGEMA_signal_6261), .Z1_t (new_AGEMA_signal_6262), .Z1_f (new_AGEMA_signal_6263) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T12_U1 ( .A0_t (RoundKey[13]), .A0_f (new_AGEMA_signal_5351), .A1_t (new_AGEMA_signal_5352), .A1_f (new_AGEMA_signal_5353), .B0_t (RoundKey[10]), .B0_f (new_AGEMA_signal_5162), .B1_t (new_AGEMA_signal_5163), .B1_f (new_AGEMA_signal_5164), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12), .Z0_f (new_AGEMA_signal_6264), .Z1_t (new_AGEMA_signal_6265), .Z1_f (new_AGEMA_signal_6266) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .A0_f (new_AGEMA_signal_6249), .A1_t (new_AGEMA_signal_6250), .A1_f (new_AGEMA_signal_6251), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .B0_f (new_AGEMA_signal_6252), .B1_t (new_AGEMA_signal_6253), .B1_f (new_AGEMA_signal_6254), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .Z0_f (new_AGEMA_signal_6856), .Z1_t (new_AGEMA_signal_6857), .Z1_f (new_AGEMA_signal_6858) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .A0_f (new_AGEMA_signal_6850), .A1_t (new_AGEMA_signal_6851), .A1_f (new_AGEMA_signal_6852), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11), .B0_f (new_AGEMA_signal_6261), .B1_t (new_AGEMA_signal_6262), .B1_f (new_AGEMA_signal_6263), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14), .Z0_f (new_AGEMA_signal_7357), .Z1_t (new_AGEMA_signal_7358), .Z1_f (new_AGEMA_signal_7359) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .A0_f (new_AGEMA_signal_6255), .A1_t (new_AGEMA_signal_6256), .A1_f (new_AGEMA_signal_6257), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11), .B0_f (new_AGEMA_signal_6261), .B1_t (new_AGEMA_signal_6262), .B1_f (new_AGEMA_signal_6263), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .Z0_f (new_AGEMA_signal_6859), .Z1_t (new_AGEMA_signal_6860), .Z1_f (new_AGEMA_signal_6861) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .A0_f (new_AGEMA_signal_6255), .A1_t (new_AGEMA_signal_6256), .A1_f (new_AGEMA_signal_6257), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12), .B0_f (new_AGEMA_signal_6264), .B1_t (new_AGEMA_signal_6265), .B1_f (new_AGEMA_signal_6266), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Z0_f (new_AGEMA_signal_6862), .Z1_t (new_AGEMA_signal_6863), .Z1_f (new_AGEMA_signal_6864) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .A0_f (new_AGEMA_signal_6853), .A1_t (new_AGEMA_signal_6854), .A1_f (new_AGEMA_signal_6855), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .B0_f (new_AGEMA_signal_6862), .B1_t (new_AGEMA_signal_6863), .B1_f (new_AGEMA_signal_6864), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .Z0_f (new_AGEMA_signal_7360), .Z1_t (new_AGEMA_signal_7361), .Z1_f (new_AGEMA_signal_7362) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T18_U1 ( .A0_t (RoundKey[12]), .A0_f (new_AGEMA_signal_5342), .A1_t (new_AGEMA_signal_5343), .A1_f (new_AGEMA_signal_5344), .B0_t (RoundKey[8]), .B0_f (new_AGEMA_signal_6107), .B1_t (new_AGEMA_signal_6108), .B1_f (new_AGEMA_signal_6109), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18), .Z0_f (new_AGEMA_signal_6267), .Z1_t (new_AGEMA_signal_6268), .Z1_f (new_AGEMA_signal_6269) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .A0_f (new_AGEMA_signal_6258), .A1_t (new_AGEMA_signal_6259), .A1_f (new_AGEMA_signal_6260), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18), .B0_f (new_AGEMA_signal_6267), .B1_t (new_AGEMA_signal_6268), .B1_f (new_AGEMA_signal_6269), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .Z0_f (new_AGEMA_signal_6865), .Z1_t (new_AGEMA_signal_6866), .Z1_f (new_AGEMA_signal_6867) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .A0_f (new_AGEMA_signal_6243), .A1_t (new_AGEMA_signal_6244), .A1_f (new_AGEMA_signal_6245), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .B0_f (new_AGEMA_signal_6865), .B1_t (new_AGEMA_signal_6866), .B1_f (new_AGEMA_signal_6867), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .Z0_f (new_AGEMA_signal_7363), .Z1_t (new_AGEMA_signal_7364), .Z1_f (new_AGEMA_signal_7365) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T21_U1 ( .A0_t (RoundKey[9]), .A0_f (new_AGEMA_signal_6206), .A1_t (new_AGEMA_signal_6207), .A1_f (new_AGEMA_signal_6208), .B0_t (RoundKey[8]), .B0_f (new_AGEMA_signal_6107), .B1_t (new_AGEMA_signal_6108), .B1_f (new_AGEMA_signal_6109), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21), .Z0_f (new_AGEMA_signal_6270), .Z1_t (new_AGEMA_signal_6271), .Z1_f (new_AGEMA_signal_6272) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .A0_f (new_AGEMA_signal_6258), .A1_t (new_AGEMA_signal_6259), .A1_f (new_AGEMA_signal_6260), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21), .B0_f (new_AGEMA_signal_6270), .B1_t (new_AGEMA_signal_6271), .B1_f (new_AGEMA_signal_6272), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .Z0_f (new_AGEMA_signal_6868), .Z1_t (new_AGEMA_signal_6869), .Z1_f (new_AGEMA_signal_6870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .A0_f (new_AGEMA_signal_6246), .A1_t (new_AGEMA_signal_6247), .A1_f (new_AGEMA_signal_6248), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .B0_f (new_AGEMA_signal_6868), .B1_t (new_AGEMA_signal_6869), .B1_f (new_AGEMA_signal_6870), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .Z0_f (new_AGEMA_signal_7366), .Z1_t (new_AGEMA_signal_7367), .Z1_f (new_AGEMA_signal_7368) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .A0_f (new_AGEMA_signal_6246), .A1_t (new_AGEMA_signal_6247), .A1_f (new_AGEMA_signal_6248), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .B0_f (new_AGEMA_signal_7354), .B1_t (new_AGEMA_signal_7355), .B1_f (new_AGEMA_signal_7356), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24), .Z0_f (new_AGEMA_signal_8123), .Z1_t (new_AGEMA_signal_8124), .Z1_f (new_AGEMA_signal_8125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .A0_f (new_AGEMA_signal_7363), .A1_t (new_AGEMA_signal_7364), .A1_f (new_AGEMA_signal_7365), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .B0_f (new_AGEMA_signal_7360), .B1_t (new_AGEMA_signal_7361), .B1_f (new_AGEMA_signal_7362), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25), .Z0_f (new_AGEMA_signal_8126), .Z1_t (new_AGEMA_signal_8127), .Z1_f (new_AGEMA_signal_8128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .A0_f (new_AGEMA_signal_6249), .A1_t (new_AGEMA_signal_6250), .A1_f (new_AGEMA_signal_6251), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .B0_f (new_AGEMA_signal_6862), .B1_t (new_AGEMA_signal_6863), .B1_f (new_AGEMA_signal_6864), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26), .Z0_f (new_AGEMA_signal_7369), .Z1_t (new_AGEMA_signal_7370), .Z1_f (new_AGEMA_signal_7371) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .A0_f (new_AGEMA_signal_6243), .A1_t (new_AGEMA_signal_6244), .A1_f (new_AGEMA_signal_6245), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12), .B0_f (new_AGEMA_signal_6264), .B1_t (new_AGEMA_signal_6265), .B1_f (new_AGEMA_signal_6266), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .Z0_f (new_AGEMA_signal_6871), .Z1_t (new_AGEMA_signal_6872), .Z1_f (new_AGEMA_signal_6873) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .A0_f (new_AGEMA_signal_6856), .A1_t (new_AGEMA_signal_6857), .A1_f (new_AGEMA_signal_6858), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .B0_f (new_AGEMA_signal_6850), .B1_t (new_AGEMA_signal_6851), .B1_f (new_AGEMA_signal_6852), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1), .Z0_f (new_AGEMA_signal_7372), .Z1_t (new_AGEMA_signal_7373), .Z1_f (new_AGEMA_signal_7374) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .A0_f (new_AGEMA_signal_7366), .A1_t (new_AGEMA_signal_7367), .A1_f (new_AGEMA_signal_7368), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .B0_f (new_AGEMA_signal_7351), .B1_t (new_AGEMA_signal_7352), .B1_f (new_AGEMA_signal_7353), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2), .Z0_f (new_AGEMA_signal_8129), .Z1_t (new_AGEMA_signal_8130), .Z1_f (new_AGEMA_signal_8131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14), .A0_f (new_AGEMA_signal_7357), .A1_t (new_AGEMA_signal_7358), .A1_f (new_AGEMA_signal_7359), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1), .B0_f (new_AGEMA_signal_7372), .B1_t (new_AGEMA_signal_7373), .B1_f (new_AGEMA_signal_7374), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3), .Z0_f (new_AGEMA_signal_8132), .Z1_t (new_AGEMA_signal_8133), .Z1_f (new_AGEMA_signal_8134) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .A0_f (new_AGEMA_signal_6865), .A1_t (new_AGEMA_signal_6866), .A1_f (new_AGEMA_signal_6867), .B0_t (RoundKey[8]), .B0_f (new_AGEMA_signal_6107), .B1_t (new_AGEMA_signal_6108), .B1_f (new_AGEMA_signal_6109), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4), .Z0_f (new_AGEMA_signal_7375), .Z1_t (new_AGEMA_signal_7376), .Z1_f (new_AGEMA_signal_7377) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4), .A0_f (new_AGEMA_signal_7375), .A1_t (new_AGEMA_signal_7376), .A1_f (new_AGEMA_signal_7377), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1), .B0_f (new_AGEMA_signal_7372), .B1_t (new_AGEMA_signal_7373), .B1_f (new_AGEMA_signal_7374), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5), .Z0_f (new_AGEMA_signal_8135), .Z1_t (new_AGEMA_signal_8136), .Z1_f (new_AGEMA_signal_8137) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .A0_f (new_AGEMA_signal_6249), .A1_t (new_AGEMA_signal_6250), .A1_f (new_AGEMA_signal_6251), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .B0_f (new_AGEMA_signal_6862), .B1_t (new_AGEMA_signal_6863), .B1_f (new_AGEMA_signal_6864), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6), .Z0_f (new_AGEMA_signal_7378), .Z1_t (new_AGEMA_signal_7379), .Z1_f (new_AGEMA_signal_7380) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .A0_f (new_AGEMA_signal_6868), .A1_t (new_AGEMA_signal_6869), .A1_f (new_AGEMA_signal_6870), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .B0_f (new_AGEMA_signal_6853), .B1_t (new_AGEMA_signal_6854), .B1_f (new_AGEMA_signal_6855), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7), .Z0_f (new_AGEMA_signal_7381), .Z1_t (new_AGEMA_signal_7382), .Z1_f (new_AGEMA_signal_7383) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26), .A0_f (new_AGEMA_signal_7369), .A1_t (new_AGEMA_signal_7370), .A1_f (new_AGEMA_signal_7371), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6), .B0_f (new_AGEMA_signal_7378), .B1_t (new_AGEMA_signal_7379), .B1_f (new_AGEMA_signal_7380), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8), .Z0_f (new_AGEMA_signal_8138), .Z1_t (new_AGEMA_signal_8139), .Z1_f (new_AGEMA_signal_8140) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .A0_f (new_AGEMA_signal_7363), .A1_t (new_AGEMA_signal_7364), .A1_f (new_AGEMA_signal_7365), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .B0_f (new_AGEMA_signal_7360), .B1_t (new_AGEMA_signal_7361), .B1_f (new_AGEMA_signal_7362), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9), .Z0_f (new_AGEMA_signal_8141), .Z1_t (new_AGEMA_signal_8142), .Z1_f (new_AGEMA_signal_8143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9), .A0_f (new_AGEMA_signal_8141), .A1_t (new_AGEMA_signal_8142), .A1_f (new_AGEMA_signal_8143), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6), .B0_f (new_AGEMA_signal_7378), .B1_t (new_AGEMA_signal_7379), .B1_f (new_AGEMA_signal_7380), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10), .Z0_f (new_AGEMA_signal_8651), .Z1_t (new_AGEMA_signal_8652), .Z1_f (new_AGEMA_signal_8653) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .A0_f (new_AGEMA_signal_6243), .A1_t (new_AGEMA_signal_6244), .A1_f (new_AGEMA_signal_6245), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .B0_f (new_AGEMA_signal_6859), .B1_t (new_AGEMA_signal_6860), .B1_f (new_AGEMA_signal_6861), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11), .Z0_f (new_AGEMA_signal_7384), .Z1_t (new_AGEMA_signal_7385), .Z1_f (new_AGEMA_signal_7386) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .A0_f (new_AGEMA_signal_6252), .A1_t (new_AGEMA_signal_6253), .A1_f (new_AGEMA_signal_6254), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .B0_f (new_AGEMA_signal_6871), .B1_t (new_AGEMA_signal_6872), .B1_f (new_AGEMA_signal_6873), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12), .Z0_f (new_AGEMA_signal_7387), .Z1_t (new_AGEMA_signal_7388), .Z1_f (new_AGEMA_signal_7389) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12), .A0_f (new_AGEMA_signal_7387), .A1_t (new_AGEMA_signal_7388), .A1_f (new_AGEMA_signal_7389), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11), .B0_f (new_AGEMA_signal_7384), .B1_t (new_AGEMA_signal_7385), .B1_f (new_AGEMA_signal_7386), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13), .Z0_f (new_AGEMA_signal_8144), .Z1_t (new_AGEMA_signal_8145), .Z1_f (new_AGEMA_signal_8146) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .A0_f (new_AGEMA_signal_6246), .A1_t (new_AGEMA_signal_6247), .A1_f (new_AGEMA_signal_6248), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .B0_f (new_AGEMA_signal_7354), .B1_t (new_AGEMA_signal_7355), .B1_f (new_AGEMA_signal_7356), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14), .Z0_f (new_AGEMA_signal_8147), .Z1_t (new_AGEMA_signal_8148), .Z1_f (new_AGEMA_signal_8149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14), .A0_f (new_AGEMA_signal_8147), .A1_t (new_AGEMA_signal_8148), .A1_f (new_AGEMA_signal_8149), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11), .B0_f (new_AGEMA_signal_7384), .B1_t (new_AGEMA_signal_7385), .B1_f (new_AGEMA_signal_7386), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15), .Z0_f (new_AGEMA_signal_8654), .Z1_t (new_AGEMA_signal_8655), .Z1_f (new_AGEMA_signal_8656) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3), .A0_f (new_AGEMA_signal_8132), .A1_t (new_AGEMA_signal_8133), .A1_f (new_AGEMA_signal_8134), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2), .B0_f (new_AGEMA_signal_8129), .B1_t (new_AGEMA_signal_8130), .B1_f (new_AGEMA_signal_8131), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16), .Z0_f (new_AGEMA_signal_8657), .Z1_t (new_AGEMA_signal_8658), .Z1_f (new_AGEMA_signal_8659) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5), .A0_f (new_AGEMA_signal_8135), .A1_t (new_AGEMA_signal_8136), .A1_f (new_AGEMA_signal_8137), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24), .B0_f (new_AGEMA_signal_8123), .B1_t (new_AGEMA_signal_8124), .B1_f (new_AGEMA_signal_8125), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17), .Z0_f (new_AGEMA_signal_8660), .Z1_t (new_AGEMA_signal_8661), .Z1_f (new_AGEMA_signal_8662) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8), .A0_f (new_AGEMA_signal_8138), .A1_t (new_AGEMA_signal_8139), .A1_f (new_AGEMA_signal_8140), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7), .B0_f (new_AGEMA_signal_7381), .B1_t (new_AGEMA_signal_7382), .B1_f (new_AGEMA_signal_7383), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18), .Z0_f (new_AGEMA_signal_8663), .Z1_t (new_AGEMA_signal_8664), .Z1_f (new_AGEMA_signal_8665) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10), .A0_f (new_AGEMA_signal_8651), .A1_t (new_AGEMA_signal_8652), .A1_f (new_AGEMA_signal_8653), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15), .B0_f (new_AGEMA_signal_8654), .B1_t (new_AGEMA_signal_8655), .B1_f (new_AGEMA_signal_8656), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19), .Z0_f (new_AGEMA_signal_8948), .Z1_t (new_AGEMA_signal_8949), .Z1_f (new_AGEMA_signal_8950) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16), .A0_f (new_AGEMA_signal_8657), .A1_t (new_AGEMA_signal_8658), .A1_f (new_AGEMA_signal_8659), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13), .B0_f (new_AGEMA_signal_8144), .B1_t (new_AGEMA_signal_8145), .B1_f (new_AGEMA_signal_8146), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .Z0_f (new_AGEMA_signal_8951), .Z1_t (new_AGEMA_signal_8952), .Z1_f (new_AGEMA_signal_8953) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17), .A0_f (new_AGEMA_signal_8660), .A1_t (new_AGEMA_signal_8661), .A1_f (new_AGEMA_signal_8662), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15), .B0_f (new_AGEMA_signal_8654), .B1_t (new_AGEMA_signal_8655), .B1_f (new_AGEMA_signal_8656), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .Z0_f (new_AGEMA_signal_8954), .Z1_t (new_AGEMA_signal_8955), .Z1_f (new_AGEMA_signal_8956) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18), .A0_f (new_AGEMA_signal_8663), .A1_t (new_AGEMA_signal_8664), .A1_f (new_AGEMA_signal_8665), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13), .B0_f (new_AGEMA_signal_8144), .B1_t (new_AGEMA_signal_8145), .B1_f (new_AGEMA_signal_8146), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .Z0_f (new_AGEMA_signal_8957), .Z1_t (new_AGEMA_signal_8958), .Z1_f (new_AGEMA_signal_8959) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19), .A0_f (new_AGEMA_signal_8948), .A1_t (new_AGEMA_signal_8949), .A1_f (new_AGEMA_signal_8950), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25), .B0_f (new_AGEMA_signal_8126), .B1_t (new_AGEMA_signal_8127), .B1_f (new_AGEMA_signal_8128), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .Z0_f (new_AGEMA_signal_9188), .Z1_t (new_AGEMA_signal_9189), .Z1_f (new_AGEMA_signal_9190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .A0_f (new_AGEMA_signal_8957), .A1_t (new_AGEMA_signal_8958), .A1_f (new_AGEMA_signal_8959), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .B0_f (new_AGEMA_signal_9188), .B1_t (new_AGEMA_signal_9189), .B1_f (new_AGEMA_signal_9190), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .Z0_f (new_AGEMA_signal_9431), .Z1_t (new_AGEMA_signal_9432), .Z1_f (new_AGEMA_signal_9433) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .A0_f (new_AGEMA_signal_8957), .A1_t (new_AGEMA_signal_8958), .A1_f (new_AGEMA_signal_8959), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .B0_f (new_AGEMA_signal_8951), .B1_t (new_AGEMA_signal_8952), .B1_f (new_AGEMA_signal_8953), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z0_f (new_AGEMA_signal_9191), .Z1_t (new_AGEMA_signal_9192), .Z1_f (new_AGEMA_signal_9193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .A0_f (new_AGEMA_signal_8954), .A1_t (new_AGEMA_signal_8955), .A1_f (new_AGEMA_signal_8956), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .B0_f (new_AGEMA_signal_9191), .B1_t (new_AGEMA_signal_9192), .B1_f (new_AGEMA_signal_9193), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26), .Z0_f (new_AGEMA_signal_9434), .Z1_t (new_AGEMA_signal_9435), .Z1_f (new_AGEMA_signal_9436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .A0_f (new_AGEMA_signal_8951), .A1_t (new_AGEMA_signal_8952), .A1_f (new_AGEMA_signal_8953), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .B0_f (new_AGEMA_signal_8954), .B1_t (new_AGEMA_signal_8955), .B1_f (new_AGEMA_signal_8956), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .Z0_f (new_AGEMA_signal_9194), .Z1_t (new_AGEMA_signal_9195), .Z1_f (new_AGEMA_signal_9196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .A0_f (new_AGEMA_signal_9188), .A1_t (new_AGEMA_signal_9189), .A1_f (new_AGEMA_signal_9190), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .B0_f (new_AGEMA_signal_9191), .B1_t (new_AGEMA_signal_9192), .B1_f (new_AGEMA_signal_9193), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28), .Z0_f (new_AGEMA_signal_9437), .Z1_t (new_AGEMA_signal_9438), .Z1_f (new_AGEMA_signal_9439) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28), .A0_f (new_AGEMA_signal_9437), .A1_t (new_AGEMA_signal_9438), .A1_f (new_AGEMA_signal_9439), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .B0_f (new_AGEMA_signal_9194), .B1_t (new_AGEMA_signal_9195), .B1_f (new_AGEMA_signal_9196), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29), .Z0_f (new_AGEMA_signal_9731), .Z1_t (new_AGEMA_signal_9732), .Z1_f (new_AGEMA_signal_9733) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M30_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26), .A0_f (new_AGEMA_signal_9434), .A1_t (new_AGEMA_signal_9435), .A1_f (new_AGEMA_signal_9436), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .B0_f (new_AGEMA_signal_9431), .B1_t (new_AGEMA_signal_9432), .B1_f (new_AGEMA_signal_9433), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30), .Z0_f (new_AGEMA_signal_9734), .Z1_t (new_AGEMA_signal_9735), .Z1_f (new_AGEMA_signal_9736) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M31_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .A0_f (new_AGEMA_signal_8951), .A1_t (new_AGEMA_signal_8952), .A1_f (new_AGEMA_signal_8953), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .B0_f (new_AGEMA_signal_9188), .B1_t (new_AGEMA_signal_9189), .B1_f (new_AGEMA_signal_9190), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31), .Z0_f (new_AGEMA_signal_9440), .Z1_t (new_AGEMA_signal_9441), .Z1_f (new_AGEMA_signal_9442) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M32_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .A0_f (new_AGEMA_signal_9194), .A1_t (new_AGEMA_signal_9195), .A1_f (new_AGEMA_signal_9196), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31), .B0_f (new_AGEMA_signal_9440), .B1_t (new_AGEMA_signal_9441), .B1_f (new_AGEMA_signal_9442), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32), .Z0_f (new_AGEMA_signal_9737), .Z1_t (new_AGEMA_signal_9738), .Z1_f (new_AGEMA_signal_9739) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M33_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .A0_f (new_AGEMA_signal_9194), .A1_t (new_AGEMA_signal_9195), .A1_f (new_AGEMA_signal_9196), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .B0_f (new_AGEMA_signal_9191), .B1_t (new_AGEMA_signal_9192), .B1_f (new_AGEMA_signal_9193), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33), .Z0_f (new_AGEMA_signal_9443), .Z1_t (new_AGEMA_signal_9444), .Z1_f (new_AGEMA_signal_9445) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M34_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .A0_f (new_AGEMA_signal_8954), .A1_t (new_AGEMA_signal_8955), .A1_f (new_AGEMA_signal_8956), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .B0_f (new_AGEMA_signal_8957), .B1_t (new_AGEMA_signal_8958), .B1_f (new_AGEMA_signal_8959), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34), .Z0_f (new_AGEMA_signal_9197), .Z1_t (new_AGEMA_signal_9198), .Z1_f (new_AGEMA_signal_9199) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M35_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .A0_f (new_AGEMA_signal_9431), .A1_t (new_AGEMA_signal_9432), .A1_f (new_AGEMA_signal_9433), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34), .B0_f (new_AGEMA_signal_9197), .B1_t (new_AGEMA_signal_9198), .B1_f (new_AGEMA_signal_9199), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35), .Z0_f (new_AGEMA_signal_9740), .Z1_t (new_AGEMA_signal_9741), .Z1_f (new_AGEMA_signal_9742) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M36_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .A0_f (new_AGEMA_signal_9431), .A1_t (new_AGEMA_signal_9432), .A1_f (new_AGEMA_signal_9433), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .B0_f (new_AGEMA_signal_9191), .B1_t (new_AGEMA_signal_9192), .B1_f (new_AGEMA_signal_9193), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36), .Z0_f (new_AGEMA_signal_9743), .Z1_t (new_AGEMA_signal_9744), .Z1_f (new_AGEMA_signal_9745) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M37_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .A0_f (new_AGEMA_signal_8954), .A1_t (new_AGEMA_signal_8955), .A1_f (new_AGEMA_signal_8956), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29), .B0_f (new_AGEMA_signal_9731), .B1_t (new_AGEMA_signal_9732), .B1_f (new_AGEMA_signal_9733), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .Z0_f (new_AGEMA_signal_10028), .Z1_t (new_AGEMA_signal_10029), .Z1_f (new_AGEMA_signal_10030) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M38_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32), .A0_f (new_AGEMA_signal_9737), .A1_t (new_AGEMA_signal_9738), .A1_f (new_AGEMA_signal_9739), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33), .B0_f (new_AGEMA_signal_9443), .B1_t (new_AGEMA_signal_9444), .B1_f (new_AGEMA_signal_9445), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .Z0_f (new_AGEMA_signal_10031), .Z1_t (new_AGEMA_signal_10032), .Z1_f (new_AGEMA_signal_10033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M39_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .A0_f (new_AGEMA_signal_9188), .A1_t (new_AGEMA_signal_9189), .A1_f (new_AGEMA_signal_9190), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30), .B0_f (new_AGEMA_signal_9734), .B1_t (new_AGEMA_signal_9735), .B1_f (new_AGEMA_signal_9736), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .Z0_f (new_AGEMA_signal_10034), .Z1_t (new_AGEMA_signal_10035), .Z1_f (new_AGEMA_signal_10036) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M40_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35), .A0_f (new_AGEMA_signal_9740), .A1_t (new_AGEMA_signal_9741), .A1_f (new_AGEMA_signal_9742), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36), .B0_f (new_AGEMA_signal_9743), .B1_t (new_AGEMA_signal_9744), .B1_f (new_AGEMA_signal_9745), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .Z0_f (new_AGEMA_signal_10037), .Z1_t (new_AGEMA_signal_10038), .Z1_f (new_AGEMA_signal_10039) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M41_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .A0_f (new_AGEMA_signal_10031), .A1_t (new_AGEMA_signal_10032), .A1_f (new_AGEMA_signal_10033), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .B0_f (new_AGEMA_signal_10037), .B1_t (new_AGEMA_signal_10038), .B1_f (new_AGEMA_signal_10039), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .Z0_f (new_AGEMA_signal_10292), .Z1_t (new_AGEMA_signal_10293), .Z1_f (new_AGEMA_signal_10294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M42_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .A0_f (new_AGEMA_signal_10028), .A1_t (new_AGEMA_signal_10029), .A1_f (new_AGEMA_signal_10030), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .B0_f (new_AGEMA_signal_10034), .B1_t (new_AGEMA_signal_10035), .B1_f (new_AGEMA_signal_10036), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .Z0_f (new_AGEMA_signal_10295), .Z1_t (new_AGEMA_signal_10296), .Z1_f (new_AGEMA_signal_10297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M43_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .A0_f (new_AGEMA_signal_10028), .A1_t (new_AGEMA_signal_10029), .A1_f (new_AGEMA_signal_10030), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .B0_f (new_AGEMA_signal_10031), .B1_t (new_AGEMA_signal_10032), .B1_f (new_AGEMA_signal_10033), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43), .Z0_f (new_AGEMA_signal_10298), .Z1_t (new_AGEMA_signal_10299), .Z1_f (new_AGEMA_signal_10300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M44_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .A0_f (new_AGEMA_signal_10034), .A1_t (new_AGEMA_signal_10035), .A1_f (new_AGEMA_signal_10036), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .B0_f (new_AGEMA_signal_10037), .B1_t (new_AGEMA_signal_10038), .B1_f (new_AGEMA_signal_10039), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44), .Z0_f (new_AGEMA_signal_10301), .Z1_t (new_AGEMA_signal_10302), .Z1_f (new_AGEMA_signal_10303) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M45_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .A0_f (new_AGEMA_signal_10295), .A1_t (new_AGEMA_signal_10296), .A1_f (new_AGEMA_signal_10297), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .B0_f (new_AGEMA_signal_10292), .B1_t (new_AGEMA_signal_10293), .B1_f (new_AGEMA_signal_10294), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45), .Z0_f (new_AGEMA_signal_11012), .Z1_t (new_AGEMA_signal_11013), .Z1_f (new_AGEMA_signal_11014) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M46_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44), .A0_f (new_AGEMA_signal_10301), .A1_t (new_AGEMA_signal_10302), .A1_f (new_AGEMA_signal_10303), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .B0_f (new_AGEMA_signal_6850), .B1_t (new_AGEMA_signal_6851), .B1_f (new_AGEMA_signal_6852), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46), .Z0_f (new_AGEMA_signal_11015), .Z1_t (new_AGEMA_signal_11016), .Z1_f (new_AGEMA_signal_11017) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M47_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .A0_f (new_AGEMA_signal_10037), .A1_t (new_AGEMA_signal_10038), .A1_f (new_AGEMA_signal_10039), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .B0_f (new_AGEMA_signal_7351), .B1_t (new_AGEMA_signal_7352), .B1_f (new_AGEMA_signal_7353), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47), .Z0_f (new_AGEMA_signal_10304), .Z1_t (new_AGEMA_signal_10305), .Z1_f (new_AGEMA_signal_10306) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M48_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .A0_f (new_AGEMA_signal_10034), .A1_t (new_AGEMA_signal_10035), .A1_f (new_AGEMA_signal_10036), .B0_t (RoundKey[8]), .B0_f (new_AGEMA_signal_6107), .B1_t (new_AGEMA_signal_6108), .B1_f (new_AGEMA_signal_6109), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48), .Z0_f (new_AGEMA_signal_10307), .Z1_t (new_AGEMA_signal_10308), .Z1_f (new_AGEMA_signal_10309) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M49_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43), .A0_f (new_AGEMA_signal_10298), .A1_t (new_AGEMA_signal_10299), .A1_f (new_AGEMA_signal_10300), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .B0_f (new_AGEMA_signal_6862), .B1_t (new_AGEMA_signal_6863), .B1_f (new_AGEMA_signal_6864), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49), .Z0_f (new_AGEMA_signal_11018), .Z1_t (new_AGEMA_signal_11019), .Z1_f (new_AGEMA_signal_11020) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M50_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .A0_f (new_AGEMA_signal_10031), .A1_t (new_AGEMA_signal_10032), .A1_f (new_AGEMA_signal_10033), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .B0_f (new_AGEMA_signal_6853), .B1_t (new_AGEMA_signal_6854), .B1_f (new_AGEMA_signal_6855), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50), .Z0_f (new_AGEMA_signal_10310), .Z1_t (new_AGEMA_signal_10311), .Z1_f (new_AGEMA_signal_10312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M51_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .A0_f (new_AGEMA_signal_10028), .A1_t (new_AGEMA_signal_10029), .A1_f (new_AGEMA_signal_10030), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .B0_f (new_AGEMA_signal_7360), .B1_t (new_AGEMA_signal_7361), .B1_f (new_AGEMA_signal_7362), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51), .Z0_f (new_AGEMA_signal_10313), .Z1_t (new_AGEMA_signal_10314), .Z1_f (new_AGEMA_signal_10315) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M52_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .A0_f (new_AGEMA_signal_10295), .A1_t (new_AGEMA_signal_10296), .A1_f (new_AGEMA_signal_10297), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .B0_f (new_AGEMA_signal_6859), .B1_t (new_AGEMA_signal_6860), .B1_f (new_AGEMA_signal_6861), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52), .Z0_f (new_AGEMA_signal_11021), .Z1_t (new_AGEMA_signal_11022), .Z1_f (new_AGEMA_signal_11023) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M53_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45), .A0_f (new_AGEMA_signal_11012), .A1_t (new_AGEMA_signal_11013), .A1_f (new_AGEMA_signal_11014), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .B0_f (new_AGEMA_signal_6871), .B1_t (new_AGEMA_signal_6872), .B1_f (new_AGEMA_signal_6873), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53), .Z0_f (new_AGEMA_signal_11726), .Z1_t (new_AGEMA_signal_11727), .Z1_f (new_AGEMA_signal_11728) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M54_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .A0_f (new_AGEMA_signal_10292), .A1_t (new_AGEMA_signal_10293), .A1_f (new_AGEMA_signal_10294), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .B0_f (new_AGEMA_signal_7354), .B1_t (new_AGEMA_signal_7355), .B1_f (new_AGEMA_signal_7356), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54), .Z0_f (new_AGEMA_signal_11024), .Z1_t (new_AGEMA_signal_11025), .Z1_f (new_AGEMA_signal_11026) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M55_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44), .A0_f (new_AGEMA_signal_10301), .A1_t (new_AGEMA_signal_10302), .A1_f (new_AGEMA_signal_10303), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .B0_f (new_AGEMA_signal_6856), .B1_t (new_AGEMA_signal_6857), .B1_f (new_AGEMA_signal_6858), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55), .Z0_f (new_AGEMA_signal_11027), .Z1_t (new_AGEMA_signal_11028), .Z1_f (new_AGEMA_signal_11029) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M56_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .A0_f (new_AGEMA_signal_10037), .A1_t (new_AGEMA_signal_10038), .A1_f (new_AGEMA_signal_10039), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .B0_f (new_AGEMA_signal_7366), .B1_t (new_AGEMA_signal_7367), .B1_f (new_AGEMA_signal_7368), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56), .Z0_f (new_AGEMA_signal_10316), .Z1_t (new_AGEMA_signal_10317), .Z1_f (new_AGEMA_signal_10318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M57_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .A0_f (new_AGEMA_signal_10034), .A1_t (new_AGEMA_signal_10035), .A1_f (new_AGEMA_signal_10036), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .B0_f (new_AGEMA_signal_6865), .B1_t (new_AGEMA_signal_6866), .B1_f (new_AGEMA_signal_6867), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57), .Z0_f (new_AGEMA_signal_10319), .Z1_t (new_AGEMA_signal_10320), .Z1_f (new_AGEMA_signal_10321) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M58_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43), .A0_f (new_AGEMA_signal_10298), .A1_t (new_AGEMA_signal_10299), .A1_f (new_AGEMA_signal_10300), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .B0_f (new_AGEMA_signal_6249), .B1_t (new_AGEMA_signal_6250), .B1_f (new_AGEMA_signal_6251), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58), .Z0_f (new_AGEMA_signal_11030), .Z1_t (new_AGEMA_signal_11031), .Z1_f (new_AGEMA_signal_11032) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M59_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .A0_f (new_AGEMA_signal_10031), .A1_t (new_AGEMA_signal_10032), .A1_f (new_AGEMA_signal_10033), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .B0_f (new_AGEMA_signal_6868), .B1_t (new_AGEMA_signal_6869), .B1_f (new_AGEMA_signal_6870), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59), .Z0_f (new_AGEMA_signal_10322), .Z1_t (new_AGEMA_signal_10323), .Z1_f (new_AGEMA_signal_10324) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M60_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .A0_f (new_AGEMA_signal_10028), .A1_t (new_AGEMA_signal_10029), .A1_f (new_AGEMA_signal_10030), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .B0_f (new_AGEMA_signal_7363), .B1_t (new_AGEMA_signal_7364), .B1_f (new_AGEMA_signal_7365), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60), .Z0_f (new_AGEMA_signal_10325), .Z1_t (new_AGEMA_signal_10326), .Z1_f (new_AGEMA_signal_10327) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M61_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .A0_f (new_AGEMA_signal_10295), .A1_t (new_AGEMA_signal_10296), .A1_f (new_AGEMA_signal_10297), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .B0_f (new_AGEMA_signal_6243), .B1_t (new_AGEMA_signal_6244), .B1_f (new_AGEMA_signal_6245), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .Z0_f (new_AGEMA_signal_11033), .Z1_t (new_AGEMA_signal_11034), .Z1_f (new_AGEMA_signal_11035) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M62_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45), .A0_f (new_AGEMA_signal_11012), .A1_t (new_AGEMA_signal_11013), .A1_f (new_AGEMA_signal_11014), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .B0_f (new_AGEMA_signal_6252), .B1_t (new_AGEMA_signal_6253), .B1_f (new_AGEMA_signal_6254), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62), .Z0_f (new_AGEMA_signal_11729), .Z1_t (new_AGEMA_signal_11730), .Z1_f (new_AGEMA_signal_11731) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M63_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .A0_f (new_AGEMA_signal_10292), .A1_t (new_AGEMA_signal_10293), .A1_f (new_AGEMA_signal_10294), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .B0_f (new_AGEMA_signal_6246), .B1_t (new_AGEMA_signal_6247), .B1_f (new_AGEMA_signal_6248), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63), .Z0_f (new_AGEMA_signal_11036), .Z1_t (new_AGEMA_signal_11037), .Z1_f (new_AGEMA_signal_11038) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .A0_f (new_AGEMA_signal_11033), .A1_t (new_AGEMA_signal_11034), .A1_f (new_AGEMA_signal_11035), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62), .B0_f (new_AGEMA_signal_11729), .B1_t (new_AGEMA_signal_11730), .B1_f (new_AGEMA_signal_11731), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .Z0_f (new_AGEMA_signal_12323), .Z1_t (new_AGEMA_signal_12324), .Z1_f (new_AGEMA_signal_12325) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50), .A0_f (new_AGEMA_signal_10310), .A1_t (new_AGEMA_signal_10311), .A1_f (new_AGEMA_signal_10312), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56), .B0_f (new_AGEMA_signal_10316), .B1_t (new_AGEMA_signal_10317), .B1_f (new_AGEMA_signal_10318), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .Z0_f (new_AGEMA_signal_11039), .Z1_t (new_AGEMA_signal_11040), .Z1_f (new_AGEMA_signal_11041) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46), .A0_f (new_AGEMA_signal_11015), .A1_t (new_AGEMA_signal_11016), .A1_f (new_AGEMA_signal_11017), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48), .B0_f (new_AGEMA_signal_10307), .B1_t (new_AGEMA_signal_10308), .B1_f (new_AGEMA_signal_10309), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2), .Z0_f (new_AGEMA_signal_11732), .Z1_t (new_AGEMA_signal_11733), .Z1_f (new_AGEMA_signal_11734) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47), .A0_f (new_AGEMA_signal_10304), .A1_t (new_AGEMA_signal_10305), .A1_f (new_AGEMA_signal_10306), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55), .B0_f (new_AGEMA_signal_11027), .B1_t (new_AGEMA_signal_11028), .B1_f (new_AGEMA_signal_11029), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3), .Z0_f (new_AGEMA_signal_11735), .Z1_t (new_AGEMA_signal_11736), .Z1_f (new_AGEMA_signal_11737) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54), .A0_f (new_AGEMA_signal_11024), .A1_t (new_AGEMA_signal_11025), .A1_f (new_AGEMA_signal_11026), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58), .B0_f (new_AGEMA_signal_11030), .B1_t (new_AGEMA_signal_11031), .B1_f (new_AGEMA_signal_11032), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4), .Z0_f (new_AGEMA_signal_11738), .Z1_t (new_AGEMA_signal_11739), .Z1_f (new_AGEMA_signal_11740) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49), .A0_f (new_AGEMA_signal_11018), .A1_t (new_AGEMA_signal_11019), .A1_f (new_AGEMA_signal_11020), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .B0_f (new_AGEMA_signal_11033), .B1_t (new_AGEMA_signal_11034), .B1_f (new_AGEMA_signal_11035), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5), .Z0_f (new_AGEMA_signal_11741), .Z1_t (new_AGEMA_signal_11742), .Z1_f (new_AGEMA_signal_11743) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62), .A0_f (new_AGEMA_signal_11729), .A1_t (new_AGEMA_signal_11730), .A1_f (new_AGEMA_signal_11731), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5), .B0_f (new_AGEMA_signal_11741), .B1_t (new_AGEMA_signal_11742), .B1_f (new_AGEMA_signal_11743), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .Z0_f (new_AGEMA_signal_12326), .Z1_t (new_AGEMA_signal_12327), .Z1_f (new_AGEMA_signal_12328) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46), .A0_f (new_AGEMA_signal_11015), .A1_t (new_AGEMA_signal_11016), .A1_f (new_AGEMA_signal_11017), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3), .B0_f (new_AGEMA_signal_11735), .B1_t (new_AGEMA_signal_11736), .B1_f (new_AGEMA_signal_11737), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7), .Z0_f (new_AGEMA_signal_12329), .Z1_t (new_AGEMA_signal_12330), .Z1_f (new_AGEMA_signal_12331) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51), .A0_f (new_AGEMA_signal_10313), .A1_t (new_AGEMA_signal_10314), .A1_f (new_AGEMA_signal_10315), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59), .B0_f (new_AGEMA_signal_10322), .B1_t (new_AGEMA_signal_10323), .B1_f (new_AGEMA_signal_10324), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8), .Z0_f (new_AGEMA_signal_11042), .Z1_t (new_AGEMA_signal_11043), .Z1_f (new_AGEMA_signal_11044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52), .A0_f (new_AGEMA_signal_11021), .A1_t (new_AGEMA_signal_11022), .A1_f (new_AGEMA_signal_11023), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53), .B0_f (new_AGEMA_signal_11726), .B1_t (new_AGEMA_signal_11727), .B1_f (new_AGEMA_signal_11728), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9), .Z0_f (new_AGEMA_signal_12332), .Z1_t (new_AGEMA_signal_12333), .Z1_f (new_AGEMA_signal_12334) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53), .A0_f (new_AGEMA_signal_11726), .A1_t (new_AGEMA_signal_11727), .A1_f (new_AGEMA_signal_11728), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4), .B0_f (new_AGEMA_signal_11738), .B1_t (new_AGEMA_signal_11739), .B1_f (new_AGEMA_signal_11740), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10), .Z0_f (new_AGEMA_signal_12335), .Z1_t (new_AGEMA_signal_12336), .Z1_f (new_AGEMA_signal_12337) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60), .A0_f (new_AGEMA_signal_10325), .A1_t (new_AGEMA_signal_10326), .A1_f (new_AGEMA_signal_10327), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2), .B0_f (new_AGEMA_signal_11732), .B1_t (new_AGEMA_signal_11733), .B1_f (new_AGEMA_signal_11734), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11), .Z0_f (new_AGEMA_signal_12338), .Z1_t (new_AGEMA_signal_12339), .Z1_f (new_AGEMA_signal_12340) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48), .A0_f (new_AGEMA_signal_10307), .A1_t (new_AGEMA_signal_10308), .A1_f (new_AGEMA_signal_10309), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51), .B0_f (new_AGEMA_signal_10313), .B1_t (new_AGEMA_signal_10314), .B1_f (new_AGEMA_signal_10315), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12), .Z0_f (new_AGEMA_signal_11045), .Z1_t (new_AGEMA_signal_11046), .Z1_f (new_AGEMA_signal_11047) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50), .A0_f (new_AGEMA_signal_10310), .A1_t (new_AGEMA_signal_10311), .A1_f (new_AGEMA_signal_10312), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .B0_f (new_AGEMA_signal_12323), .B1_t (new_AGEMA_signal_12324), .B1_f (new_AGEMA_signal_12325), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13), .Z0_f (new_AGEMA_signal_12869), .Z1_t (new_AGEMA_signal_12870), .Z1_f (new_AGEMA_signal_12871) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52), .A0_f (new_AGEMA_signal_11021), .A1_t (new_AGEMA_signal_11022), .A1_f (new_AGEMA_signal_11023), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .B0_f (new_AGEMA_signal_11033), .B1_t (new_AGEMA_signal_11034), .B1_f (new_AGEMA_signal_11035), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14), .Z0_f (new_AGEMA_signal_11744), .Z1_t (new_AGEMA_signal_11745), .Z1_f (new_AGEMA_signal_11746) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55), .A0_f (new_AGEMA_signal_11027), .A1_t (new_AGEMA_signal_11028), .A1_f (new_AGEMA_signal_11029), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .B0_f (new_AGEMA_signal_11039), .B1_t (new_AGEMA_signal_11040), .B1_f (new_AGEMA_signal_11041), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15), .Z0_f (new_AGEMA_signal_11747), .Z1_t (new_AGEMA_signal_11748), .Z1_f (new_AGEMA_signal_11749) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56), .A0_f (new_AGEMA_signal_10316), .A1_t (new_AGEMA_signal_10317), .A1_f (new_AGEMA_signal_10318), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .B0_f (new_AGEMA_signal_12323), .B1_t (new_AGEMA_signal_12324), .B1_f (new_AGEMA_signal_12325), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16), .Z0_f (new_AGEMA_signal_12872), .Z1_t (new_AGEMA_signal_12873), .Z1_f (new_AGEMA_signal_12874) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57), .A0_f (new_AGEMA_signal_10319), .A1_t (new_AGEMA_signal_10320), .A1_f (new_AGEMA_signal_10321), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .B0_f (new_AGEMA_signal_11039), .B1_t (new_AGEMA_signal_11040), .B1_f (new_AGEMA_signal_11041), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17), .Z0_f (new_AGEMA_signal_11750), .Z1_t (new_AGEMA_signal_11751), .Z1_f (new_AGEMA_signal_11752) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58), .A0_f (new_AGEMA_signal_11030), .A1_t (new_AGEMA_signal_11031), .A1_f (new_AGEMA_signal_11032), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8), .B0_f (new_AGEMA_signal_11042), .B1_t (new_AGEMA_signal_11043), .B1_f (new_AGEMA_signal_11044), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18), .Z0_f (new_AGEMA_signal_11753), .Z1_t (new_AGEMA_signal_11754), .Z1_f (new_AGEMA_signal_11755) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63), .A0_f (new_AGEMA_signal_11036), .A1_t (new_AGEMA_signal_11037), .A1_f (new_AGEMA_signal_11038), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4), .B0_f (new_AGEMA_signal_11738), .B1_t (new_AGEMA_signal_11739), .B1_f (new_AGEMA_signal_11740), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19), .Z0_f (new_AGEMA_signal_12341), .Z1_t (new_AGEMA_signal_12342), .Z1_f (new_AGEMA_signal_12343) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .A0_f (new_AGEMA_signal_12323), .A1_t (new_AGEMA_signal_12324), .A1_f (new_AGEMA_signal_12325), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .B0_f (new_AGEMA_signal_11039), .B1_t (new_AGEMA_signal_11040), .B1_f (new_AGEMA_signal_11041), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20), .Z0_f (new_AGEMA_signal_12875), .Z1_t (new_AGEMA_signal_12876), .Z1_f (new_AGEMA_signal_12877) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .A0_f (new_AGEMA_signal_11039), .A1_t (new_AGEMA_signal_11040), .A1_f (new_AGEMA_signal_11041), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7), .B0_f (new_AGEMA_signal_12329), .B1_t (new_AGEMA_signal_12330), .B1_f (new_AGEMA_signal_12331), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21), .Z0_f (new_AGEMA_signal_12878), .Z1_t (new_AGEMA_signal_12879), .Z1_f (new_AGEMA_signal_12880) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3), .A0_f (new_AGEMA_signal_11735), .A1_t (new_AGEMA_signal_11736), .A1_f (new_AGEMA_signal_11737), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12), .B0_f (new_AGEMA_signal_11045), .B1_t (new_AGEMA_signal_11046), .B1_f (new_AGEMA_signal_11047), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22), .Z0_f (new_AGEMA_signal_12344), .Z1_t (new_AGEMA_signal_12345), .Z1_f (new_AGEMA_signal_12346) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18), .A0_f (new_AGEMA_signal_11753), .A1_t (new_AGEMA_signal_11754), .A1_f (new_AGEMA_signal_11755), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2), .B0_f (new_AGEMA_signal_11732), .B1_t (new_AGEMA_signal_11733), .B1_f (new_AGEMA_signal_11734), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23), .Z0_f (new_AGEMA_signal_12347), .Z1_t (new_AGEMA_signal_12348), .Z1_f (new_AGEMA_signal_12349) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15), .A0_f (new_AGEMA_signal_11747), .A1_t (new_AGEMA_signal_11748), .A1_f (new_AGEMA_signal_11749), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9), .B0_f (new_AGEMA_signal_12332), .B1_t (new_AGEMA_signal_12333), .B1_f (new_AGEMA_signal_12334), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24), .Z0_f (new_AGEMA_signal_12881), .Z1_t (new_AGEMA_signal_12882), .Z1_f (new_AGEMA_signal_12883) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .A0_f (new_AGEMA_signal_12326), .A1_t (new_AGEMA_signal_12327), .A1_f (new_AGEMA_signal_12328), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10), .B0_f (new_AGEMA_signal_12335), .B1_t (new_AGEMA_signal_12336), .B1_f (new_AGEMA_signal_12337), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25), .Z0_f (new_AGEMA_signal_12884), .Z1_t (new_AGEMA_signal_12885), .Z1_f (new_AGEMA_signal_12886) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7), .A0_f (new_AGEMA_signal_12329), .A1_t (new_AGEMA_signal_12330), .A1_f (new_AGEMA_signal_12331), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9), .B0_f (new_AGEMA_signal_12332), .B1_t (new_AGEMA_signal_12333), .B1_f (new_AGEMA_signal_12334), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26), .Z0_f (new_AGEMA_signal_12887), .Z1_t (new_AGEMA_signal_12888), .Z1_f (new_AGEMA_signal_12889) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8), .A0_f (new_AGEMA_signal_11042), .A1_t (new_AGEMA_signal_11043), .A1_f (new_AGEMA_signal_11044), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10), .B0_f (new_AGEMA_signal_12335), .B1_t (new_AGEMA_signal_12336), .B1_f (new_AGEMA_signal_12337), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27), .Z0_f (new_AGEMA_signal_12890), .Z1_t (new_AGEMA_signal_12891), .Z1_f (new_AGEMA_signal_12892) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11), .A0_f (new_AGEMA_signal_12338), .A1_t (new_AGEMA_signal_12339), .A1_f (new_AGEMA_signal_12340), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14), .B0_f (new_AGEMA_signal_11744), .B1_t (new_AGEMA_signal_11745), .B1_f (new_AGEMA_signal_11746), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28), .Z0_f (new_AGEMA_signal_12893), .Z1_t (new_AGEMA_signal_12894), .Z1_f (new_AGEMA_signal_12895) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11), .A0_f (new_AGEMA_signal_12338), .A1_t (new_AGEMA_signal_12339), .A1_f (new_AGEMA_signal_12340), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17), .B0_f (new_AGEMA_signal_11750), .B1_t (new_AGEMA_signal_11751), .B1_f (new_AGEMA_signal_11752), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29), .Z0_f (new_AGEMA_signal_12896), .Z1_t (new_AGEMA_signal_12897), .Z1_f (new_AGEMA_signal_12898) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .A0_f (new_AGEMA_signal_12326), .A1_t (new_AGEMA_signal_12327), .A1_f (new_AGEMA_signal_12328), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24), .B0_f (new_AGEMA_signal_12881), .B1_t (new_AGEMA_signal_12882), .B1_f (new_AGEMA_signal_12883), .Z0_t (KeyExpansionIns_tmp[23]), .Z0_f (new_AGEMA_signal_13529), .Z1_t (new_AGEMA_signal_13530), .Z1_f (new_AGEMA_signal_13531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16), .A0_f (new_AGEMA_signal_12872), .A1_t (new_AGEMA_signal_12873), .A1_f (new_AGEMA_signal_12874), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26), .B0_f (new_AGEMA_signal_12887), .B1_t (new_AGEMA_signal_12888), .B1_f (new_AGEMA_signal_12889), .Z0_t (KeyExpansionIns_tmp[22]), .Z0_f (new_AGEMA_signal_13532), .Z1_t (new_AGEMA_signal_13533), .Z1_f (new_AGEMA_signal_13534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19), .A0_f (new_AGEMA_signal_12341), .A1_t (new_AGEMA_signal_12342), .A1_f (new_AGEMA_signal_12343), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28), .B0_f (new_AGEMA_signal_12893), .B1_t (new_AGEMA_signal_12894), .B1_f (new_AGEMA_signal_12895), .Z0_t (KeyExpansionIns_tmp[21]), .Z0_f (new_AGEMA_signal_13535), .Z1_t (new_AGEMA_signal_13536), .Z1_f (new_AGEMA_signal_13537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .A0_f (new_AGEMA_signal_12326), .A1_t (new_AGEMA_signal_12327), .A1_f (new_AGEMA_signal_12328), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21), .B0_f (new_AGEMA_signal_12878), .B1_t (new_AGEMA_signal_12879), .B1_f (new_AGEMA_signal_12880), .Z0_t (KeyExpansionIns_tmp[20]), .Z0_f (new_AGEMA_signal_13538), .Z1_t (new_AGEMA_signal_13539), .Z1_f (new_AGEMA_signal_13540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20), .A0_f (new_AGEMA_signal_12875), .A1_t (new_AGEMA_signal_12876), .A1_f (new_AGEMA_signal_12877), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22), .B0_f (new_AGEMA_signal_12344), .B1_t (new_AGEMA_signal_12345), .B1_f (new_AGEMA_signal_12346), .Z0_t (KeyExpansionIns_tmp[19]), .Z0_f (new_AGEMA_signal_13541), .Z1_t (new_AGEMA_signal_13542), .Z1_f (new_AGEMA_signal_13543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25), .A0_f (new_AGEMA_signal_12884), .A1_t (new_AGEMA_signal_12885), .A1_f (new_AGEMA_signal_12886), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29), .B0_f (new_AGEMA_signal_12896), .B1_t (new_AGEMA_signal_12897), .B1_f (new_AGEMA_signal_12898), .Z0_t (KeyExpansionIns_tmp[18]), .Z0_f (new_AGEMA_signal_13544), .Z1_t (new_AGEMA_signal_13545), .Z1_f (new_AGEMA_signal_13546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13), .A0_f (new_AGEMA_signal_12869), .A1_t (new_AGEMA_signal_12870), .A1_f (new_AGEMA_signal_12871), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27), .B0_f (new_AGEMA_signal_12890), .B1_t (new_AGEMA_signal_12891), .B1_f (new_AGEMA_signal_12892), .Z0_t (KeyExpansionIns_tmp[17]), .Z0_f (new_AGEMA_signal_13547), .Z1_t (new_AGEMA_signal_13548), .Z1_f (new_AGEMA_signal_13549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .A0_f (new_AGEMA_signal_12326), .A1_t (new_AGEMA_signal_12327), .A1_f (new_AGEMA_signal_12328), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23), .B0_f (new_AGEMA_signal_12347), .B1_t (new_AGEMA_signal_12348), .B1_f (new_AGEMA_signal_12349), .Z0_t (KeyExpansionIns_tmp[16]), .Z0_f (new_AGEMA_signal_12899), .Z1_t (new_AGEMA_signal_12900), .Z1_f (new_AGEMA_signal_12901) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T1_U1 ( .A0_t (RoundKey[7]), .A0_f (new_AGEMA_signal_6008), .A1_t (new_AGEMA_signal_6009), .A1_f (new_AGEMA_signal_6010), .B0_t (RoundKey[4]), .B0_f (new_AGEMA_signal_5711), .B1_t (new_AGEMA_signal_5712), .B1_f (new_AGEMA_signal_5713), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .Z0_f (new_AGEMA_signal_6273), .Z1_t (new_AGEMA_signal_6274), .Z1_f (new_AGEMA_signal_6275) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T2_U1 ( .A0_t (RoundKey[7]), .A0_f (new_AGEMA_signal_6008), .A1_t (new_AGEMA_signal_6009), .A1_f (new_AGEMA_signal_6010), .B0_t (RoundKey[2]), .B0_f (new_AGEMA_signal_5513), .B1_t (new_AGEMA_signal_5514), .B1_f (new_AGEMA_signal_5515), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .Z0_f (new_AGEMA_signal_6276), .Z1_t (new_AGEMA_signal_6277), .Z1_f (new_AGEMA_signal_6278) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T3_U1 ( .A0_t (RoundKey[7]), .A0_f (new_AGEMA_signal_6008), .A1_t (new_AGEMA_signal_6009), .A1_f (new_AGEMA_signal_6010), .B0_t (RoundKey[1]), .B0_f (new_AGEMA_signal_5414), .B1_t (new_AGEMA_signal_5415), .B1_f (new_AGEMA_signal_5416), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .Z0_f (new_AGEMA_signal_6279), .Z1_t (new_AGEMA_signal_6280), .Z1_f (new_AGEMA_signal_6281) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T4_U1 ( .A0_t (RoundKey[4]), .A0_f (new_AGEMA_signal_5711), .A1_t (new_AGEMA_signal_5712), .A1_f (new_AGEMA_signal_5713), .B0_t (RoundKey[2]), .B0_f (new_AGEMA_signal_5513), .B1_t (new_AGEMA_signal_5514), .B1_f (new_AGEMA_signal_5515), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .Z0_f (new_AGEMA_signal_6282), .Z1_t (new_AGEMA_signal_6283), .Z1_f (new_AGEMA_signal_6284) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T5_U1 ( .A0_t (RoundKey[3]), .A0_f (new_AGEMA_signal_5612), .A1_t (new_AGEMA_signal_5613), .A1_f (new_AGEMA_signal_5614), .B0_t (RoundKey[1]), .B0_f (new_AGEMA_signal_5414), .B1_t (new_AGEMA_signal_5415), .B1_f (new_AGEMA_signal_5416), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .Z0_f (new_AGEMA_signal_6285), .Z1_t (new_AGEMA_signal_6286), .Z1_f (new_AGEMA_signal_6287) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .A0_f (new_AGEMA_signal_6273), .A1_t (new_AGEMA_signal_6274), .A1_f (new_AGEMA_signal_6275), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .B0_f (new_AGEMA_signal_6285), .B1_t (new_AGEMA_signal_6286), .B1_f (new_AGEMA_signal_6287), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .Z0_f (new_AGEMA_signal_6874), .Z1_t (new_AGEMA_signal_6875), .Z1_f (new_AGEMA_signal_6876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T7_U1 ( .A0_t (RoundKey[6]), .A0_f (new_AGEMA_signal_5909), .A1_t (new_AGEMA_signal_5910), .A1_f (new_AGEMA_signal_5911), .B0_t (RoundKey[5]), .B0_f (new_AGEMA_signal_5810), .B1_t (new_AGEMA_signal_5811), .B1_f (new_AGEMA_signal_5812), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .Z0_f (new_AGEMA_signal_6288), .Z1_t (new_AGEMA_signal_6289), .Z1_f (new_AGEMA_signal_6290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T8_U1 ( .A0_t (RoundKey[0]), .A0_f (new_AGEMA_signal_5063), .A1_t (new_AGEMA_signal_5064), .A1_f (new_AGEMA_signal_5065), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .B0_f (new_AGEMA_signal_6874), .B1_t (new_AGEMA_signal_6875), .B1_f (new_AGEMA_signal_6876), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .Z0_f (new_AGEMA_signal_7390), .Z1_t (new_AGEMA_signal_7391), .Z1_f (new_AGEMA_signal_7392) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T9_U1 ( .A0_t (RoundKey[0]), .A0_f (new_AGEMA_signal_5063), .A1_t (new_AGEMA_signal_5064), .A1_f (new_AGEMA_signal_5065), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .B0_f (new_AGEMA_signal_6288), .B1_t (new_AGEMA_signal_6289), .B1_f (new_AGEMA_signal_6290), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .Z0_f (new_AGEMA_signal_6877), .Z1_t (new_AGEMA_signal_6878), .Z1_f (new_AGEMA_signal_6879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .A0_f (new_AGEMA_signal_6874), .A1_t (new_AGEMA_signal_6875), .A1_f (new_AGEMA_signal_6876), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .B0_f (new_AGEMA_signal_6288), .B1_t (new_AGEMA_signal_6289), .B1_f (new_AGEMA_signal_6290), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .Z0_f (new_AGEMA_signal_7393), .Z1_t (new_AGEMA_signal_7394), .Z1_f (new_AGEMA_signal_7395) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T11_U1 ( .A0_t (RoundKey[6]), .A0_f (new_AGEMA_signal_5909), .A1_t (new_AGEMA_signal_5910), .A1_f (new_AGEMA_signal_5911), .B0_t (RoundKey[2]), .B0_f (new_AGEMA_signal_5513), .B1_t (new_AGEMA_signal_5514), .B1_f (new_AGEMA_signal_5515), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11), .Z0_f (new_AGEMA_signal_6291), .Z1_t (new_AGEMA_signal_6292), .Z1_f (new_AGEMA_signal_6293) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T12_U1 ( .A0_t (RoundKey[5]), .A0_f (new_AGEMA_signal_5810), .A1_t (new_AGEMA_signal_5811), .A1_f (new_AGEMA_signal_5812), .B0_t (RoundKey[2]), .B0_f (new_AGEMA_signal_5513), .B1_t (new_AGEMA_signal_5514), .B1_f (new_AGEMA_signal_5515), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12), .Z0_f (new_AGEMA_signal_6294), .Z1_t (new_AGEMA_signal_6295), .Z1_f (new_AGEMA_signal_6296) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .A0_f (new_AGEMA_signal_6279), .A1_t (new_AGEMA_signal_6280), .A1_f (new_AGEMA_signal_6281), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .B0_f (new_AGEMA_signal_6282), .B1_t (new_AGEMA_signal_6283), .B1_f (new_AGEMA_signal_6284), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .Z0_f (new_AGEMA_signal_6880), .Z1_t (new_AGEMA_signal_6881), .Z1_f (new_AGEMA_signal_6882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .A0_f (new_AGEMA_signal_6874), .A1_t (new_AGEMA_signal_6875), .A1_f (new_AGEMA_signal_6876), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11), .B0_f (new_AGEMA_signal_6291), .B1_t (new_AGEMA_signal_6292), .B1_f (new_AGEMA_signal_6293), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14), .Z0_f (new_AGEMA_signal_7396), .Z1_t (new_AGEMA_signal_7397), .Z1_f (new_AGEMA_signal_7398) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .A0_f (new_AGEMA_signal_6285), .A1_t (new_AGEMA_signal_6286), .A1_f (new_AGEMA_signal_6287), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11), .B0_f (new_AGEMA_signal_6291), .B1_t (new_AGEMA_signal_6292), .B1_f (new_AGEMA_signal_6293), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .Z0_f (new_AGEMA_signal_6883), .Z1_t (new_AGEMA_signal_6884), .Z1_f (new_AGEMA_signal_6885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .A0_f (new_AGEMA_signal_6285), .A1_t (new_AGEMA_signal_6286), .A1_f (new_AGEMA_signal_6287), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12), .B0_f (new_AGEMA_signal_6294), .B1_t (new_AGEMA_signal_6295), .B1_f (new_AGEMA_signal_6296), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Z0_f (new_AGEMA_signal_6886), .Z1_t (new_AGEMA_signal_6887), .Z1_f (new_AGEMA_signal_6888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .A0_f (new_AGEMA_signal_6877), .A1_t (new_AGEMA_signal_6878), .A1_f (new_AGEMA_signal_6879), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .B0_f (new_AGEMA_signal_6886), .B1_t (new_AGEMA_signal_6887), .B1_f (new_AGEMA_signal_6888), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .Z0_f (new_AGEMA_signal_7399), .Z1_t (new_AGEMA_signal_7400), .Z1_f (new_AGEMA_signal_7401) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T18_U1 ( .A0_t (RoundKey[4]), .A0_f (new_AGEMA_signal_5711), .A1_t (new_AGEMA_signal_5712), .A1_f (new_AGEMA_signal_5713), .B0_t (RoundKey[0]), .B0_f (new_AGEMA_signal_5063), .B1_t (new_AGEMA_signal_5064), .B1_f (new_AGEMA_signal_5065), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18), .Z0_f (new_AGEMA_signal_6297), .Z1_t (new_AGEMA_signal_6298), .Z1_f (new_AGEMA_signal_6299) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .A0_f (new_AGEMA_signal_6288), .A1_t (new_AGEMA_signal_6289), .A1_f (new_AGEMA_signal_6290), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18), .B0_f (new_AGEMA_signal_6297), .B1_t (new_AGEMA_signal_6298), .B1_f (new_AGEMA_signal_6299), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .Z0_f (new_AGEMA_signal_6889), .Z1_t (new_AGEMA_signal_6890), .Z1_f (new_AGEMA_signal_6891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .A0_f (new_AGEMA_signal_6273), .A1_t (new_AGEMA_signal_6274), .A1_f (new_AGEMA_signal_6275), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .B0_f (new_AGEMA_signal_6889), .B1_t (new_AGEMA_signal_6890), .B1_f (new_AGEMA_signal_6891), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .Z0_f (new_AGEMA_signal_7402), .Z1_t (new_AGEMA_signal_7403), .Z1_f (new_AGEMA_signal_7404) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T21_U1 ( .A0_t (RoundKey[1]), .A0_f (new_AGEMA_signal_5414), .A1_t (new_AGEMA_signal_5415), .A1_f (new_AGEMA_signal_5416), .B0_t (RoundKey[0]), .B0_f (new_AGEMA_signal_5063), .B1_t (new_AGEMA_signal_5064), .B1_f (new_AGEMA_signal_5065), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21), .Z0_f (new_AGEMA_signal_6300), .Z1_t (new_AGEMA_signal_6301), .Z1_f (new_AGEMA_signal_6302) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .A0_f (new_AGEMA_signal_6288), .A1_t (new_AGEMA_signal_6289), .A1_f (new_AGEMA_signal_6290), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21), .B0_f (new_AGEMA_signal_6300), .B1_t (new_AGEMA_signal_6301), .B1_f (new_AGEMA_signal_6302), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .Z0_f (new_AGEMA_signal_6892), .Z1_t (new_AGEMA_signal_6893), .Z1_f (new_AGEMA_signal_6894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .A0_f (new_AGEMA_signal_6276), .A1_t (new_AGEMA_signal_6277), .A1_f (new_AGEMA_signal_6278), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .B0_f (new_AGEMA_signal_6892), .B1_t (new_AGEMA_signal_6893), .B1_f (new_AGEMA_signal_6894), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .Z0_f (new_AGEMA_signal_7405), .Z1_t (new_AGEMA_signal_7406), .Z1_f (new_AGEMA_signal_7407) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .A0_f (new_AGEMA_signal_6276), .A1_t (new_AGEMA_signal_6277), .A1_f (new_AGEMA_signal_6278), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .B0_f (new_AGEMA_signal_7393), .B1_t (new_AGEMA_signal_7394), .B1_f (new_AGEMA_signal_7395), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24), .Z0_f (new_AGEMA_signal_8150), .Z1_t (new_AGEMA_signal_8151), .Z1_f (new_AGEMA_signal_8152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .A0_f (new_AGEMA_signal_7402), .A1_t (new_AGEMA_signal_7403), .A1_f (new_AGEMA_signal_7404), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .B0_f (new_AGEMA_signal_7399), .B1_t (new_AGEMA_signal_7400), .B1_f (new_AGEMA_signal_7401), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25), .Z0_f (new_AGEMA_signal_8153), .Z1_t (new_AGEMA_signal_8154), .Z1_f (new_AGEMA_signal_8155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .A0_f (new_AGEMA_signal_6279), .A1_t (new_AGEMA_signal_6280), .A1_f (new_AGEMA_signal_6281), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .B0_f (new_AGEMA_signal_6886), .B1_t (new_AGEMA_signal_6887), .B1_f (new_AGEMA_signal_6888), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26), .Z0_f (new_AGEMA_signal_7408), .Z1_t (new_AGEMA_signal_7409), .Z1_f (new_AGEMA_signal_7410) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .A0_f (new_AGEMA_signal_6273), .A1_t (new_AGEMA_signal_6274), .A1_f (new_AGEMA_signal_6275), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12), .B0_f (new_AGEMA_signal_6294), .B1_t (new_AGEMA_signal_6295), .B1_f (new_AGEMA_signal_6296), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .Z0_f (new_AGEMA_signal_6895), .Z1_t (new_AGEMA_signal_6896), .Z1_f (new_AGEMA_signal_6897) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .A0_f (new_AGEMA_signal_6880), .A1_t (new_AGEMA_signal_6881), .A1_f (new_AGEMA_signal_6882), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .B0_f (new_AGEMA_signal_6874), .B1_t (new_AGEMA_signal_6875), .B1_f (new_AGEMA_signal_6876), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1), .Z0_f (new_AGEMA_signal_7411), .Z1_t (new_AGEMA_signal_7412), .Z1_f (new_AGEMA_signal_7413) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .A0_f (new_AGEMA_signal_7405), .A1_t (new_AGEMA_signal_7406), .A1_f (new_AGEMA_signal_7407), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .B0_f (new_AGEMA_signal_7390), .B1_t (new_AGEMA_signal_7391), .B1_f (new_AGEMA_signal_7392), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2), .Z0_f (new_AGEMA_signal_8156), .Z1_t (new_AGEMA_signal_8157), .Z1_f (new_AGEMA_signal_8158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14), .A0_f (new_AGEMA_signal_7396), .A1_t (new_AGEMA_signal_7397), .A1_f (new_AGEMA_signal_7398), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1), .B0_f (new_AGEMA_signal_7411), .B1_t (new_AGEMA_signal_7412), .B1_f (new_AGEMA_signal_7413), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3), .Z0_f (new_AGEMA_signal_8159), .Z1_t (new_AGEMA_signal_8160), .Z1_f (new_AGEMA_signal_8161) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .A0_f (new_AGEMA_signal_6889), .A1_t (new_AGEMA_signal_6890), .A1_f (new_AGEMA_signal_6891), .B0_t (RoundKey[0]), .B0_f (new_AGEMA_signal_5063), .B1_t (new_AGEMA_signal_5064), .B1_f (new_AGEMA_signal_5065), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4), .Z0_f (new_AGEMA_signal_7414), .Z1_t (new_AGEMA_signal_7415), .Z1_f (new_AGEMA_signal_7416) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4), .A0_f (new_AGEMA_signal_7414), .A1_t (new_AGEMA_signal_7415), .A1_f (new_AGEMA_signal_7416), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1), .B0_f (new_AGEMA_signal_7411), .B1_t (new_AGEMA_signal_7412), .B1_f (new_AGEMA_signal_7413), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5), .Z0_f (new_AGEMA_signal_8162), .Z1_t (new_AGEMA_signal_8163), .Z1_f (new_AGEMA_signal_8164) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .A0_f (new_AGEMA_signal_6279), .A1_t (new_AGEMA_signal_6280), .A1_f (new_AGEMA_signal_6281), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .B0_f (new_AGEMA_signal_6886), .B1_t (new_AGEMA_signal_6887), .B1_f (new_AGEMA_signal_6888), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6), .Z0_f (new_AGEMA_signal_7417), .Z1_t (new_AGEMA_signal_7418), .Z1_f (new_AGEMA_signal_7419) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .A0_f (new_AGEMA_signal_6892), .A1_t (new_AGEMA_signal_6893), .A1_f (new_AGEMA_signal_6894), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .B0_f (new_AGEMA_signal_6877), .B1_t (new_AGEMA_signal_6878), .B1_f (new_AGEMA_signal_6879), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7), .Z0_f (new_AGEMA_signal_7420), .Z1_t (new_AGEMA_signal_7421), .Z1_f (new_AGEMA_signal_7422) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26), .A0_f (new_AGEMA_signal_7408), .A1_t (new_AGEMA_signal_7409), .A1_f (new_AGEMA_signal_7410), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6), .B0_f (new_AGEMA_signal_7417), .B1_t (new_AGEMA_signal_7418), .B1_f (new_AGEMA_signal_7419), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8), .Z0_f (new_AGEMA_signal_8165), .Z1_t (new_AGEMA_signal_8166), .Z1_f (new_AGEMA_signal_8167) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .A0_f (new_AGEMA_signal_7402), .A1_t (new_AGEMA_signal_7403), .A1_f (new_AGEMA_signal_7404), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .B0_f (new_AGEMA_signal_7399), .B1_t (new_AGEMA_signal_7400), .B1_f (new_AGEMA_signal_7401), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9), .Z0_f (new_AGEMA_signal_8168), .Z1_t (new_AGEMA_signal_8169), .Z1_f (new_AGEMA_signal_8170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9), .A0_f (new_AGEMA_signal_8168), .A1_t (new_AGEMA_signal_8169), .A1_f (new_AGEMA_signal_8170), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6), .B0_f (new_AGEMA_signal_7417), .B1_t (new_AGEMA_signal_7418), .B1_f (new_AGEMA_signal_7419), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10), .Z0_f (new_AGEMA_signal_8666), .Z1_t (new_AGEMA_signal_8667), .Z1_f (new_AGEMA_signal_8668) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .A0_f (new_AGEMA_signal_6273), .A1_t (new_AGEMA_signal_6274), .A1_f (new_AGEMA_signal_6275), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .B0_f (new_AGEMA_signal_6883), .B1_t (new_AGEMA_signal_6884), .B1_f (new_AGEMA_signal_6885), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11), .Z0_f (new_AGEMA_signal_7423), .Z1_t (new_AGEMA_signal_7424), .Z1_f (new_AGEMA_signal_7425) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .A0_f (new_AGEMA_signal_6282), .A1_t (new_AGEMA_signal_6283), .A1_f (new_AGEMA_signal_6284), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .B0_f (new_AGEMA_signal_6895), .B1_t (new_AGEMA_signal_6896), .B1_f (new_AGEMA_signal_6897), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12), .Z0_f (new_AGEMA_signal_7426), .Z1_t (new_AGEMA_signal_7427), .Z1_f (new_AGEMA_signal_7428) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12), .A0_f (new_AGEMA_signal_7426), .A1_t (new_AGEMA_signal_7427), .A1_f (new_AGEMA_signal_7428), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11), .B0_f (new_AGEMA_signal_7423), .B1_t (new_AGEMA_signal_7424), .B1_f (new_AGEMA_signal_7425), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13), .Z0_f (new_AGEMA_signal_8171), .Z1_t (new_AGEMA_signal_8172), .Z1_f (new_AGEMA_signal_8173) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .A0_f (new_AGEMA_signal_6276), .A1_t (new_AGEMA_signal_6277), .A1_f (new_AGEMA_signal_6278), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .B0_f (new_AGEMA_signal_7393), .B1_t (new_AGEMA_signal_7394), .B1_f (new_AGEMA_signal_7395), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14), .Z0_f (new_AGEMA_signal_8174), .Z1_t (new_AGEMA_signal_8175), .Z1_f (new_AGEMA_signal_8176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14), .A0_f (new_AGEMA_signal_8174), .A1_t (new_AGEMA_signal_8175), .A1_f (new_AGEMA_signal_8176), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11), .B0_f (new_AGEMA_signal_7423), .B1_t (new_AGEMA_signal_7424), .B1_f (new_AGEMA_signal_7425), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15), .Z0_f (new_AGEMA_signal_8669), .Z1_t (new_AGEMA_signal_8670), .Z1_f (new_AGEMA_signal_8671) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3), .A0_f (new_AGEMA_signal_8159), .A1_t (new_AGEMA_signal_8160), .A1_f (new_AGEMA_signal_8161), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2), .B0_f (new_AGEMA_signal_8156), .B1_t (new_AGEMA_signal_8157), .B1_f (new_AGEMA_signal_8158), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16), .Z0_f (new_AGEMA_signal_8672), .Z1_t (new_AGEMA_signal_8673), .Z1_f (new_AGEMA_signal_8674) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5), .A0_f (new_AGEMA_signal_8162), .A1_t (new_AGEMA_signal_8163), .A1_f (new_AGEMA_signal_8164), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24), .B0_f (new_AGEMA_signal_8150), .B1_t (new_AGEMA_signal_8151), .B1_f (new_AGEMA_signal_8152), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17), .Z0_f (new_AGEMA_signal_8675), .Z1_t (new_AGEMA_signal_8676), .Z1_f (new_AGEMA_signal_8677) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8), .A0_f (new_AGEMA_signal_8165), .A1_t (new_AGEMA_signal_8166), .A1_f (new_AGEMA_signal_8167), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7), .B0_f (new_AGEMA_signal_7420), .B1_t (new_AGEMA_signal_7421), .B1_f (new_AGEMA_signal_7422), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18), .Z0_f (new_AGEMA_signal_8678), .Z1_t (new_AGEMA_signal_8679), .Z1_f (new_AGEMA_signal_8680) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10), .A0_f (new_AGEMA_signal_8666), .A1_t (new_AGEMA_signal_8667), .A1_f (new_AGEMA_signal_8668), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15), .B0_f (new_AGEMA_signal_8669), .B1_t (new_AGEMA_signal_8670), .B1_f (new_AGEMA_signal_8671), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19), .Z0_f (new_AGEMA_signal_8960), .Z1_t (new_AGEMA_signal_8961), .Z1_f (new_AGEMA_signal_8962) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16), .A0_f (new_AGEMA_signal_8672), .A1_t (new_AGEMA_signal_8673), .A1_f (new_AGEMA_signal_8674), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13), .B0_f (new_AGEMA_signal_8171), .B1_t (new_AGEMA_signal_8172), .B1_f (new_AGEMA_signal_8173), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .Z0_f (new_AGEMA_signal_8963), .Z1_t (new_AGEMA_signal_8964), .Z1_f (new_AGEMA_signal_8965) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17), .A0_f (new_AGEMA_signal_8675), .A1_t (new_AGEMA_signal_8676), .A1_f (new_AGEMA_signal_8677), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15), .B0_f (new_AGEMA_signal_8669), .B1_t (new_AGEMA_signal_8670), .B1_f (new_AGEMA_signal_8671), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .Z0_f (new_AGEMA_signal_8966), .Z1_t (new_AGEMA_signal_8967), .Z1_f (new_AGEMA_signal_8968) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18), .A0_f (new_AGEMA_signal_8678), .A1_t (new_AGEMA_signal_8679), .A1_f (new_AGEMA_signal_8680), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13), .B0_f (new_AGEMA_signal_8171), .B1_t (new_AGEMA_signal_8172), .B1_f (new_AGEMA_signal_8173), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .Z0_f (new_AGEMA_signal_8969), .Z1_t (new_AGEMA_signal_8970), .Z1_f (new_AGEMA_signal_8971) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19), .A0_f (new_AGEMA_signal_8960), .A1_t (new_AGEMA_signal_8961), .A1_f (new_AGEMA_signal_8962), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25), .B0_f (new_AGEMA_signal_8153), .B1_t (new_AGEMA_signal_8154), .B1_f (new_AGEMA_signal_8155), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .Z0_f (new_AGEMA_signal_9200), .Z1_t (new_AGEMA_signal_9201), .Z1_f (new_AGEMA_signal_9202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .A0_f (new_AGEMA_signal_8969), .A1_t (new_AGEMA_signal_8970), .A1_f (new_AGEMA_signal_8971), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .B0_f (new_AGEMA_signal_9200), .B1_t (new_AGEMA_signal_9201), .B1_f (new_AGEMA_signal_9202), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .Z0_f (new_AGEMA_signal_9446), .Z1_t (new_AGEMA_signal_9447), .Z1_f (new_AGEMA_signal_9448) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .A0_f (new_AGEMA_signal_8969), .A1_t (new_AGEMA_signal_8970), .A1_f (new_AGEMA_signal_8971), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .B0_f (new_AGEMA_signal_8963), .B1_t (new_AGEMA_signal_8964), .B1_f (new_AGEMA_signal_8965), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z0_f (new_AGEMA_signal_9203), .Z1_t (new_AGEMA_signal_9204), .Z1_f (new_AGEMA_signal_9205) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .A0_f (new_AGEMA_signal_8966), .A1_t (new_AGEMA_signal_8967), .A1_f (new_AGEMA_signal_8968), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .B0_f (new_AGEMA_signal_9203), .B1_t (new_AGEMA_signal_9204), .B1_f (new_AGEMA_signal_9205), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26), .Z0_f (new_AGEMA_signal_9449), .Z1_t (new_AGEMA_signal_9450), .Z1_f (new_AGEMA_signal_9451) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .A0_f (new_AGEMA_signal_8963), .A1_t (new_AGEMA_signal_8964), .A1_f (new_AGEMA_signal_8965), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .B0_f (new_AGEMA_signal_8966), .B1_t (new_AGEMA_signal_8967), .B1_f (new_AGEMA_signal_8968), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .Z0_f (new_AGEMA_signal_9206), .Z1_t (new_AGEMA_signal_9207), .Z1_f (new_AGEMA_signal_9208) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .A0_f (new_AGEMA_signal_9200), .A1_t (new_AGEMA_signal_9201), .A1_f (new_AGEMA_signal_9202), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .B0_f (new_AGEMA_signal_9203), .B1_t (new_AGEMA_signal_9204), .B1_f (new_AGEMA_signal_9205), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28), .Z0_f (new_AGEMA_signal_9452), .Z1_t (new_AGEMA_signal_9453), .Z1_f (new_AGEMA_signal_9454) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28), .A0_f (new_AGEMA_signal_9452), .A1_t (new_AGEMA_signal_9453), .A1_f (new_AGEMA_signal_9454), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .B0_f (new_AGEMA_signal_9206), .B1_t (new_AGEMA_signal_9207), .B1_f (new_AGEMA_signal_9208), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29), .Z0_f (new_AGEMA_signal_9746), .Z1_t (new_AGEMA_signal_9747), .Z1_f (new_AGEMA_signal_9748) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M30_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26), .A0_f (new_AGEMA_signal_9449), .A1_t (new_AGEMA_signal_9450), .A1_f (new_AGEMA_signal_9451), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .B0_f (new_AGEMA_signal_9446), .B1_t (new_AGEMA_signal_9447), .B1_f (new_AGEMA_signal_9448), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30), .Z0_f (new_AGEMA_signal_9749), .Z1_t (new_AGEMA_signal_9750), .Z1_f (new_AGEMA_signal_9751) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M31_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .A0_f (new_AGEMA_signal_8963), .A1_t (new_AGEMA_signal_8964), .A1_f (new_AGEMA_signal_8965), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .B0_f (new_AGEMA_signal_9200), .B1_t (new_AGEMA_signal_9201), .B1_f (new_AGEMA_signal_9202), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31), .Z0_f (new_AGEMA_signal_9455), .Z1_t (new_AGEMA_signal_9456), .Z1_f (new_AGEMA_signal_9457) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M32_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .A0_f (new_AGEMA_signal_9206), .A1_t (new_AGEMA_signal_9207), .A1_f (new_AGEMA_signal_9208), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31), .B0_f (new_AGEMA_signal_9455), .B1_t (new_AGEMA_signal_9456), .B1_f (new_AGEMA_signal_9457), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32), .Z0_f (new_AGEMA_signal_9752), .Z1_t (new_AGEMA_signal_9753), .Z1_f (new_AGEMA_signal_9754) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M33_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .A0_f (new_AGEMA_signal_9206), .A1_t (new_AGEMA_signal_9207), .A1_f (new_AGEMA_signal_9208), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .B0_f (new_AGEMA_signal_9203), .B1_t (new_AGEMA_signal_9204), .B1_f (new_AGEMA_signal_9205), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33), .Z0_f (new_AGEMA_signal_9458), .Z1_t (new_AGEMA_signal_9459), .Z1_f (new_AGEMA_signal_9460) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M34_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .A0_f (new_AGEMA_signal_8966), .A1_t (new_AGEMA_signal_8967), .A1_f (new_AGEMA_signal_8968), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .B0_f (new_AGEMA_signal_8969), .B1_t (new_AGEMA_signal_8970), .B1_f (new_AGEMA_signal_8971), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34), .Z0_f (new_AGEMA_signal_9209), .Z1_t (new_AGEMA_signal_9210), .Z1_f (new_AGEMA_signal_9211) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M35_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .A0_f (new_AGEMA_signal_9446), .A1_t (new_AGEMA_signal_9447), .A1_f (new_AGEMA_signal_9448), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34), .B0_f (new_AGEMA_signal_9209), .B1_t (new_AGEMA_signal_9210), .B1_f (new_AGEMA_signal_9211), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35), .Z0_f (new_AGEMA_signal_9755), .Z1_t (new_AGEMA_signal_9756), .Z1_f (new_AGEMA_signal_9757) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M36_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .A0_f (new_AGEMA_signal_9446), .A1_t (new_AGEMA_signal_9447), .A1_f (new_AGEMA_signal_9448), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .B0_f (new_AGEMA_signal_9203), .B1_t (new_AGEMA_signal_9204), .B1_f (new_AGEMA_signal_9205), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36), .Z0_f (new_AGEMA_signal_9758), .Z1_t (new_AGEMA_signal_9759), .Z1_f (new_AGEMA_signal_9760) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M37_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .A0_f (new_AGEMA_signal_8966), .A1_t (new_AGEMA_signal_8967), .A1_f (new_AGEMA_signal_8968), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29), .B0_f (new_AGEMA_signal_9746), .B1_t (new_AGEMA_signal_9747), .B1_f (new_AGEMA_signal_9748), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .Z0_f (new_AGEMA_signal_10040), .Z1_t (new_AGEMA_signal_10041), .Z1_f (new_AGEMA_signal_10042) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M38_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32), .A0_f (new_AGEMA_signal_9752), .A1_t (new_AGEMA_signal_9753), .A1_f (new_AGEMA_signal_9754), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33), .B0_f (new_AGEMA_signal_9458), .B1_t (new_AGEMA_signal_9459), .B1_f (new_AGEMA_signal_9460), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .Z0_f (new_AGEMA_signal_10043), .Z1_t (new_AGEMA_signal_10044), .Z1_f (new_AGEMA_signal_10045) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M39_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .A0_f (new_AGEMA_signal_9200), .A1_t (new_AGEMA_signal_9201), .A1_f (new_AGEMA_signal_9202), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30), .B0_f (new_AGEMA_signal_9749), .B1_t (new_AGEMA_signal_9750), .B1_f (new_AGEMA_signal_9751), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .Z0_f (new_AGEMA_signal_10046), .Z1_t (new_AGEMA_signal_10047), .Z1_f (new_AGEMA_signal_10048) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M40_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35), .A0_f (new_AGEMA_signal_9755), .A1_t (new_AGEMA_signal_9756), .A1_f (new_AGEMA_signal_9757), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36), .B0_f (new_AGEMA_signal_9758), .B1_t (new_AGEMA_signal_9759), .B1_f (new_AGEMA_signal_9760), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .Z0_f (new_AGEMA_signal_10049), .Z1_t (new_AGEMA_signal_10050), .Z1_f (new_AGEMA_signal_10051) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M41_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .A0_f (new_AGEMA_signal_10043), .A1_t (new_AGEMA_signal_10044), .A1_f (new_AGEMA_signal_10045), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .B0_f (new_AGEMA_signal_10049), .B1_t (new_AGEMA_signal_10050), .B1_f (new_AGEMA_signal_10051), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .Z0_f (new_AGEMA_signal_10328), .Z1_t (new_AGEMA_signal_10329), .Z1_f (new_AGEMA_signal_10330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M42_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .A0_f (new_AGEMA_signal_10040), .A1_t (new_AGEMA_signal_10041), .A1_f (new_AGEMA_signal_10042), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .B0_f (new_AGEMA_signal_10046), .B1_t (new_AGEMA_signal_10047), .B1_f (new_AGEMA_signal_10048), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .Z0_f (new_AGEMA_signal_10331), .Z1_t (new_AGEMA_signal_10332), .Z1_f (new_AGEMA_signal_10333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M43_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .A0_f (new_AGEMA_signal_10040), .A1_t (new_AGEMA_signal_10041), .A1_f (new_AGEMA_signal_10042), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .B0_f (new_AGEMA_signal_10043), .B1_t (new_AGEMA_signal_10044), .B1_f (new_AGEMA_signal_10045), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43), .Z0_f (new_AGEMA_signal_10334), .Z1_t (new_AGEMA_signal_10335), .Z1_f (new_AGEMA_signal_10336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M44_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .A0_f (new_AGEMA_signal_10046), .A1_t (new_AGEMA_signal_10047), .A1_f (new_AGEMA_signal_10048), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .B0_f (new_AGEMA_signal_10049), .B1_t (new_AGEMA_signal_10050), .B1_f (new_AGEMA_signal_10051), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44), .Z0_f (new_AGEMA_signal_10337), .Z1_t (new_AGEMA_signal_10338), .Z1_f (new_AGEMA_signal_10339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M45_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .A0_f (new_AGEMA_signal_10331), .A1_t (new_AGEMA_signal_10332), .A1_f (new_AGEMA_signal_10333), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .B0_f (new_AGEMA_signal_10328), .B1_t (new_AGEMA_signal_10329), .B1_f (new_AGEMA_signal_10330), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45), .Z0_f (new_AGEMA_signal_11048), .Z1_t (new_AGEMA_signal_11049), .Z1_f (new_AGEMA_signal_11050) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M46_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44), .A0_f (new_AGEMA_signal_10337), .A1_t (new_AGEMA_signal_10338), .A1_f (new_AGEMA_signal_10339), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .B0_f (new_AGEMA_signal_6874), .B1_t (new_AGEMA_signal_6875), .B1_f (new_AGEMA_signal_6876), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46), .Z0_f (new_AGEMA_signal_11051), .Z1_t (new_AGEMA_signal_11052), .Z1_f (new_AGEMA_signal_11053) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M47_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .A0_f (new_AGEMA_signal_10049), .A1_t (new_AGEMA_signal_10050), .A1_f (new_AGEMA_signal_10051), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .B0_f (new_AGEMA_signal_7390), .B1_t (new_AGEMA_signal_7391), .B1_f (new_AGEMA_signal_7392), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47), .Z0_f (new_AGEMA_signal_10340), .Z1_t (new_AGEMA_signal_10341), .Z1_f (new_AGEMA_signal_10342) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M48_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .A0_f (new_AGEMA_signal_10046), .A1_t (new_AGEMA_signal_10047), .A1_f (new_AGEMA_signal_10048), .B0_t (RoundKey[0]), .B0_f (new_AGEMA_signal_5063), .B1_t (new_AGEMA_signal_5064), .B1_f (new_AGEMA_signal_5065), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48), .Z0_f (new_AGEMA_signal_10343), .Z1_t (new_AGEMA_signal_10344), .Z1_f (new_AGEMA_signal_10345) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M49_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43), .A0_f (new_AGEMA_signal_10334), .A1_t (new_AGEMA_signal_10335), .A1_f (new_AGEMA_signal_10336), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .B0_f (new_AGEMA_signal_6886), .B1_t (new_AGEMA_signal_6887), .B1_f (new_AGEMA_signal_6888), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49), .Z0_f (new_AGEMA_signal_11054), .Z1_t (new_AGEMA_signal_11055), .Z1_f (new_AGEMA_signal_11056) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M50_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .A0_f (new_AGEMA_signal_10043), .A1_t (new_AGEMA_signal_10044), .A1_f (new_AGEMA_signal_10045), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .B0_f (new_AGEMA_signal_6877), .B1_t (new_AGEMA_signal_6878), .B1_f (new_AGEMA_signal_6879), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50), .Z0_f (new_AGEMA_signal_10346), .Z1_t (new_AGEMA_signal_10347), .Z1_f (new_AGEMA_signal_10348) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M51_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .A0_f (new_AGEMA_signal_10040), .A1_t (new_AGEMA_signal_10041), .A1_f (new_AGEMA_signal_10042), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .B0_f (new_AGEMA_signal_7399), .B1_t (new_AGEMA_signal_7400), .B1_f (new_AGEMA_signal_7401), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51), .Z0_f (new_AGEMA_signal_10349), .Z1_t (new_AGEMA_signal_10350), .Z1_f (new_AGEMA_signal_10351) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M52_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .A0_f (new_AGEMA_signal_10331), .A1_t (new_AGEMA_signal_10332), .A1_f (new_AGEMA_signal_10333), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .B0_f (new_AGEMA_signal_6883), .B1_t (new_AGEMA_signal_6884), .B1_f (new_AGEMA_signal_6885), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52), .Z0_f (new_AGEMA_signal_11057), .Z1_t (new_AGEMA_signal_11058), .Z1_f (new_AGEMA_signal_11059) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M53_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45), .A0_f (new_AGEMA_signal_11048), .A1_t (new_AGEMA_signal_11049), .A1_f (new_AGEMA_signal_11050), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .B0_f (new_AGEMA_signal_6895), .B1_t (new_AGEMA_signal_6896), .B1_f (new_AGEMA_signal_6897), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53), .Z0_f (new_AGEMA_signal_11756), .Z1_t (new_AGEMA_signal_11757), .Z1_f (new_AGEMA_signal_11758) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M54_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .A0_f (new_AGEMA_signal_10328), .A1_t (new_AGEMA_signal_10329), .A1_f (new_AGEMA_signal_10330), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .B0_f (new_AGEMA_signal_7393), .B1_t (new_AGEMA_signal_7394), .B1_f (new_AGEMA_signal_7395), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54), .Z0_f (new_AGEMA_signal_11060), .Z1_t (new_AGEMA_signal_11061), .Z1_f (new_AGEMA_signal_11062) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M55_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44), .A0_f (new_AGEMA_signal_10337), .A1_t (new_AGEMA_signal_10338), .A1_f (new_AGEMA_signal_10339), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .B0_f (new_AGEMA_signal_6880), .B1_t (new_AGEMA_signal_6881), .B1_f (new_AGEMA_signal_6882), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55), .Z0_f (new_AGEMA_signal_11063), .Z1_t (new_AGEMA_signal_11064), .Z1_f (new_AGEMA_signal_11065) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M56_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .A0_f (new_AGEMA_signal_10049), .A1_t (new_AGEMA_signal_10050), .A1_f (new_AGEMA_signal_10051), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .B0_f (new_AGEMA_signal_7405), .B1_t (new_AGEMA_signal_7406), .B1_f (new_AGEMA_signal_7407), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56), .Z0_f (new_AGEMA_signal_10352), .Z1_t (new_AGEMA_signal_10353), .Z1_f (new_AGEMA_signal_10354) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M57_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .A0_f (new_AGEMA_signal_10046), .A1_t (new_AGEMA_signal_10047), .A1_f (new_AGEMA_signal_10048), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .B0_f (new_AGEMA_signal_6889), .B1_t (new_AGEMA_signal_6890), .B1_f (new_AGEMA_signal_6891), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57), .Z0_f (new_AGEMA_signal_10355), .Z1_t (new_AGEMA_signal_10356), .Z1_f (new_AGEMA_signal_10357) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M58_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43), .A0_f (new_AGEMA_signal_10334), .A1_t (new_AGEMA_signal_10335), .A1_f (new_AGEMA_signal_10336), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .B0_f (new_AGEMA_signal_6279), .B1_t (new_AGEMA_signal_6280), .B1_f (new_AGEMA_signal_6281), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58), .Z0_f (new_AGEMA_signal_11066), .Z1_t (new_AGEMA_signal_11067), .Z1_f (new_AGEMA_signal_11068) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M59_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .A0_f (new_AGEMA_signal_10043), .A1_t (new_AGEMA_signal_10044), .A1_f (new_AGEMA_signal_10045), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .B0_f (new_AGEMA_signal_6892), .B1_t (new_AGEMA_signal_6893), .B1_f (new_AGEMA_signal_6894), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59), .Z0_f (new_AGEMA_signal_10358), .Z1_t (new_AGEMA_signal_10359), .Z1_f (new_AGEMA_signal_10360) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M60_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .A0_f (new_AGEMA_signal_10040), .A1_t (new_AGEMA_signal_10041), .A1_f (new_AGEMA_signal_10042), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .B0_f (new_AGEMA_signal_7402), .B1_t (new_AGEMA_signal_7403), .B1_f (new_AGEMA_signal_7404), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60), .Z0_f (new_AGEMA_signal_10361), .Z1_t (new_AGEMA_signal_10362), .Z1_f (new_AGEMA_signal_10363) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M61_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .A0_f (new_AGEMA_signal_10331), .A1_t (new_AGEMA_signal_10332), .A1_f (new_AGEMA_signal_10333), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .B0_f (new_AGEMA_signal_6273), .B1_t (new_AGEMA_signal_6274), .B1_f (new_AGEMA_signal_6275), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .Z0_f (new_AGEMA_signal_11069), .Z1_t (new_AGEMA_signal_11070), .Z1_f (new_AGEMA_signal_11071) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M62_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45), .A0_f (new_AGEMA_signal_11048), .A1_t (new_AGEMA_signal_11049), .A1_f (new_AGEMA_signal_11050), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .B0_f (new_AGEMA_signal_6282), .B1_t (new_AGEMA_signal_6283), .B1_f (new_AGEMA_signal_6284), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62), .Z0_f (new_AGEMA_signal_11759), .Z1_t (new_AGEMA_signal_11760), .Z1_f (new_AGEMA_signal_11761) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M63_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .A0_f (new_AGEMA_signal_10328), .A1_t (new_AGEMA_signal_10329), .A1_f (new_AGEMA_signal_10330), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .B0_f (new_AGEMA_signal_6276), .B1_t (new_AGEMA_signal_6277), .B1_f (new_AGEMA_signal_6278), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63), .Z0_f (new_AGEMA_signal_11072), .Z1_t (new_AGEMA_signal_11073), .Z1_f (new_AGEMA_signal_11074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .A0_f (new_AGEMA_signal_11069), .A1_t (new_AGEMA_signal_11070), .A1_f (new_AGEMA_signal_11071), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62), .B0_f (new_AGEMA_signal_11759), .B1_t (new_AGEMA_signal_11760), .B1_f (new_AGEMA_signal_11761), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .Z0_f (new_AGEMA_signal_12350), .Z1_t (new_AGEMA_signal_12351), .Z1_f (new_AGEMA_signal_12352) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50), .A0_f (new_AGEMA_signal_10346), .A1_t (new_AGEMA_signal_10347), .A1_f (new_AGEMA_signal_10348), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56), .B0_f (new_AGEMA_signal_10352), .B1_t (new_AGEMA_signal_10353), .B1_f (new_AGEMA_signal_10354), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .Z0_f (new_AGEMA_signal_11075), .Z1_t (new_AGEMA_signal_11076), .Z1_f (new_AGEMA_signal_11077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46), .A0_f (new_AGEMA_signal_11051), .A1_t (new_AGEMA_signal_11052), .A1_f (new_AGEMA_signal_11053), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48), .B0_f (new_AGEMA_signal_10343), .B1_t (new_AGEMA_signal_10344), .B1_f (new_AGEMA_signal_10345), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2), .Z0_f (new_AGEMA_signal_11762), .Z1_t (new_AGEMA_signal_11763), .Z1_f (new_AGEMA_signal_11764) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47), .A0_f (new_AGEMA_signal_10340), .A1_t (new_AGEMA_signal_10341), .A1_f (new_AGEMA_signal_10342), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55), .B0_f (new_AGEMA_signal_11063), .B1_t (new_AGEMA_signal_11064), .B1_f (new_AGEMA_signal_11065), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3), .Z0_f (new_AGEMA_signal_11765), .Z1_t (new_AGEMA_signal_11766), .Z1_f (new_AGEMA_signal_11767) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54), .A0_f (new_AGEMA_signal_11060), .A1_t (new_AGEMA_signal_11061), .A1_f (new_AGEMA_signal_11062), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58), .B0_f (new_AGEMA_signal_11066), .B1_t (new_AGEMA_signal_11067), .B1_f (new_AGEMA_signal_11068), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4), .Z0_f (new_AGEMA_signal_11768), .Z1_t (new_AGEMA_signal_11769), .Z1_f (new_AGEMA_signal_11770) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49), .A0_f (new_AGEMA_signal_11054), .A1_t (new_AGEMA_signal_11055), .A1_f (new_AGEMA_signal_11056), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .B0_f (new_AGEMA_signal_11069), .B1_t (new_AGEMA_signal_11070), .B1_f (new_AGEMA_signal_11071), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5), .Z0_f (new_AGEMA_signal_11771), .Z1_t (new_AGEMA_signal_11772), .Z1_f (new_AGEMA_signal_11773) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62), .A0_f (new_AGEMA_signal_11759), .A1_t (new_AGEMA_signal_11760), .A1_f (new_AGEMA_signal_11761), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5), .B0_f (new_AGEMA_signal_11771), .B1_t (new_AGEMA_signal_11772), .B1_f (new_AGEMA_signal_11773), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .Z0_f (new_AGEMA_signal_12353), .Z1_t (new_AGEMA_signal_12354), .Z1_f (new_AGEMA_signal_12355) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46), .A0_f (new_AGEMA_signal_11051), .A1_t (new_AGEMA_signal_11052), .A1_f (new_AGEMA_signal_11053), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3), .B0_f (new_AGEMA_signal_11765), .B1_t (new_AGEMA_signal_11766), .B1_f (new_AGEMA_signal_11767), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7), .Z0_f (new_AGEMA_signal_12356), .Z1_t (new_AGEMA_signal_12357), .Z1_f (new_AGEMA_signal_12358) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51), .A0_f (new_AGEMA_signal_10349), .A1_t (new_AGEMA_signal_10350), .A1_f (new_AGEMA_signal_10351), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59), .B0_f (new_AGEMA_signal_10358), .B1_t (new_AGEMA_signal_10359), .B1_f (new_AGEMA_signal_10360), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8), .Z0_f (new_AGEMA_signal_11078), .Z1_t (new_AGEMA_signal_11079), .Z1_f (new_AGEMA_signal_11080) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52), .A0_f (new_AGEMA_signal_11057), .A1_t (new_AGEMA_signal_11058), .A1_f (new_AGEMA_signal_11059), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53), .B0_f (new_AGEMA_signal_11756), .B1_t (new_AGEMA_signal_11757), .B1_f (new_AGEMA_signal_11758), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9), .Z0_f (new_AGEMA_signal_12359), .Z1_t (new_AGEMA_signal_12360), .Z1_f (new_AGEMA_signal_12361) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53), .A0_f (new_AGEMA_signal_11756), .A1_t (new_AGEMA_signal_11757), .A1_f (new_AGEMA_signal_11758), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4), .B0_f (new_AGEMA_signal_11768), .B1_t (new_AGEMA_signal_11769), .B1_f (new_AGEMA_signal_11770), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10), .Z0_f (new_AGEMA_signal_12362), .Z1_t (new_AGEMA_signal_12363), .Z1_f (new_AGEMA_signal_12364) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60), .A0_f (new_AGEMA_signal_10361), .A1_t (new_AGEMA_signal_10362), .A1_f (new_AGEMA_signal_10363), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2), .B0_f (new_AGEMA_signal_11762), .B1_t (new_AGEMA_signal_11763), .B1_f (new_AGEMA_signal_11764), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11), .Z0_f (new_AGEMA_signal_12365), .Z1_t (new_AGEMA_signal_12366), .Z1_f (new_AGEMA_signal_12367) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48), .A0_f (new_AGEMA_signal_10343), .A1_t (new_AGEMA_signal_10344), .A1_f (new_AGEMA_signal_10345), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51), .B0_f (new_AGEMA_signal_10349), .B1_t (new_AGEMA_signal_10350), .B1_f (new_AGEMA_signal_10351), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12), .Z0_f (new_AGEMA_signal_11081), .Z1_t (new_AGEMA_signal_11082), .Z1_f (new_AGEMA_signal_11083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50), .A0_f (new_AGEMA_signal_10346), .A1_t (new_AGEMA_signal_10347), .A1_f (new_AGEMA_signal_10348), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .B0_f (new_AGEMA_signal_12350), .B1_t (new_AGEMA_signal_12351), .B1_f (new_AGEMA_signal_12352), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13), .Z0_f (new_AGEMA_signal_12902), .Z1_t (new_AGEMA_signal_12903), .Z1_f (new_AGEMA_signal_12904) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52), .A0_f (new_AGEMA_signal_11057), .A1_t (new_AGEMA_signal_11058), .A1_f (new_AGEMA_signal_11059), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .B0_f (new_AGEMA_signal_11069), .B1_t (new_AGEMA_signal_11070), .B1_f (new_AGEMA_signal_11071), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14), .Z0_f (new_AGEMA_signal_11774), .Z1_t (new_AGEMA_signal_11775), .Z1_f (new_AGEMA_signal_11776) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55), .A0_f (new_AGEMA_signal_11063), .A1_t (new_AGEMA_signal_11064), .A1_f (new_AGEMA_signal_11065), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .B0_f (new_AGEMA_signal_11075), .B1_t (new_AGEMA_signal_11076), .B1_f (new_AGEMA_signal_11077), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15), .Z0_f (new_AGEMA_signal_11777), .Z1_t (new_AGEMA_signal_11778), .Z1_f (new_AGEMA_signal_11779) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56), .A0_f (new_AGEMA_signal_10352), .A1_t (new_AGEMA_signal_10353), .A1_f (new_AGEMA_signal_10354), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .B0_f (new_AGEMA_signal_12350), .B1_t (new_AGEMA_signal_12351), .B1_f (new_AGEMA_signal_12352), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16), .Z0_f (new_AGEMA_signal_12905), .Z1_t (new_AGEMA_signal_12906), .Z1_f (new_AGEMA_signal_12907) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57), .A0_f (new_AGEMA_signal_10355), .A1_t (new_AGEMA_signal_10356), .A1_f (new_AGEMA_signal_10357), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .B0_f (new_AGEMA_signal_11075), .B1_t (new_AGEMA_signal_11076), .B1_f (new_AGEMA_signal_11077), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17), .Z0_f (new_AGEMA_signal_11780), .Z1_t (new_AGEMA_signal_11781), .Z1_f (new_AGEMA_signal_11782) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58), .A0_f (new_AGEMA_signal_11066), .A1_t (new_AGEMA_signal_11067), .A1_f (new_AGEMA_signal_11068), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8), .B0_f (new_AGEMA_signal_11078), .B1_t (new_AGEMA_signal_11079), .B1_f (new_AGEMA_signal_11080), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18), .Z0_f (new_AGEMA_signal_11783), .Z1_t (new_AGEMA_signal_11784), .Z1_f (new_AGEMA_signal_11785) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63), .A0_f (new_AGEMA_signal_11072), .A1_t (new_AGEMA_signal_11073), .A1_f (new_AGEMA_signal_11074), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4), .B0_f (new_AGEMA_signal_11768), .B1_t (new_AGEMA_signal_11769), .B1_f (new_AGEMA_signal_11770), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19), .Z0_f (new_AGEMA_signal_12368), .Z1_t (new_AGEMA_signal_12369), .Z1_f (new_AGEMA_signal_12370) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .A0_f (new_AGEMA_signal_12350), .A1_t (new_AGEMA_signal_12351), .A1_f (new_AGEMA_signal_12352), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .B0_f (new_AGEMA_signal_11075), .B1_t (new_AGEMA_signal_11076), .B1_f (new_AGEMA_signal_11077), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20), .Z0_f (new_AGEMA_signal_12908), .Z1_t (new_AGEMA_signal_12909), .Z1_f (new_AGEMA_signal_12910) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .A0_f (new_AGEMA_signal_11075), .A1_t (new_AGEMA_signal_11076), .A1_f (new_AGEMA_signal_11077), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7), .B0_f (new_AGEMA_signal_12356), .B1_t (new_AGEMA_signal_12357), .B1_f (new_AGEMA_signal_12358), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21), .Z0_f (new_AGEMA_signal_12911), .Z1_t (new_AGEMA_signal_12912), .Z1_f (new_AGEMA_signal_12913) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3), .A0_f (new_AGEMA_signal_11765), .A1_t (new_AGEMA_signal_11766), .A1_f (new_AGEMA_signal_11767), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12), .B0_f (new_AGEMA_signal_11081), .B1_t (new_AGEMA_signal_11082), .B1_f (new_AGEMA_signal_11083), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22), .Z0_f (new_AGEMA_signal_12371), .Z1_t (new_AGEMA_signal_12372), .Z1_f (new_AGEMA_signal_12373) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18), .A0_f (new_AGEMA_signal_11783), .A1_t (new_AGEMA_signal_11784), .A1_f (new_AGEMA_signal_11785), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2), .B0_f (new_AGEMA_signal_11762), .B1_t (new_AGEMA_signal_11763), .B1_f (new_AGEMA_signal_11764), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23), .Z0_f (new_AGEMA_signal_12374), .Z1_t (new_AGEMA_signal_12375), .Z1_f (new_AGEMA_signal_12376) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15), .A0_f (new_AGEMA_signal_11777), .A1_t (new_AGEMA_signal_11778), .A1_f (new_AGEMA_signal_11779), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9), .B0_f (new_AGEMA_signal_12359), .B1_t (new_AGEMA_signal_12360), .B1_f (new_AGEMA_signal_12361), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24), .Z0_f (new_AGEMA_signal_12914), .Z1_t (new_AGEMA_signal_12915), .Z1_f (new_AGEMA_signal_12916) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .A0_f (new_AGEMA_signal_12353), .A1_t (new_AGEMA_signal_12354), .A1_f (new_AGEMA_signal_12355), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10), .B0_f (new_AGEMA_signal_12362), .B1_t (new_AGEMA_signal_12363), .B1_f (new_AGEMA_signal_12364), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25), .Z0_f (new_AGEMA_signal_12917), .Z1_t (new_AGEMA_signal_12918), .Z1_f (new_AGEMA_signal_12919) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7), .A0_f (new_AGEMA_signal_12356), .A1_t (new_AGEMA_signal_12357), .A1_f (new_AGEMA_signal_12358), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9), .B0_f (new_AGEMA_signal_12359), .B1_t (new_AGEMA_signal_12360), .B1_f (new_AGEMA_signal_12361), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26), .Z0_f (new_AGEMA_signal_12920), .Z1_t (new_AGEMA_signal_12921), .Z1_f (new_AGEMA_signal_12922) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8), .A0_f (new_AGEMA_signal_11078), .A1_t (new_AGEMA_signal_11079), .A1_f (new_AGEMA_signal_11080), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10), .B0_f (new_AGEMA_signal_12362), .B1_t (new_AGEMA_signal_12363), .B1_f (new_AGEMA_signal_12364), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27), .Z0_f (new_AGEMA_signal_12923), .Z1_t (new_AGEMA_signal_12924), .Z1_f (new_AGEMA_signal_12925) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11), .A0_f (new_AGEMA_signal_12365), .A1_t (new_AGEMA_signal_12366), .A1_f (new_AGEMA_signal_12367), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14), .B0_f (new_AGEMA_signal_11774), .B1_t (new_AGEMA_signal_11775), .B1_f (new_AGEMA_signal_11776), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28), .Z0_f (new_AGEMA_signal_12926), .Z1_t (new_AGEMA_signal_12927), .Z1_f (new_AGEMA_signal_12928) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11), .A0_f (new_AGEMA_signal_12365), .A1_t (new_AGEMA_signal_12366), .A1_f (new_AGEMA_signal_12367), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17), .B0_f (new_AGEMA_signal_11780), .B1_t (new_AGEMA_signal_11781), .B1_f (new_AGEMA_signal_11782), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29), .Z0_f (new_AGEMA_signal_12929), .Z1_t (new_AGEMA_signal_12930), .Z1_f (new_AGEMA_signal_12931) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .A0_f (new_AGEMA_signal_12353), .A1_t (new_AGEMA_signal_12354), .A1_f (new_AGEMA_signal_12355), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24), .B0_f (new_AGEMA_signal_12914), .B1_t (new_AGEMA_signal_12915), .B1_f (new_AGEMA_signal_12916), .Z0_t (KeyExpansionIns_tmp[15]), .Z0_f (new_AGEMA_signal_13550), .Z1_t (new_AGEMA_signal_13551), .Z1_f (new_AGEMA_signal_13552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16), .A0_f (new_AGEMA_signal_12905), .A1_t (new_AGEMA_signal_12906), .A1_f (new_AGEMA_signal_12907), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26), .B0_f (new_AGEMA_signal_12920), .B1_t (new_AGEMA_signal_12921), .B1_f (new_AGEMA_signal_12922), .Z0_t (KeyExpansionIns_tmp[14]), .Z0_f (new_AGEMA_signal_13553), .Z1_t (new_AGEMA_signal_13554), .Z1_f (new_AGEMA_signal_13555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19), .A0_f (new_AGEMA_signal_12368), .A1_t (new_AGEMA_signal_12369), .A1_f (new_AGEMA_signal_12370), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28), .B0_f (new_AGEMA_signal_12926), .B1_t (new_AGEMA_signal_12927), .B1_f (new_AGEMA_signal_12928), .Z0_t (KeyExpansionIns_tmp[13]), .Z0_f (new_AGEMA_signal_13556), .Z1_t (new_AGEMA_signal_13557), .Z1_f (new_AGEMA_signal_13558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .A0_f (new_AGEMA_signal_12353), .A1_t (new_AGEMA_signal_12354), .A1_f (new_AGEMA_signal_12355), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21), .B0_f (new_AGEMA_signal_12911), .B1_t (new_AGEMA_signal_12912), .B1_f (new_AGEMA_signal_12913), .Z0_t (KeyExpansionIns_tmp[12]), .Z0_f (new_AGEMA_signal_13559), .Z1_t (new_AGEMA_signal_13560), .Z1_f (new_AGEMA_signal_13561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20), .A0_f (new_AGEMA_signal_12908), .A1_t (new_AGEMA_signal_12909), .A1_f (new_AGEMA_signal_12910), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22), .B0_f (new_AGEMA_signal_12371), .B1_t (new_AGEMA_signal_12372), .B1_f (new_AGEMA_signal_12373), .Z0_t (KeyExpansionIns_tmp[11]), .Z0_f (new_AGEMA_signal_13562), .Z1_t (new_AGEMA_signal_13563), .Z1_f (new_AGEMA_signal_13564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25), .A0_f (new_AGEMA_signal_12917), .A1_t (new_AGEMA_signal_12918), .A1_f (new_AGEMA_signal_12919), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29), .B0_f (new_AGEMA_signal_12929), .B1_t (new_AGEMA_signal_12930), .B1_f (new_AGEMA_signal_12931), .Z0_t (KeyExpansionIns_tmp[10]), .Z0_f (new_AGEMA_signal_13565), .Z1_t (new_AGEMA_signal_13566), .Z1_f (new_AGEMA_signal_13567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13), .A0_f (new_AGEMA_signal_12902), .A1_t (new_AGEMA_signal_12903), .A1_f (new_AGEMA_signal_12904), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27), .B0_f (new_AGEMA_signal_12923), .B1_t (new_AGEMA_signal_12924), .B1_f (new_AGEMA_signal_12925), .Z0_t (KeyExpansionIns_tmp[9]), .Z0_f (new_AGEMA_signal_13568), .Z1_t (new_AGEMA_signal_13569), .Z1_f (new_AGEMA_signal_13570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .A0_f (new_AGEMA_signal_12353), .A1_t (new_AGEMA_signal_12354), .A1_f (new_AGEMA_signal_12355), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23), .B0_f (new_AGEMA_signal_12374), .B1_t (new_AGEMA_signal_12375), .B1_f (new_AGEMA_signal_12376), .Z0_t (KeyExpansionIns_tmp[8]), .Z0_f (new_AGEMA_signal_12932), .Z1_t (new_AGEMA_signal_12933), .Z1_f (new_AGEMA_signal_12934) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T1_U1 ( .A0_t (RoundKey[31]), .A0_f (new_AGEMA_signal_5531), .A1_t (new_AGEMA_signal_5532), .A1_f (new_AGEMA_signal_5533), .B0_t (RoundKey[28]), .B0_f (new_AGEMA_signal_5495), .B1_t (new_AGEMA_signal_5496), .B1_f (new_AGEMA_signal_5497), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .Z0_f (new_AGEMA_signal_6303), .Z1_t (new_AGEMA_signal_6304), .Z1_f (new_AGEMA_signal_6305) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T2_U1 ( .A0_t (RoundKey[31]), .A0_f (new_AGEMA_signal_5531), .A1_t (new_AGEMA_signal_5532), .A1_f (new_AGEMA_signal_5533), .B0_t (RoundKey[26]), .B0_f (new_AGEMA_signal_5477), .B1_t (new_AGEMA_signal_5478), .B1_f (new_AGEMA_signal_5479), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .Z0_f (new_AGEMA_signal_6306), .Z1_t (new_AGEMA_signal_6307), .Z1_f (new_AGEMA_signal_6308) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T3_U1 ( .A0_t (RoundKey[31]), .A0_f (new_AGEMA_signal_5531), .A1_t (new_AGEMA_signal_5532), .A1_f (new_AGEMA_signal_5533), .B0_t (RoundKey[25]), .B0_f (new_AGEMA_signal_5468), .B1_t (new_AGEMA_signal_5469), .B1_f (new_AGEMA_signal_5470), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .Z0_f (new_AGEMA_signal_6309), .Z1_t (new_AGEMA_signal_6310), .Z1_f (new_AGEMA_signal_6311) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T4_U1 ( .A0_t (RoundKey[28]), .A0_f (new_AGEMA_signal_5495), .A1_t (new_AGEMA_signal_5496), .A1_f (new_AGEMA_signal_5497), .B0_t (RoundKey[26]), .B0_f (new_AGEMA_signal_5477), .B1_t (new_AGEMA_signal_5478), .B1_f (new_AGEMA_signal_5479), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .Z0_f (new_AGEMA_signal_6312), .Z1_t (new_AGEMA_signal_6313), .Z1_f (new_AGEMA_signal_6314) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T5_U1 ( .A0_t (RoundKey[27]), .A0_f (new_AGEMA_signal_5486), .A1_t (new_AGEMA_signal_5487), .A1_f (new_AGEMA_signal_5488), .B0_t (RoundKey[25]), .B0_f (new_AGEMA_signal_5468), .B1_t (new_AGEMA_signal_5469), .B1_f (new_AGEMA_signal_5470), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .Z0_f (new_AGEMA_signal_6315), .Z1_t (new_AGEMA_signal_6316), .Z1_f (new_AGEMA_signal_6317) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .A0_f (new_AGEMA_signal_6303), .A1_t (new_AGEMA_signal_6304), .A1_f (new_AGEMA_signal_6305), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .B0_f (new_AGEMA_signal_6315), .B1_t (new_AGEMA_signal_6316), .B1_f (new_AGEMA_signal_6317), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .Z0_f (new_AGEMA_signal_6898), .Z1_t (new_AGEMA_signal_6899), .Z1_f (new_AGEMA_signal_6900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T7_U1 ( .A0_t (RoundKey[30]), .A0_f (new_AGEMA_signal_5522), .A1_t (new_AGEMA_signal_5523), .A1_f (new_AGEMA_signal_5524), .B0_t (RoundKey[29]), .B0_f (new_AGEMA_signal_5504), .B1_t (new_AGEMA_signal_5505), .B1_f (new_AGEMA_signal_5506), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .Z0_f (new_AGEMA_signal_6318), .Z1_t (new_AGEMA_signal_6319), .Z1_f (new_AGEMA_signal_6320) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T8_U1 ( .A0_t (RoundKey[24]), .A0_f (new_AGEMA_signal_5459), .A1_t (new_AGEMA_signal_5460), .A1_f (new_AGEMA_signal_5461), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .B0_f (new_AGEMA_signal_6898), .B1_t (new_AGEMA_signal_6899), .B1_f (new_AGEMA_signal_6900), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .Z0_f (new_AGEMA_signal_7429), .Z1_t (new_AGEMA_signal_7430), .Z1_f (new_AGEMA_signal_7431) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T9_U1 ( .A0_t (RoundKey[24]), .A0_f (new_AGEMA_signal_5459), .A1_t (new_AGEMA_signal_5460), .A1_f (new_AGEMA_signal_5461), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .B0_f (new_AGEMA_signal_6318), .B1_t (new_AGEMA_signal_6319), .B1_f (new_AGEMA_signal_6320), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .Z0_f (new_AGEMA_signal_6901), .Z1_t (new_AGEMA_signal_6902), .Z1_f (new_AGEMA_signal_6903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .A0_f (new_AGEMA_signal_6898), .A1_t (new_AGEMA_signal_6899), .A1_f (new_AGEMA_signal_6900), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .B0_f (new_AGEMA_signal_6318), .B1_t (new_AGEMA_signal_6319), .B1_f (new_AGEMA_signal_6320), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .Z0_f (new_AGEMA_signal_7432), .Z1_t (new_AGEMA_signal_7433), .Z1_f (new_AGEMA_signal_7434) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T11_U1 ( .A0_t (RoundKey[30]), .A0_f (new_AGEMA_signal_5522), .A1_t (new_AGEMA_signal_5523), .A1_f (new_AGEMA_signal_5524), .B0_t (RoundKey[26]), .B0_f (new_AGEMA_signal_5477), .B1_t (new_AGEMA_signal_5478), .B1_f (new_AGEMA_signal_5479), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11), .Z0_f (new_AGEMA_signal_6321), .Z1_t (new_AGEMA_signal_6322), .Z1_f (new_AGEMA_signal_6323) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T12_U1 ( .A0_t (RoundKey[29]), .A0_f (new_AGEMA_signal_5504), .A1_t (new_AGEMA_signal_5505), .A1_f (new_AGEMA_signal_5506), .B0_t (RoundKey[26]), .B0_f (new_AGEMA_signal_5477), .B1_t (new_AGEMA_signal_5478), .B1_f (new_AGEMA_signal_5479), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12), .Z0_f (new_AGEMA_signal_6324), .Z1_t (new_AGEMA_signal_6325), .Z1_f (new_AGEMA_signal_6326) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .A0_f (new_AGEMA_signal_6309), .A1_t (new_AGEMA_signal_6310), .A1_f (new_AGEMA_signal_6311), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .B0_f (new_AGEMA_signal_6312), .B1_t (new_AGEMA_signal_6313), .B1_f (new_AGEMA_signal_6314), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .Z0_f (new_AGEMA_signal_6904), .Z1_t (new_AGEMA_signal_6905), .Z1_f (new_AGEMA_signal_6906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .A0_f (new_AGEMA_signal_6898), .A1_t (new_AGEMA_signal_6899), .A1_f (new_AGEMA_signal_6900), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11), .B0_f (new_AGEMA_signal_6321), .B1_t (new_AGEMA_signal_6322), .B1_f (new_AGEMA_signal_6323), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14), .Z0_f (new_AGEMA_signal_7435), .Z1_t (new_AGEMA_signal_7436), .Z1_f (new_AGEMA_signal_7437) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .A0_f (new_AGEMA_signal_6315), .A1_t (new_AGEMA_signal_6316), .A1_f (new_AGEMA_signal_6317), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11), .B0_f (new_AGEMA_signal_6321), .B1_t (new_AGEMA_signal_6322), .B1_f (new_AGEMA_signal_6323), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .Z0_f (new_AGEMA_signal_6907), .Z1_t (new_AGEMA_signal_6908), .Z1_f (new_AGEMA_signal_6909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .A0_f (new_AGEMA_signal_6315), .A1_t (new_AGEMA_signal_6316), .A1_f (new_AGEMA_signal_6317), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12), .B0_f (new_AGEMA_signal_6324), .B1_t (new_AGEMA_signal_6325), .B1_f (new_AGEMA_signal_6326), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Z0_f (new_AGEMA_signal_6910), .Z1_t (new_AGEMA_signal_6911), .Z1_f (new_AGEMA_signal_6912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .A0_f (new_AGEMA_signal_6901), .A1_t (new_AGEMA_signal_6902), .A1_f (new_AGEMA_signal_6903), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .B0_f (new_AGEMA_signal_6910), .B1_t (new_AGEMA_signal_6911), .B1_f (new_AGEMA_signal_6912), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .Z0_f (new_AGEMA_signal_7438), .Z1_t (new_AGEMA_signal_7439), .Z1_f (new_AGEMA_signal_7440) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T18_U1 ( .A0_t (RoundKey[28]), .A0_f (new_AGEMA_signal_5495), .A1_t (new_AGEMA_signal_5496), .A1_f (new_AGEMA_signal_5497), .B0_t (RoundKey[24]), .B0_f (new_AGEMA_signal_5459), .B1_t (new_AGEMA_signal_5460), .B1_f (new_AGEMA_signal_5461), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18), .Z0_f (new_AGEMA_signal_6327), .Z1_t (new_AGEMA_signal_6328), .Z1_f (new_AGEMA_signal_6329) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .A0_f (new_AGEMA_signal_6318), .A1_t (new_AGEMA_signal_6319), .A1_f (new_AGEMA_signal_6320), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18), .B0_f (new_AGEMA_signal_6327), .B1_t (new_AGEMA_signal_6328), .B1_f (new_AGEMA_signal_6329), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .Z0_f (new_AGEMA_signal_6913), .Z1_t (new_AGEMA_signal_6914), .Z1_f (new_AGEMA_signal_6915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .A0_f (new_AGEMA_signal_6303), .A1_t (new_AGEMA_signal_6304), .A1_f (new_AGEMA_signal_6305), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .B0_f (new_AGEMA_signal_6913), .B1_t (new_AGEMA_signal_6914), .B1_f (new_AGEMA_signal_6915), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .Z0_f (new_AGEMA_signal_7441), .Z1_t (new_AGEMA_signal_7442), .Z1_f (new_AGEMA_signal_7443) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T21_U1 ( .A0_t (RoundKey[25]), .A0_f (new_AGEMA_signal_5468), .A1_t (new_AGEMA_signal_5469), .A1_f (new_AGEMA_signal_5470), .B0_t (RoundKey[24]), .B0_f (new_AGEMA_signal_5459), .B1_t (new_AGEMA_signal_5460), .B1_f (new_AGEMA_signal_5461), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21), .Z0_f (new_AGEMA_signal_6330), .Z1_t (new_AGEMA_signal_6331), .Z1_f (new_AGEMA_signal_6332) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .A0_f (new_AGEMA_signal_6318), .A1_t (new_AGEMA_signal_6319), .A1_f (new_AGEMA_signal_6320), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21), .B0_f (new_AGEMA_signal_6330), .B1_t (new_AGEMA_signal_6331), .B1_f (new_AGEMA_signal_6332), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .Z0_f (new_AGEMA_signal_6916), .Z1_t (new_AGEMA_signal_6917), .Z1_f (new_AGEMA_signal_6918) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .A0_f (new_AGEMA_signal_6306), .A1_t (new_AGEMA_signal_6307), .A1_f (new_AGEMA_signal_6308), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .B0_f (new_AGEMA_signal_6916), .B1_t (new_AGEMA_signal_6917), .B1_f (new_AGEMA_signal_6918), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .Z0_f (new_AGEMA_signal_7444), .Z1_t (new_AGEMA_signal_7445), .Z1_f (new_AGEMA_signal_7446) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .A0_f (new_AGEMA_signal_6306), .A1_t (new_AGEMA_signal_6307), .A1_f (new_AGEMA_signal_6308), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .B0_f (new_AGEMA_signal_7432), .B1_t (new_AGEMA_signal_7433), .B1_f (new_AGEMA_signal_7434), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24), .Z0_f (new_AGEMA_signal_8177), .Z1_t (new_AGEMA_signal_8178), .Z1_f (new_AGEMA_signal_8179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .A0_f (new_AGEMA_signal_7441), .A1_t (new_AGEMA_signal_7442), .A1_f (new_AGEMA_signal_7443), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .B0_f (new_AGEMA_signal_7438), .B1_t (new_AGEMA_signal_7439), .B1_f (new_AGEMA_signal_7440), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25), .Z0_f (new_AGEMA_signal_8180), .Z1_t (new_AGEMA_signal_8181), .Z1_f (new_AGEMA_signal_8182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .A0_f (new_AGEMA_signal_6309), .A1_t (new_AGEMA_signal_6310), .A1_f (new_AGEMA_signal_6311), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .B0_f (new_AGEMA_signal_6910), .B1_t (new_AGEMA_signal_6911), .B1_f (new_AGEMA_signal_6912), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26), .Z0_f (new_AGEMA_signal_7447), .Z1_t (new_AGEMA_signal_7448), .Z1_f (new_AGEMA_signal_7449) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .A0_f (new_AGEMA_signal_6303), .A1_t (new_AGEMA_signal_6304), .A1_f (new_AGEMA_signal_6305), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12), .B0_f (new_AGEMA_signal_6324), .B1_t (new_AGEMA_signal_6325), .B1_f (new_AGEMA_signal_6326), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .Z0_f (new_AGEMA_signal_6919), .Z1_t (new_AGEMA_signal_6920), .Z1_f (new_AGEMA_signal_6921) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .A0_f (new_AGEMA_signal_6904), .A1_t (new_AGEMA_signal_6905), .A1_f (new_AGEMA_signal_6906), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .B0_f (new_AGEMA_signal_6898), .B1_t (new_AGEMA_signal_6899), .B1_f (new_AGEMA_signal_6900), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1), .Z0_f (new_AGEMA_signal_7450), .Z1_t (new_AGEMA_signal_7451), .Z1_f (new_AGEMA_signal_7452) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .A0_f (new_AGEMA_signal_7444), .A1_t (new_AGEMA_signal_7445), .A1_f (new_AGEMA_signal_7446), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .B0_f (new_AGEMA_signal_7429), .B1_t (new_AGEMA_signal_7430), .B1_f (new_AGEMA_signal_7431), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2), .Z0_f (new_AGEMA_signal_8183), .Z1_t (new_AGEMA_signal_8184), .Z1_f (new_AGEMA_signal_8185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14), .A0_f (new_AGEMA_signal_7435), .A1_t (new_AGEMA_signal_7436), .A1_f (new_AGEMA_signal_7437), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1), .B0_f (new_AGEMA_signal_7450), .B1_t (new_AGEMA_signal_7451), .B1_f (new_AGEMA_signal_7452), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3), .Z0_f (new_AGEMA_signal_8186), .Z1_t (new_AGEMA_signal_8187), .Z1_f (new_AGEMA_signal_8188) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .A0_f (new_AGEMA_signal_6913), .A1_t (new_AGEMA_signal_6914), .A1_f (new_AGEMA_signal_6915), .B0_t (RoundKey[24]), .B0_f (new_AGEMA_signal_5459), .B1_t (new_AGEMA_signal_5460), .B1_f (new_AGEMA_signal_5461), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4), .Z0_f (new_AGEMA_signal_7453), .Z1_t (new_AGEMA_signal_7454), .Z1_f (new_AGEMA_signal_7455) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4), .A0_f (new_AGEMA_signal_7453), .A1_t (new_AGEMA_signal_7454), .A1_f (new_AGEMA_signal_7455), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1), .B0_f (new_AGEMA_signal_7450), .B1_t (new_AGEMA_signal_7451), .B1_f (new_AGEMA_signal_7452), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5), .Z0_f (new_AGEMA_signal_8189), .Z1_t (new_AGEMA_signal_8190), .Z1_f (new_AGEMA_signal_8191) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .A0_f (new_AGEMA_signal_6309), .A1_t (new_AGEMA_signal_6310), .A1_f (new_AGEMA_signal_6311), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .B0_f (new_AGEMA_signal_6910), .B1_t (new_AGEMA_signal_6911), .B1_f (new_AGEMA_signal_6912), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6), .Z0_f (new_AGEMA_signal_7456), .Z1_t (new_AGEMA_signal_7457), .Z1_f (new_AGEMA_signal_7458) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .A0_f (new_AGEMA_signal_6916), .A1_t (new_AGEMA_signal_6917), .A1_f (new_AGEMA_signal_6918), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .B0_f (new_AGEMA_signal_6901), .B1_t (new_AGEMA_signal_6902), .B1_f (new_AGEMA_signal_6903), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7), .Z0_f (new_AGEMA_signal_7459), .Z1_t (new_AGEMA_signal_7460), .Z1_f (new_AGEMA_signal_7461) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26), .A0_f (new_AGEMA_signal_7447), .A1_t (new_AGEMA_signal_7448), .A1_f (new_AGEMA_signal_7449), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6), .B0_f (new_AGEMA_signal_7456), .B1_t (new_AGEMA_signal_7457), .B1_f (new_AGEMA_signal_7458), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8), .Z0_f (new_AGEMA_signal_8192), .Z1_t (new_AGEMA_signal_8193), .Z1_f (new_AGEMA_signal_8194) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .A0_f (new_AGEMA_signal_7441), .A1_t (new_AGEMA_signal_7442), .A1_f (new_AGEMA_signal_7443), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .B0_f (new_AGEMA_signal_7438), .B1_t (new_AGEMA_signal_7439), .B1_f (new_AGEMA_signal_7440), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9), .Z0_f (new_AGEMA_signal_8195), .Z1_t (new_AGEMA_signal_8196), .Z1_f (new_AGEMA_signal_8197) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9), .A0_f (new_AGEMA_signal_8195), .A1_t (new_AGEMA_signal_8196), .A1_f (new_AGEMA_signal_8197), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6), .B0_f (new_AGEMA_signal_7456), .B1_t (new_AGEMA_signal_7457), .B1_f (new_AGEMA_signal_7458), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10), .Z0_f (new_AGEMA_signal_8681), .Z1_t (new_AGEMA_signal_8682), .Z1_f (new_AGEMA_signal_8683) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .A0_f (new_AGEMA_signal_6303), .A1_t (new_AGEMA_signal_6304), .A1_f (new_AGEMA_signal_6305), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .B0_f (new_AGEMA_signal_6907), .B1_t (new_AGEMA_signal_6908), .B1_f (new_AGEMA_signal_6909), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11), .Z0_f (new_AGEMA_signal_7462), .Z1_t (new_AGEMA_signal_7463), .Z1_f (new_AGEMA_signal_7464) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .A0_f (new_AGEMA_signal_6312), .A1_t (new_AGEMA_signal_6313), .A1_f (new_AGEMA_signal_6314), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .B0_f (new_AGEMA_signal_6919), .B1_t (new_AGEMA_signal_6920), .B1_f (new_AGEMA_signal_6921), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12), .Z0_f (new_AGEMA_signal_7465), .Z1_t (new_AGEMA_signal_7466), .Z1_f (new_AGEMA_signal_7467) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12), .A0_f (new_AGEMA_signal_7465), .A1_t (new_AGEMA_signal_7466), .A1_f (new_AGEMA_signal_7467), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11), .B0_f (new_AGEMA_signal_7462), .B1_t (new_AGEMA_signal_7463), .B1_f (new_AGEMA_signal_7464), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13), .Z0_f (new_AGEMA_signal_8198), .Z1_t (new_AGEMA_signal_8199), .Z1_f (new_AGEMA_signal_8200) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .A0_f (new_AGEMA_signal_6306), .A1_t (new_AGEMA_signal_6307), .A1_f (new_AGEMA_signal_6308), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .B0_f (new_AGEMA_signal_7432), .B1_t (new_AGEMA_signal_7433), .B1_f (new_AGEMA_signal_7434), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14), .Z0_f (new_AGEMA_signal_8201), .Z1_t (new_AGEMA_signal_8202), .Z1_f (new_AGEMA_signal_8203) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14), .A0_f (new_AGEMA_signal_8201), .A1_t (new_AGEMA_signal_8202), .A1_f (new_AGEMA_signal_8203), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11), .B0_f (new_AGEMA_signal_7462), .B1_t (new_AGEMA_signal_7463), .B1_f (new_AGEMA_signal_7464), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15), .Z0_f (new_AGEMA_signal_8684), .Z1_t (new_AGEMA_signal_8685), .Z1_f (new_AGEMA_signal_8686) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3), .A0_f (new_AGEMA_signal_8186), .A1_t (new_AGEMA_signal_8187), .A1_f (new_AGEMA_signal_8188), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2), .B0_f (new_AGEMA_signal_8183), .B1_t (new_AGEMA_signal_8184), .B1_f (new_AGEMA_signal_8185), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16), .Z0_f (new_AGEMA_signal_8687), .Z1_t (new_AGEMA_signal_8688), .Z1_f (new_AGEMA_signal_8689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5), .A0_f (new_AGEMA_signal_8189), .A1_t (new_AGEMA_signal_8190), .A1_f (new_AGEMA_signal_8191), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24), .B0_f (new_AGEMA_signal_8177), .B1_t (new_AGEMA_signal_8178), .B1_f (new_AGEMA_signal_8179), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17), .Z0_f (new_AGEMA_signal_8690), .Z1_t (new_AGEMA_signal_8691), .Z1_f (new_AGEMA_signal_8692) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8), .A0_f (new_AGEMA_signal_8192), .A1_t (new_AGEMA_signal_8193), .A1_f (new_AGEMA_signal_8194), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7), .B0_f (new_AGEMA_signal_7459), .B1_t (new_AGEMA_signal_7460), .B1_f (new_AGEMA_signal_7461), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18), .Z0_f (new_AGEMA_signal_8693), .Z1_t (new_AGEMA_signal_8694), .Z1_f (new_AGEMA_signal_8695) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10), .A0_f (new_AGEMA_signal_8681), .A1_t (new_AGEMA_signal_8682), .A1_f (new_AGEMA_signal_8683), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15), .B0_f (new_AGEMA_signal_8684), .B1_t (new_AGEMA_signal_8685), .B1_f (new_AGEMA_signal_8686), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19), .Z0_f (new_AGEMA_signal_8972), .Z1_t (new_AGEMA_signal_8973), .Z1_f (new_AGEMA_signal_8974) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16), .A0_f (new_AGEMA_signal_8687), .A1_t (new_AGEMA_signal_8688), .A1_f (new_AGEMA_signal_8689), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13), .B0_f (new_AGEMA_signal_8198), .B1_t (new_AGEMA_signal_8199), .B1_f (new_AGEMA_signal_8200), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .Z0_f (new_AGEMA_signal_8975), .Z1_t (new_AGEMA_signal_8976), .Z1_f (new_AGEMA_signal_8977) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17), .A0_f (new_AGEMA_signal_8690), .A1_t (new_AGEMA_signal_8691), .A1_f (new_AGEMA_signal_8692), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15), .B0_f (new_AGEMA_signal_8684), .B1_t (new_AGEMA_signal_8685), .B1_f (new_AGEMA_signal_8686), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .Z0_f (new_AGEMA_signal_8978), .Z1_t (new_AGEMA_signal_8979), .Z1_f (new_AGEMA_signal_8980) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18), .A0_f (new_AGEMA_signal_8693), .A1_t (new_AGEMA_signal_8694), .A1_f (new_AGEMA_signal_8695), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13), .B0_f (new_AGEMA_signal_8198), .B1_t (new_AGEMA_signal_8199), .B1_f (new_AGEMA_signal_8200), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .Z0_f (new_AGEMA_signal_8981), .Z1_t (new_AGEMA_signal_8982), .Z1_f (new_AGEMA_signal_8983) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19), .A0_f (new_AGEMA_signal_8972), .A1_t (new_AGEMA_signal_8973), .A1_f (new_AGEMA_signal_8974), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25), .B0_f (new_AGEMA_signal_8180), .B1_t (new_AGEMA_signal_8181), .B1_f (new_AGEMA_signal_8182), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .Z0_f (new_AGEMA_signal_9212), .Z1_t (new_AGEMA_signal_9213), .Z1_f (new_AGEMA_signal_9214) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .A0_f (new_AGEMA_signal_8981), .A1_t (new_AGEMA_signal_8982), .A1_f (new_AGEMA_signal_8983), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .B0_f (new_AGEMA_signal_9212), .B1_t (new_AGEMA_signal_9213), .B1_f (new_AGEMA_signal_9214), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .Z0_f (new_AGEMA_signal_9461), .Z1_t (new_AGEMA_signal_9462), .Z1_f (new_AGEMA_signal_9463) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .A0_f (new_AGEMA_signal_8981), .A1_t (new_AGEMA_signal_8982), .A1_f (new_AGEMA_signal_8983), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .B0_f (new_AGEMA_signal_8975), .B1_t (new_AGEMA_signal_8976), .B1_f (new_AGEMA_signal_8977), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z0_f (new_AGEMA_signal_9215), .Z1_t (new_AGEMA_signal_9216), .Z1_f (new_AGEMA_signal_9217) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .A0_f (new_AGEMA_signal_8978), .A1_t (new_AGEMA_signal_8979), .A1_f (new_AGEMA_signal_8980), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .B0_f (new_AGEMA_signal_9215), .B1_t (new_AGEMA_signal_9216), .B1_f (new_AGEMA_signal_9217), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26), .Z0_f (new_AGEMA_signal_9464), .Z1_t (new_AGEMA_signal_9465), .Z1_f (new_AGEMA_signal_9466) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .A0_f (new_AGEMA_signal_8975), .A1_t (new_AGEMA_signal_8976), .A1_f (new_AGEMA_signal_8977), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .B0_f (new_AGEMA_signal_8978), .B1_t (new_AGEMA_signal_8979), .B1_f (new_AGEMA_signal_8980), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .Z0_f (new_AGEMA_signal_9218), .Z1_t (new_AGEMA_signal_9219), .Z1_f (new_AGEMA_signal_9220) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .A0_f (new_AGEMA_signal_9212), .A1_t (new_AGEMA_signal_9213), .A1_f (new_AGEMA_signal_9214), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .B0_f (new_AGEMA_signal_9215), .B1_t (new_AGEMA_signal_9216), .B1_f (new_AGEMA_signal_9217), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28), .Z0_f (new_AGEMA_signal_9467), .Z1_t (new_AGEMA_signal_9468), .Z1_f (new_AGEMA_signal_9469) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28), .A0_f (new_AGEMA_signal_9467), .A1_t (new_AGEMA_signal_9468), .A1_f (new_AGEMA_signal_9469), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .B0_f (new_AGEMA_signal_9218), .B1_t (new_AGEMA_signal_9219), .B1_f (new_AGEMA_signal_9220), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29), .Z0_f (new_AGEMA_signal_9761), .Z1_t (new_AGEMA_signal_9762), .Z1_f (new_AGEMA_signal_9763) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M30_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26), .A0_f (new_AGEMA_signal_9464), .A1_t (new_AGEMA_signal_9465), .A1_f (new_AGEMA_signal_9466), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .B0_f (new_AGEMA_signal_9461), .B1_t (new_AGEMA_signal_9462), .B1_f (new_AGEMA_signal_9463), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30), .Z0_f (new_AGEMA_signal_9764), .Z1_t (new_AGEMA_signal_9765), .Z1_f (new_AGEMA_signal_9766) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M31_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .A0_f (new_AGEMA_signal_8975), .A1_t (new_AGEMA_signal_8976), .A1_f (new_AGEMA_signal_8977), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .B0_f (new_AGEMA_signal_9212), .B1_t (new_AGEMA_signal_9213), .B1_f (new_AGEMA_signal_9214), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31), .Z0_f (new_AGEMA_signal_9470), .Z1_t (new_AGEMA_signal_9471), .Z1_f (new_AGEMA_signal_9472) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M32_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .A0_f (new_AGEMA_signal_9218), .A1_t (new_AGEMA_signal_9219), .A1_f (new_AGEMA_signal_9220), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31), .B0_f (new_AGEMA_signal_9470), .B1_t (new_AGEMA_signal_9471), .B1_f (new_AGEMA_signal_9472), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32), .Z0_f (new_AGEMA_signal_9767), .Z1_t (new_AGEMA_signal_9768), .Z1_f (new_AGEMA_signal_9769) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M33_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .A0_f (new_AGEMA_signal_9218), .A1_t (new_AGEMA_signal_9219), .A1_f (new_AGEMA_signal_9220), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .B0_f (new_AGEMA_signal_9215), .B1_t (new_AGEMA_signal_9216), .B1_f (new_AGEMA_signal_9217), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33), .Z0_f (new_AGEMA_signal_9473), .Z1_t (new_AGEMA_signal_9474), .Z1_f (new_AGEMA_signal_9475) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M34_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .A0_f (new_AGEMA_signal_8978), .A1_t (new_AGEMA_signal_8979), .A1_f (new_AGEMA_signal_8980), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .B0_f (new_AGEMA_signal_8981), .B1_t (new_AGEMA_signal_8982), .B1_f (new_AGEMA_signal_8983), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34), .Z0_f (new_AGEMA_signal_9221), .Z1_t (new_AGEMA_signal_9222), .Z1_f (new_AGEMA_signal_9223) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M35_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .A0_f (new_AGEMA_signal_9461), .A1_t (new_AGEMA_signal_9462), .A1_f (new_AGEMA_signal_9463), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34), .B0_f (new_AGEMA_signal_9221), .B1_t (new_AGEMA_signal_9222), .B1_f (new_AGEMA_signal_9223), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35), .Z0_f (new_AGEMA_signal_9770), .Z1_t (new_AGEMA_signal_9771), .Z1_f (new_AGEMA_signal_9772) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M36_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .A0_f (new_AGEMA_signal_9461), .A1_t (new_AGEMA_signal_9462), .A1_f (new_AGEMA_signal_9463), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .B0_f (new_AGEMA_signal_9215), .B1_t (new_AGEMA_signal_9216), .B1_f (new_AGEMA_signal_9217), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36), .Z0_f (new_AGEMA_signal_9773), .Z1_t (new_AGEMA_signal_9774), .Z1_f (new_AGEMA_signal_9775) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M37_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .A0_f (new_AGEMA_signal_8978), .A1_t (new_AGEMA_signal_8979), .A1_f (new_AGEMA_signal_8980), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29), .B0_f (new_AGEMA_signal_9761), .B1_t (new_AGEMA_signal_9762), .B1_f (new_AGEMA_signal_9763), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .Z0_f (new_AGEMA_signal_10052), .Z1_t (new_AGEMA_signal_10053), .Z1_f (new_AGEMA_signal_10054) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M38_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32), .A0_f (new_AGEMA_signal_9767), .A1_t (new_AGEMA_signal_9768), .A1_f (new_AGEMA_signal_9769), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33), .B0_f (new_AGEMA_signal_9473), .B1_t (new_AGEMA_signal_9474), .B1_f (new_AGEMA_signal_9475), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .Z0_f (new_AGEMA_signal_10055), .Z1_t (new_AGEMA_signal_10056), .Z1_f (new_AGEMA_signal_10057) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M39_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .A0_f (new_AGEMA_signal_9212), .A1_t (new_AGEMA_signal_9213), .A1_f (new_AGEMA_signal_9214), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30), .B0_f (new_AGEMA_signal_9764), .B1_t (new_AGEMA_signal_9765), .B1_f (new_AGEMA_signal_9766), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .Z0_f (new_AGEMA_signal_10058), .Z1_t (new_AGEMA_signal_10059), .Z1_f (new_AGEMA_signal_10060) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M40_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35), .A0_f (new_AGEMA_signal_9770), .A1_t (new_AGEMA_signal_9771), .A1_f (new_AGEMA_signal_9772), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36), .B0_f (new_AGEMA_signal_9773), .B1_t (new_AGEMA_signal_9774), .B1_f (new_AGEMA_signal_9775), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .Z0_f (new_AGEMA_signal_10061), .Z1_t (new_AGEMA_signal_10062), .Z1_f (new_AGEMA_signal_10063) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M41_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .A0_f (new_AGEMA_signal_10055), .A1_t (new_AGEMA_signal_10056), .A1_f (new_AGEMA_signal_10057), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .B0_f (new_AGEMA_signal_10061), .B1_t (new_AGEMA_signal_10062), .B1_f (new_AGEMA_signal_10063), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .Z0_f (new_AGEMA_signal_10364), .Z1_t (new_AGEMA_signal_10365), .Z1_f (new_AGEMA_signal_10366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M42_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .A0_f (new_AGEMA_signal_10052), .A1_t (new_AGEMA_signal_10053), .A1_f (new_AGEMA_signal_10054), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .B0_f (new_AGEMA_signal_10058), .B1_t (new_AGEMA_signal_10059), .B1_f (new_AGEMA_signal_10060), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .Z0_f (new_AGEMA_signal_10367), .Z1_t (new_AGEMA_signal_10368), .Z1_f (new_AGEMA_signal_10369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M43_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .A0_f (new_AGEMA_signal_10052), .A1_t (new_AGEMA_signal_10053), .A1_f (new_AGEMA_signal_10054), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .B0_f (new_AGEMA_signal_10055), .B1_t (new_AGEMA_signal_10056), .B1_f (new_AGEMA_signal_10057), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43), .Z0_f (new_AGEMA_signal_10370), .Z1_t (new_AGEMA_signal_10371), .Z1_f (new_AGEMA_signal_10372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M44_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .A0_f (new_AGEMA_signal_10058), .A1_t (new_AGEMA_signal_10059), .A1_f (new_AGEMA_signal_10060), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .B0_f (new_AGEMA_signal_10061), .B1_t (new_AGEMA_signal_10062), .B1_f (new_AGEMA_signal_10063), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44), .Z0_f (new_AGEMA_signal_10373), .Z1_t (new_AGEMA_signal_10374), .Z1_f (new_AGEMA_signal_10375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M45_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .A0_f (new_AGEMA_signal_10367), .A1_t (new_AGEMA_signal_10368), .A1_f (new_AGEMA_signal_10369), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .B0_f (new_AGEMA_signal_10364), .B1_t (new_AGEMA_signal_10365), .B1_f (new_AGEMA_signal_10366), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45), .Z0_f (new_AGEMA_signal_11084), .Z1_t (new_AGEMA_signal_11085), .Z1_f (new_AGEMA_signal_11086) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M46_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44), .A0_f (new_AGEMA_signal_10373), .A1_t (new_AGEMA_signal_10374), .A1_f (new_AGEMA_signal_10375), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .B0_f (new_AGEMA_signal_6898), .B1_t (new_AGEMA_signal_6899), .B1_f (new_AGEMA_signal_6900), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46), .Z0_f (new_AGEMA_signal_11087), .Z1_t (new_AGEMA_signal_11088), .Z1_f (new_AGEMA_signal_11089) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M47_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .A0_f (new_AGEMA_signal_10061), .A1_t (new_AGEMA_signal_10062), .A1_f (new_AGEMA_signal_10063), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .B0_f (new_AGEMA_signal_7429), .B1_t (new_AGEMA_signal_7430), .B1_f (new_AGEMA_signal_7431), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47), .Z0_f (new_AGEMA_signal_10376), .Z1_t (new_AGEMA_signal_10377), .Z1_f (new_AGEMA_signal_10378) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M48_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .A0_f (new_AGEMA_signal_10058), .A1_t (new_AGEMA_signal_10059), .A1_f (new_AGEMA_signal_10060), .B0_t (RoundKey[24]), .B0_f (new_AGEMA_signal_5459), .B1_t (new_AGEMA_signal_5460), .B1_f (new_AGEMA_signal_5461), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48), .Z0_f (new_AGEMA_signal_10379), .Z1_t (new_AGEMA_signal_10380), .Z1_f (new_AGEMA_signal_10381) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M49_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43), .A0_f (new_AGEMA_signal_10370), .A1_t (new_AGEMA_signal_10371), .A1_f (new_AGEMA_signal_10372), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .B0_f (new_AGEMA_signal_6910), .B1_t (new_AGEMA_signal_6911), .B1_f (new_AGEMA_signal_6912), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49), .Z0_f (new_AGEMA_signal_11090), .Z1_t (new_AGEMA_signal_11091), .Z1_f (new_AGEMA_signal_11092) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M50_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .A0_f (new_AGEMA_signal_10055), .A1_t (new_AGEMA_signal_10056), .A1_f (new_AGEMA_signal_10057), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .B0_f (new_AGEMA_signal_6901), .B1_t (new_AGEMA_signal_6902), .B1_f (new_AGEMA_signal_6903), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50), .Z0_f (new_AGEMA_signal_10382), .Z1_t (new_AGEMA_signal_10383), .Z1_f (new_AGEMA_signal_10384) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M51_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .A0_f (new_AGEMA_signal_10052), .A1_t (new_AGEMA_signal_10053), .A1_f (new_AGEMA_signal_10054), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .B0_f (new_AGEMA_signal_7438), .B1_t (new_AGEMA_signal_7439), .B1_f (new_AGEMA_signal_7440), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51), .Z0_f (new_AGEMA_signal_10385), .Z1_t (new_AGEMA_signal_10386), .Z1_f (new_AGEMA_signal_10387) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M52_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .A0_f (new_AGEMA_signal_10367), .A1_t (new_AGEMA_signal_10368), .A1_f (new_AGEMA_signal_10369), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .B0_f (new_AGEMA_signal_6907), .B1_t (new_AGEMA_signal_6908), .B1_f (new_AGEMA_signal_6909), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52), .Z0_f (new_AGEMA_signal_11093), .Z1_t (new_AGEMA_signal_11094), .Z1_f (new_AGEMA_signal_11095) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M53_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45), .A0_f (new_AGEMA_signal_11084), .A1_t (new_AGEMA_signal_11085), .A1_f (new_AGEMA_signal_11086), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .B0_f (new_AGEMA_signal_6919), .B1_t (new_AGEMA_signal_6920), .B1_f (new_AGEMA_signal_6921), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53), .Z0_f (new_AGEMA_signal_11786), .Z1_t (new_AGEMA_signal_11787), .Z1_f (new_AGEMA_signal_11788) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M54_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .A0_f (new_AGEMA_signal_10364), .A1_t (new_AGEMA_signal_10365), .A1_f (new_AGEMA_signal_10366), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .B0_f (new_AGEMA_signal_7432), .B1_t (new_AGEMA_signal_7433), .B1_f (new_AGEMA_signal_7434), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54), .Z0_f (new_AGEMA_signal_11096), .Z1_t (new_AGEMA_signal_11097), .Z1_f (new_AGEMA_signal_11098) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M55_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44), .A0_f (new_AGEMA_signal_10373), .A1_t (new_AGEMA_signal_10374), .A1_f (new_AGEMA_signal_10375), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .B0_f (new_AGEMA_signal_6904), .B1_t (new_AGEMA_signal_6905), .B1_f (new_AGEMA_signal_6906), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55), .Z0_f (new_AGEMA_signal_11099), .Z1_t (new_AGEMA_signal_11100), .Z1_f (new_AGEMA_signal_11101) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M56_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .A0_f (new_AGEMA_signal_10061), .A1_t (new_AGEMA_signal_10062), .A1_f (new_AGEMA_signal_10063), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .B0_f (new_AGEMA_signal_7444), .B1_t (new_AGEMA_signal_7445), .B1_f (new_AGEMA_signal_7446), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56), .Z0_f (new_AGEMA_signal_10388), .Z1_t (new_AGEMA_signal_10389), .Z1_f (new_AGEMA_signal_10390) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M57_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .A0_f (new_AGEMA_signal_10058), .A1_t (new_AGEMA_signal_10059), .A1_f (new_AGEMA_signal_10060), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .B0_f (new_AGEMA_signal_6913), .B1_t (new_AGEMA_signal_6914), .B1_f (new_AGEMA_signal_6915), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57), .Z0_f (new_AGEMA_signal_10391), .Z1_t (new_AGEMA_signal_10392), .Z1_f (new_AGEMA_signal_10393) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M58_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43), .A0_f (new_AGEMA_signal_10370), .A1_t (new_AGEMA_signal_10371), .A1_f (new_AGEMA_signal_10372), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .B0_f (new_AGEMA_signal_6309), .B1_t (new_AGEMA_signal_6310), .B1_f (new_AGEMA_signal_6311), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58), .Z0_f (new_AGEMA_signal_11102), .Z1_t (new_AGEMA_signal_11103), .Z1_f (new_AGEMA_signal_11104) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M59_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .A0_f (new_AGEMA_signal_10055), .A1_t (new_AGEMA_signal_10056), .A1_f (new_AGEMA_signal_10057), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .B0_f (new_AGEMA_signal_6916), .B1_t (new_AGEMA_signal_6917), .B1_f (new_AGEMA_signal_6918), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59), .Z0_f (new_AGEMA_signal_10394), .Z1_t (new_AGEMA_signal_10395), .Z1_f (new_AGEMA_signal_10396) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M60_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .A0_f (new_AGEMA_signal_10052), .A1_t (new_AGEMA_signal_10053), .A1_f (new_AGEMA_signal_10054), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .B0_f (new_AGEMA_signal_7441), .B1_t (new_AGEMA_signal_7442), .B1_f (new_AGEMA_signal_7443), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60), .Z0_f (new_AGEMA_signal_10397), .Z1_t (new_AGEMA_signal_10398), .Z1_f (new_AGEMA_signal_10399) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M61_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .A0_f (new_AGEMA_signal_10367), .A1_t (new_AGEMA_signal_10368), .A1_f (new_AGEMA_signal_10369), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .B0_f (new_AGEMA_signal_6303), .B1_t (new_AGEMA_signal_6304), .B1_f (new_AGEMA_signal_6305), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .Z0_f (new_AGEMA_signal_11105), .Z1_t (new_AGEMA_signal_11106), .Z1_f (new_AGEMA_signal_11107) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M62_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45), .A0_f (new_AGEMA_signal_11084), .A1_t (new_AGEMA_signal_11085), .A1_f (new_AGEMA_signal_11086), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .B0_f (new_AGEMA_signal_6312), .B1_t (new_AGEMA_signal_6313), .B1_f (new_AGEMA_signal_6314), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62), .Z0_f (new_AGEMA_signal_11789), .Z1_t (new_AGEMA_signal_11790), .Z1_f (new_AGEMA_signal_11791) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M63_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .A0_f (new_AGEMA_signal_10364), .A1_t (new_AGEMA_signal_10365), .A1_f (new_AGEMA_signal_10366), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .B0_f (new_AGEMA_signal_6306), .B1_t (new_AGEMA_signal_6307), .B1_f (new_AGEMA_signal_6308), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63), .Z0_f (new_AGEMA_signal_11108), .Z1_t (new_AGEMA_signal_11109), .Z1_f (new_AGEMA_signal_11110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .A0_f (new_AGEMA_signal_11105), .A1_t (new_AGEMA_signal_11106), .A1_f (new_AGEMA_signal_11107), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62), .B0_f (new_AGEMA_signal_11789), .B1_t (new_AGEMA_signal_11790), .B1_f (new_AGEMA_signal_11791), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .Z0_f (new_AGEMA_signal_12377), .Z1_t (new_AGEMA_signal_12378), .Z1_f (new_AGEMA_signal_12379) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50), .A0_f (new_AGEMA_signal_10382), .A1_t (new_AGEMA_signal_10383), .A1_f (new_AGEMA_signal_10384), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56), .B0_f (new_AGEMA_signal_10388), .B1_t (new_AGEMA_signal_10389), .B1_f (new_AGEMA_signal_10390), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .Z0_f (new_AGEMA_signal_11111), .Z1_t (new_AGEMA_signal_11112), .Z1_f (new_AGEMA_signal_11113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46), .A0_f (new_AGEMA_signal_11087), .A1_t (new_AGEMA_signal_11088), .A1_f (new_AGEMA_signal_11089), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48), .B0_f (new_AGEMA_signal_10379), .B1_t (new_AGEMA_signal_10380), .B1_f (new_AGEMA_signal_10381), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2), .Z0_f (new_AGEMA_signal_11792), .Z1_t (new_AGEMA_signal_11793), .Z1_f (new_AGEMA_signal_11794) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47), .A0_f (new_AGEMA_signal_10376), .A1_t (new_AGEMA_signal_10377), .A1_f (new_AGEMA_signal_10378), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55), .B0_f (new_AGEMA_signal_11099), .B1_t (new_AGEMA_signal_11100), .B1_f (new_AGEMA_signal_11101), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3), .Z0_f (new_AGEMA_signal_11795), .Z1_t (new_AGEMA_signal_11796), .Z1_f (new_AGEMA_signal_11797) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54), .A0_f (new_AGEMA_signal_11096), .A1_t (new_AGEMA_signal_11097), .A1_f (new_AGEMA_signal_11098), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58), .B0_f (new_AGEMA_signal_11102), .B1_t (new_AGEMA_signal_11103), .B1_f (new_AGEMA_signal_11104), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4), .Z0_f (new_AGEMA_signal_11798), .Z1_t (new_AGEMA_signal_11799), .Z1_f (new_AGEMA_signal_11800) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49), .A0_f (new_AGEMA_signal_11090), .A1_t (new_AGEMA_signal_11091), .A1_f (new_AGEMA_signal_11092), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .B0_f (new_AGEMA_signal_11105), .B1_t (new_AGEMA_signal_11106), .B1_f (new_AGEMA_signal_11107), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5), .Z0_f (new_AGEMA_signal_11801), .Z1_t (new_AGEMA_signal_11802), .Z1_f (new_AGEMA_signal_11803) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62), .A0_f (new_AGEMA_signal_11789), .A1_t (new_AGEMA_signal_11790), .A1_f (new_AGEMA_signal_11791), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5), .B0_f (new_AGEMA_signal_11801), .B1_t (new_AGEMA_signal_11802), .B1_f (new_AGEMA_signal_11803), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .Z0_f (new_AGEMA_signal_12380), .Z1_t (new_AGEMA_signal_12381), .Z1_f (new_AGEMA_signal_12382) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46), .A0_f (new_AGEMA_signal_11087), .A1_t (new_AGEMA_signal_11088), .A1_f (new_AGEMA_signal_11089), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3), .B0_f (new_AGEMA_signal_11795), .B1_t (new_AGEMA_signal_11796), .B1_f (new_AGEMA_signal_11797), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7), .Z0_f (new_AGEMA_signal_12383), .Z1_t (new_AGEMA_signal_12384), .Z1_f (new_AGEMA_signal_12385) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51), .A0_f (new_AGEMA_signal_10385), .A1_t (new_AGEMA_signal_10386), .A1_f (new_AGEMA_signal_10387), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59), .B0_f (new_AGEMA_signal_10394), .B1_t (new_AGEMA_signal_10395), .B1_f (new_AGEMA_signal_10396), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8), .Z0_f (new_AGEMA_signal_11114), .Z1_t (new_AGEMA_signal_11115), .Z1_f (new_AGEMA_signal_11116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52), .A0_f (new_AGEMA_signal_11093), .A1_t (new_AGEMA_signal_11094), .A1_f (new_AGEMA_signal_11095), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53), .B0_f (new_AGEMA_signal_11786), .B1_t (new_AGEMA_signal_11787), .B1_f (new_AGEMA_signal_11788), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9), .Z0_f (new_AGEMA_signal_12386), .Z1_t (new_AGEMA_signal_12387), .Z1_f (new_AGEMA_signal_12388) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53), .A0_f (new_AGEMA_signal_11786), .A1_t (new_AGEMA_signal_11787), .A1_f (new_AGEMA_signal_11788), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4), .B0_f (new_AGEMA_signal_11798), .B1_t (new_AGEMA_signal_11799), .B1_f (new_AGEMA_signal_11800), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10), .Z0_f (new_AGEMA_signal_12389), .Z1_t (new_AGEMA_signal_12390), .Z1_f (new_AGEMA_signal_12391) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60), .A0_f (new_AGEMA_signal_10397), .A1_t (new_AGEMA_signal_10398), .A1_f (new_AGEMA_signal_10399), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2), .B0_f (new_AGEMA_signal_11792), .B1_t (new_AGEMA_signal_11793), .B1_f (new_AGEMA_signal_11794), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11), .Z0_f (new_AGEMA_signal_12392), .Z1_t (new_AGEMA_signal_12393), .Z1_f (new_AGEMA_signal_12394) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48), .A0_f (new_AGEMA_signal_10379), .A1_t (new_AGEMA_signal_10380), .A1_f (new_AGEMA_signal_10381), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51), .B0_f (new_AGEMA_signal_10385), .B1_t (new_AGEMA_signal_10386), .B1_f (new_AGEMA_signal_10387), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12), .Z0_f (new_AGEMA_signal_11117), .Z1_t (new_AGEMA_signal_11118), .Z1_f (new_AGEMA_signal_11119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50), .A0_f (new_AGEMA_signal_10382), .A1_t (new_AGEMA_signal_10383), .A1_f (new_AGEMA_signal_10384), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .B0_f (new_AGEMA_signal_12377), .B1_t (new_AGEMA_signal_12378), .B1_f (new_AGEMA_signal_12379), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13), .Z0_f (new_AGEMA_signal_12935), .Z1_t (new_AGEMA_signal_12936), .Z1_f (new_AGEMA_signal_12937) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52), .A0_f (new_AGEMA_signal_11093), .A1_t (new_AGEMA_signal_11094), .A1_f (new_AGEMA_signal_11095), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .B0_f (new_AGEMA_signal_11105), .B1_t (new_AGEMA_signal_11106), .B1_f (new_AGEMA_signal_11107), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14), .Z0_f (new_AGEMA_signal_11804), .Z1_t (new_AGEMA_signal_11805), .Z1_f (new_AGEMA_signal_11806) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55), .A0_f (new_AGEMA_signal_11099), .A1_t (new_AGEMA_signal_11100), .A1_f (new_AGEMA_signal_11101), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .B0_f (new_AGEMA_signal_11111), .B1_t (new_AGEMA_signal_11112), .B1_f (new_AGEMA_signal_11113), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15), .Z0_f (new_AGEMA_signal_11807), .Z1_t (new_AGEMA_signal_11808), .Z1_f (new_AGEMA_signal_11809) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56), .A0_f (new_AGEMA_signal_10388), .A1_t (new_AGEMA_signal_10389), .A1_f (new_AGEMA_signal_10390), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .B0_f (new_AGEMA_signal_12377), .B1_t (new_AGEMA_signal_12378), .B1_f (new_AGEMA_signal_12379), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16), .Z0_f (new_AGEMA_signal_12938), .Z1_t (new_AGEMA_signal_12939), .Z1_f (new_AGEMA_signal_12940) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57), .A0_f (new_AGEMA_signal_10391), .A1_t (new_AGEMA_signal_10392), .A1_f (new_AGEMA_signal_10393), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .B0_f (new_AGEMA_signal_11111), .B1_t (new_AGEMA_signal_11112), .B1_f (new_AGEMA_signal_11113), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17), .Z0_f (new_AGEMA_signal_11810), .Z1_t (new_AGEMA_signal_11811), .Z1_f (new_AGEMA_signal_11812) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58), .A0_f (new_AGEMA_signal_11102), .A1_t (new_AGEMA_signal_11103), .A1_f (new_AGEMA_signal_11104), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8), .B0_f (new_AGEMA_signal_11114), .B1_t (new_AGEMA_signal_11115), .B1_f (new_AGEMA_signal_11116), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18), .Z0_f (new_AGEMA_signal_11813), .Z1_t (new_AGEMA_signal_11814), .Z1_f (new_AGEMA_signal_11815) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63), .A0_f (new_AGEMA_signal_11108), .A1_t (new_AGEMA_signal_11109), .A1_f (new_AGEMA_signal_11110), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4), .B0_f (new_AGEMA_signal_11798), .B1_t (new_AGEMA_signal_11799), .B1_f (new_AGEMA_signal_11800), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19), .Z0_f (new_AGEMA_signal_12395), .Z1_t (new_AGEMA_signal_12396), .Z1_f (new_AGEMA_signal_12397) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .A0_f (new_AGEMA_signal_12377), .A1_t (new_AGEMA_signal_12378), .A1_f (new_AGEMA_signal_12379), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .B0_f (new_AGEMA_signal_11111), .B1_t (new_AGEMA_signal_11112), .B1_f (new_AGEMA_signal_11113), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20), .Z0_f (new_AGEMA_signal_12941), .Z1_t (new_AGEMA_signal_12942), .Z1_f (new_AGEMA_signal_12943) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .A0_f (new_AGEMA_signal_11111), .A1_t (new_AGEMA_signal_11112), .A1_f (new_AGEMA_signal_11113), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7), .B0_f (new_AGEMA_signal_12383), .B1_t (new_AGEMA_signal_12384), .B1_f (new_AGEMA_signal_12385), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21), .Z0_f (new_AGEMA_signal_12944), .Z1_t (new_AGEMA_signal_12945), .Z1_f (new_AGEMA_signal_12946) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3), .A0_f (new_AGEMA_signal_11795), .A1_t (new_AGEMA_signal_11796), .A1_f (new_AGEMA_signal_11797), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12), .B0_f (new_AGEMA_signal_11117), .B1_t (new_AGEMA_signal_11118), .B1_f (new_AGEMA_signal_11119), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22), .Z0_f (new_AGEMA_signal_12398), .Z1_t (new_AGEMA_signal_12399), .Z1_f (new_AGEMA_signal_12400) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18), .A0_f (new_AGEMA_signal_11813), .A1_t (new_AGEMA_signal_11814), .A1_f (new_AGEMA_signal_11815), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2), .B0_f (new_AGEMA_signal_11792), .B1_t (new_AGEMA_signal_11793), .B1_f (new_AGEMA_signal_11794), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23), .Z0_f (new_AGEMA_signal_12401), .Z1_t (new_AGEMA_signal_12402), .Z1_f (new_AGEMA_signal_12403) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15), .A0_f (new_AGEMA_signal_11807), .A1_t (new_AGEMA_signal_11808), .A1_f (new_AGEMA_signal_11809), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9), .B0_f (new_AGEMA_signal_12386), .B1_t (new_AGEMA_signal_12387), .B1_f (new_AGEMA_signal_12388), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24), .Z0_f (new_AGEMA_signal_12947), .Z1_t (new_AGEMA_signal_12948), .Z1_f (new_AGEMA_signal_12949) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .A0_f (new_AGEMA_signal_12380), .A1_t (new_AGEMA_signal_12381), .A1_f (new_AGEMA_signal_12382), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10), .B0_f (new_AGEMA_signal_12389), .B1_t (new_AGEMA_signal_12390), .B1_f (new_AGEMA_signal_12391), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25), .Z0_f (new_AGEMA_signal_12950), .Z1_t (new_AGEMA_signal_12951), .Z1_f (new_AGEMA_signal_12952) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7), .A0_f (new_AGEMA_signal_12383), .A1_t (new_AGEMA_signal_12384), .A1_f (new_AGEMA_signal_12385), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9), .B0_f (new_AGEMA_signal_12386), .B1_t (new_AGEMA_signal_12387), .B1_f (new_AGEMA_signal_12388), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26), .Z0_f (new_AGEMA_signal_12953), .Z1_t (new_AGEMA_signal_12954), .Z1_f (new_AGEMA_signal_12955) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8), .A0_f (new_AGEMA_signal_11114), .A1_t (new_AGEMA_signal_11115), .A1_f (new_AGEMA_signal_11116), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10), .B0_f (new_AGEMA_signal_12389), .B1_t (new_AGEMA_signal_12390), .B1_f (new_AGEMA_signal_12391), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27), .Z0_f (new_AGEMA_signal_12956), .Z1_t (new_AGEMA_signal_12957), .Z1_f (new_AGEMA_signal_12958) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11), .A0_f (new_AGEMA_signal_12392), .A1_t (new_AGEMA_signal_12393), .A1_f (new_AGEMA_signal_12394), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14), .B0_f (new_AGEMA_signal_11804), .B1_t (new_AGEMA_signal_11805), .B1_f (new_AGEMA_signal_11806), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28), .Z0_f (new_AGEMA_signal_12959), .Z1_t (new_AGEMA_signal_12960), .Z1_f (new_AGEMA_signal_12961) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11), .A0_f (new_AGEMA_signal_12392), .A1_t (new_AGEMA_signal_12393), .A1_f (new_AGEMA_signal_12394), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17), .B0_f (new_AGEMA_signal_11810), .B1_t (new_AGEMA_signal_11811), .B1_f (new_AGEMA_signal_11812), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29), .Z0_f (new_AGEMA_signal_12962), .Z1_t (new_AGEMA_signal_12963), .Z1_f (new_AGEMA_signal_12964) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .A0_f (new_AGEMA_signal_12380), .A1_t (new_AGEMA_signal_12381), .A1_f (new_AGEMA_signal_12382), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24), .B0_f (new_AGEMA_signal_12947), .B1_t (new_AGEMA_signal_12948), .B1_f (new_AGEMA_signal_12949), .Z0_t (KeyExpansionIns_tmp[7]), .Z0_f (new_AGEMA_signal_13571), .Z1_t (new_AGEMA_signal_13572), .Z1_f (new_AGEMA_signal_13573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16), .A0_f (new_AGEMA_signal_12938), .A1_t (new_AGEMA_signal_12939), .A1_f (new_AGEMA_signal_12940), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26), .B0_f (new_AGEMA_signal_12953), .B1_t (new_AGEMA_signal_12954), .B1_f (new_AGEMA_signal_12955), .Z0_t (KeyExpansionIns_tmp[6]), .Z0_f (new_AGEMA_signal_13574), .Z1_t (new_AGEMA_signal_13575), .Z1_f (new_AGEMA_signal_13576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19), .A0_f (new_AGEMA_signal_12395), .A1_t (new_AGEMA_signal_12396), .A1_f (new_AGEMA_signal_12397), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28), .B0_f (new_AGEMA_signal_12959), .B1_t (new_AGEMA_signal_12960), .B1_f (new_AGEMA_signal_12961), .Z0_t (KeyExpansionIns_tmp[5]), .Z0_f (new_AGEMA_signal_13577), .Z1_t (new_AGEMA_signal_13578), .Z1_f (new_AGEMA_signal_13579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .A0_f (new_AGEMA_signal_12380), .A1_t (new_AGEMA_signal_12381), .A1_f (new_AGEMA_signal_12382), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21), .B0_f (new_AGEMA_signal_12944), .B1_t (new_AGEMA_signal_12945), .B1_f (new_AGEMA_signal_12946), .Z0_t (KeyExpansionIns_tmp[4]), .Z0_f (new_AGEMA_signal_13580), .Z1_t (new_AGEMA_signal_13581), .Z1_f (new_AGEMA_signal_13582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20), .A0_f (new_AGEMA_signal_12941), .A1_t (new_AGEMA_signal_12942), .A1_f (new_AGEMA_signal_12943), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22), .B0_f (new_AGEMA_signal_12398), .B1_t (new_AGEMA_signal_12399), .B1_f (new_AGEMA_signal_12400), .Z0_t (KeyExpansionIns_tmp[3]), .Z0_f (new_AGEMA_signal_13583), .Z1_t (new_AGEMA_signal_13584), .Z1_f (new_AGEMA_signal_13585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25), .A0_f (new_AGEMA_signal_12950), .A1_t (new_AGEMA_signal_12951), .A1_f (new_AGEMA_signal_12952), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29), .B0_f (new_AGEMA_signal_12962), .B1_t (new_AGEMA_signal_12963), .B1_f (new_AGEMA_signal_12964), .Z0_t (KeyExpansionIns_tmp[2]), .Z0_f (new_AGEMA_signal_13586), .Z1_t (new_AGEMA_signal_13587), .Z1_f (new_AGEMA_signal_13588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13), .A0_f (new_AGEMA_signal_12935), .A1_t (new_AGEMA_signal_12936), .A1_f (new_AGEMA_signal_12937), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27), .B0_f (new_AGEMA_signal_12956), .B1_t (new_AGEMA_signal_12957), .B1_f (new_AGEMA_signal_12958), .Z0_t (KeyExpansionIns_tmp[1]), .Z0_f (new_AGEMA_signal_13589), .Z1_t (new_AGEMA_signal_13590), .Z1_f (new_AGEMA_signal_13591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .A0_f (new_AGEMA_signal_12380), .A1_t (new_AGEMA_signal_12381), .A1_f (new_AGEMA_signal_12382), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23), .B0_f (new_AGEMA_signal_12401), .B1_t (new_AGEMA_signal_12402), .B1_f (new_AGEMA_signal_12403), .Z0_t (KeyExpansionIns_tmp[0]), .Z0_f (new_AGEMA_signal_12965), .Z1_t (new_AGEMA_signal_12966), .Z1_f (new_AGEMA_signal_12967) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) RoundCounterIns_U11 ( .A0_t (start_t), .A0_f (start_f), .B0_t (RoundCounterIns_n5), .B0_f (new_AGEMA_signal_6922), .Z0_t (RoundCounter[2]), .Z0_f (new_AGEMA_signal_5052) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) RoundCounterIns_U10 ( .A0_t (RoundCounter[2]), .A0_f (new_AGEMA_signal_5052), .B0_t (RoundCounterIns_n4), .B0_f (new_AGEMA_signal_6334), .Z0_t (RoundCounterIns_n5), .Z0_f (new_AGEMA_signal_6922) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) RoundCounterIns_U9 ( .A0_t (start_t), .A0_f (start_f), .B0_t (RoundCounterIns_n3), .B0_f (new_AGEMA_signal_6333), .Z0_t (RoundCounter[1]), .Z0_f (new_AGEMA_signal_5051) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) RoundCounterIns_U8 ( .A0_t (RoundCounter[1]), .A0_f (new_AGEMA_signal_5051), .B0_t (RoundCounter[0]), .B0_f (new_AGEMA_signal_5054), .Z0_t (RoundCounterIns_n3), .Z0_f (new_AGEMA_signal_6333) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) RoundCounterIns_U7 ( .A0_t (start_t), .A0_f (start_f), .B0_t (RoundCounterIns_n2), .B0_f (new_AGEMA_signal_7468), .Z0_t (RoundCounter[3]), .Z0_f (new_AGEMA_signal_5055) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) RoundCounterIns_U6 ( .A0_t (RoundCounter[3]), .A0_f (new_AGEMA_signal_5055), .B0_t (RoundCounterIns_n1), .B0_f (new_AGEMA_signal_6923), .Z0_t (RoundCounterIns_n2), .Z0_f (new_AGEMA_signal_7468) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) RoundCounterIns_U5 ( .A0_t (RoundCounterIns_n4), .A0_f (new_AGEMA_signal_6334), .B0_t (RoundCounter[2]), .B0_f (new_AGEMA_signal_5052), .Z0_t (RoundCounterIns_n1), .Z0_f (new_AGEMA_signal_6923) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) RoundCounterIns_U4 ( .A0_t (RoundCounter[0]), .A0_f (new_AGEMA_signal_5054), .B0_t (RoundCounter[1]), .B0_f (new_AGEMA_signal_5051), .Z0_t (RoundCounterIns_n4), .Z0_f (new_AGEMA_signal_6334) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) RoundCounterIns_U3 ( .A0_t (start_t), .A0_f (start_f), .B0_t (RoundCounter[0]), .B0_f (new_AGEMA_signal_5054), .Z0_t (RoundCounter[0]), .Z0_f (new_AGEMA_signal_5054) ) ;

    /* register cells */
endmodule
