module eFPGA_top
    #(
        parameter include_eFPGA=1,
        parameter NumberOfRows=23,
        parameter NumberOfCols=11,
        parameter FrameBitsPerRow=32,
        parameter MaxFramesPerCol=20,
        parameter desync_flag=20,
        parameter FrameSelectWidth=7,
        parameter RowSelectWidth=7
    )
    (
        //External IO port
        output [92-1:0] A_config_C,
        output [92-1:0] B_config_C,
        output [23-1:0] I_top_0_t,
        output [23-1:0] I_top_0_f,
        output [23-1:0] I_top_1_t,
        output [23-1:0] I_top_1_f,
        output [23-1:0] T_top,
        input [23-1:0] O_top_0_t,
        input [23-1:0] O_top_0_f,
        input [23-1:0] O_top_1_t,
        input [23-1:0] O_top_1_f,
        output [23-1:0] ctrl_I_top_0_t,
        output [23-1:0] ctrl_I_top_0_f,
        output [23-1:0] ctrl_T_top,
        input [23-1:0] ctrl_O_top_0_t,
        input [23-1:0] ctrl_O_top_0_f,

        //Custom ports (*SAUBER*)
        input rst,
        output f_detected,
        output prech1,
        output prech2,
        input prng_rst,
        input [79:0] key_t,
        input [79:0] key_f,
        input [79:0] iv_t,
        input [79:0] iv_f,

        //Config related ports
        input CLK,
        input resetn,
        input SelfWriteStrobe,
        input [31:0] SelfWriteData,
        input Rx,
        output ComActive,
        output ReceiveLED,
        input s_clk,
        input s_data
);

 //Custom signal declarations for SAUBER
wire[22:0] F_masked1_top;
wire[22:0] F_masked2_top;
wire[22:0] F_ctrl_top;
wire[574:0] R_t_top;
wire[574:0] R_f_top;


 //Signal declarations
wire[(NumberOfRows*FrameBitsPerRow)-1:0] FrameRegister;
wire[(MaxFramesPerCol*NumberOfCols)-1:0] FrameSelect;
wire[(FrameBitsPerRow*(NumberOfRows+2))-1:0] FrameData;
wire[FrameBitsPerRow-1:0] FrameAddressRegister;
wire LongFrameStrobe;
wire[31:0] LocalWriteData;
wire LocalWriteStrobe;
wire[RowSelectWidth-1:0] RowSelect;
wire resten;
`ifndef EMULATION

eFPGA_Config
    #(
    .RowSelectWidth(RowSelectWidth),
    .NumberOfRows(NumberOfRows),
    .desync_flag(desync_flag),
    .FrameBitsPerRow(FrameBitsPerRow)
    )
    eFPGA_Config_inst
    (
    .CLK(CLK),
    .resetn(resetn),
    .Rx(Rx),
    .ComActive(ComActive),
    .ReceiveLED(ReceiveLED),
    .s_clk(s_clk),
    .s_data(s_data),
    .SelfWriteData(SelfWriteData),
    .SelfWriteStrobe(SelfWriteStrobe),
    .ConfigWriteData(LocalWriteData),
    .ConfigWriteStrobe(LocalWriteStrobe),
    .FrameAddressRegister(FrameAddressRegister),
    .LongFrameStrobe(LongFrameStrobe),
    .RowSelect(RowSelect)
);


Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(1)
    )
    inst_Frame_Data_Reg_0
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[0*FrameBitsPerRow+FrameBitsPerRow-1:0*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(2)
    )
    inst_Frame_Data_Reg_1
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[1*FrameBitsPerRow+FrameBitsPerRow-1:1*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(3)
    )
    inst_Frame_Data_Reg_2
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[2*FrameBitsPerRow+FrameBitsPerRow-1:2*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(4)
    )
    inst_Frame_Data_Reg_3
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[3*FrameBitsPerRow+FrameBitsPerRow-1:3*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(5)
    )
    inst_Frame_Data_Reg_4
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[4*FrameBitsPerRow+FrameBitsPerRow-1:4*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(6)
    )
    inst_Frame_Data_Reg_5
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[5*FrameBitsPerRow+FrameBitsPerRow-1:5*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(7)
    )
    inst_Frame_Data_Reg_6
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[6*FrameBitsPerRow+FrameBitsPerRow-1:6*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(8)
    )
    inst_Frame_Data_Reg_7
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[7*FrameBitsPerRow+FrameBitsPerRow-1:7*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(9)
    )
    inst_Frame_Data_Reg_8
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[8*FrameBitsPerRow+FrameBitsPerRow-1:8*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(10)
    )
    inst_Frame_Data_Reg_9
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[9*FrameBitsPerRow+FrameBitsPerRow-1:9*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(11)
    )
    inst_Frame_Data_Reg_10
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[10*FrameBitsPerRow+FrameBitsPerRow-1:10*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(12)
    )
    inst_Frame_Data_Reg_11
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[11*FrameBitsPerRow+FrameBitsPerRow-1:11*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(13)
    )
    inst_Frame_Data_Reg_12
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[12*FrameBitsPerRow+FrameBitsPerRow-1:12*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(14)
    )
    inst_Frame_Data_Reg_13
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[13*FrameBitsPerRow+FrameBitsPerRow-1:13*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(15)
    )
    inst_Frame_Data_Reg_14
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[14*FrameBitsPerRow+FrameBitsPerRow-1:14*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(16)
    )
    inst_Frame_Data_Reg_15
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[15*FrameBitsPerRow+FrameBitsPerRow-1:15*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(17)
    )
    inst_Frame_Data_Reg_16
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[16*FrameBitsPerRow+FrameBitsPerRow-1:16*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(18)
    )
    inst_Frame_Data_Reg_17
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[17*FrameBitsPerRow+FrameBitsPerRow-1:17*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(19)
    )
    inst_Frame_Data_Reg_18
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[18*FrameBitsPerRow+FrameBitsPerRow-1:18*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(20)
    )
    inst_Frame_Data_Reg_19
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[19*FrameBitsPerRow+FrameBitsPerRow-1:19*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(21)
    )
    inst_Frame_Data_Reg_20
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[20*FrameBitsPerRow+FrameBitsPerRow-1:20*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(22)
    )
    inst_Frame_Data_Reg_21
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[21*FrameBitsPerRow+FrameBitsPerRow-1:21*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(23)
    )
    inst_Frame_Data_Reg_22
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[22*FrameBitsPerRow+FrameBitsPerRow-1:22*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);


Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(0)
    )
    inst_Frame_Select_0
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[0*MaxFramesPerCol+MaxFramesPerCol-1:0*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(1)
    )
    inst_Frame_Select_1
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[1*MaxFramesPerCol+MaxFramesPerCol-1:1*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(2)
    )
    inst_Frame_Select_2
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[2*MaxFramesPerCol+MaxFramesPerCol-1:2*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(3)
    )
    inst_Frame_Select_3
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[3*MaxFramesPerCol+MaxFramesPerCol-1:3*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(4)
    )
    inst_Frame_Select_4
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[4*MaxFramesPerCol+MaxFramesPerCol-1:4*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(5)
    )
    inst_Frame_Select_5
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[5*MaxFramesPerCol+MaxFramesPerCol-1:5*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(6)
    )
    inst_Frame_Select_6
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[6*MaxFramesPerCol+MaxFramesPerCol-1:6*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(7)
    )
    inst_Frame_Select_7
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[7*MaxFramesPerCol+MaxFramesPerCol-1:7*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(8)
    )
    inst_Frame_Select_8
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[8*MaxFramesPerCol+MaxFramesPerCol-1:8*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(9)
    )
    inst_Frame_Select_9
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[9*MaxFramesPerCol+MaxFramesPerCol-1:9*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(10)
    )
    inst_Frame_Select_10
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[10*MaxFramesPerCol+MaxFramesPerCol-1:10*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);


`endif
eFPGA eFPGA_inst (
    .Tile_X3Y1_R_t(R_t_top[0]),
    .Tile_X3Y1_R_f(R_f_top[0]),
    .Tile_X6Y1_R_t(R_t_top[1]),
    .Tile_X6Y1_R_f(R_f_top[1]),
    .Tile_X9Y1_R_t(R_t_top[2]),
    .Tile_X9Y1_R_f(R_f_top[2]),
    .Tile_X12Y1_R_t(R_t_top[3]),
    .Tile_X12Y1_R_f(R_f_top[3]),
    .Tile_X15Y1_R_t(R_t_top[4]),
    .Tile_X15Y1_R_f(R_f_top[4]),
    .Tile_X18Y1_R_t(R_t_top[5]),
    .Tile_X18Y1_R_f(R_f_top[5]),
    .Tile_X21Y1_R_t(R_t_top[6]),
    .Tile_X21Y1_R_f(R_f_top[6]),
    .Tile_X24Y1_R_t(R_t_top[7]),
    .Tile_X24Y1_R_f(R_f_top[7]),
    .Tile_X27Y1_R_t(R_t_top[8]),
    .Tile_X27Y1_R_f(R_f_top[8]),
    .Tile_X30Y1_R_t(R_t_top[9]),
    .Tile_X30Y1_R_f(R_f_top[9]),
    .Tile_X33Y1_R_t(R_t_top[10]),
    .Tile_X33Y1_R_f(R_f_top[10]),
    .Tile_X36Y1_R_t(R_t_top[11]),
    .Tile_X36Y1_R_f(R_f_top[11]),
    .Tile_X39Y1_R_t(R_t_top[12]),
    .Tile_X39Y1_R_f(R_f_top[12]),
    .Tile_X42Y1_R_t(R_t_top[13]),
    .Tile_X42Y1_R_f(R_f_top[13]),
    .Tile_X45Y1_R_t(R_t_top[14]),
    .Tile_X45Y1_R_f(R_f_top[14]),
    .Tile_X48Y1_R_t(R_t_top[15]),
    .Tile_X48Y1_R_f(R_f_top[15]),
    .Tile_X51Y1_R_t(R_t_top[16]),
    .Tile_X51Y1_R_f(R_f_top[16]),
    .Tile_X54Y1_R_t(R_t_top[17]),
    .Tile_X54Y1_R_f(R_f_top[17]),
    .Tile_X57Y1_R_t(R_t_top[18]),
    .Tile_X57Y1_R_f(R_f_top[18]),
    .Tile_X60Y1_R_t(R_t_top[19]),
    .Tile_X60Y1_R_f(R_f_top[19]),
    .Tile_X63Y1_R_t(R_t_top[20]),
    .Tile_X63Y1_R_f(R_f_top[20]),
    .Tile_X66Y1_R_t(R_t_top[21]),
    .Tile_X66Y1_R_f(R_f_top[21]),
    .Tile_X69Y1_R_t(R_t_top[22]),
    .Tile_X69Y1_R_f(R_f_top[22]),
    .Tile_X72Y1_R_t(R_t_top[23]),
    .Tile_X72Y1_R_f(R_f_top[23]),
    .Tile_X75Y1_R_t(R_t_top[24]),
    .Tile_X75Y1_R_f(R_f_top[24]),
    .Tile_X3Y2_R_t(R_t_top[25]),
    .Tile_X3Y2_R_f(R_f_top[25]),
    .Tile_X6Y2_R_t(R_t_top[26]),
    .Tile_X6Y2_R_f(R_f_top[26]),
    .Tile_X9Y2_R_t(R_t_top[27]),
    .Tile_X9Y2_R_f(R_f_top[27]),
    .Tile_X12Y2_R_t(R_t_top[28]),
    .Tile_X12Y2_R_f(R_f_top[28]),
    .Tile_X15Y2_R_t(R_t_top[29]),
    .Tile_X15Y2_R_f(R_f_top[29]),
    .Tile_X18Y2_R_t(R_t_top[30]),
    .Tile_X18Y2_R_f(R_f_top[30]),
    .Tile_X21Y2_R_t(R_t_top[31]),
    .Tile_X21Y2_R_f(R_f_top[31]),
    .Tile_X24Y2_R_t(R_t_top[32]),
    .Tile_X24Y2_R_f(R_f_top[32]),
    .Tile_X27Y2_R_t(R_t_top[33]),
    .Tile_X27Y2_R_f(R_f_top[33]),
    .Tile_X30Y2_R_t(R_t_top[34]),
    .Tile_X30Y2_R_f(R_f_top[34]),
    .Tile_X33Y2_R_t(R_t_top[35]),
    .Tile_X33Y2_R_f(R_f_top[35]),
    .Tile_X36Y2_R_t(R_t_top[36]),
    .Tile_X36Y2_R_f(R_f_top[36]),
    .Tile_X39Y2_R_t(R_t_top[37]),
    .Tile_X39Y2_R_f(R_f_top[37]),
    .Tile_X42Y2_R_t(R_t_top[38]),
    .Tile_X42Y2_R_f(R_f_top[38]),
    .Tile_X45Y2_R_t(R_t_top[39]),
    .Tile_X45Y2_R_f(R_f_top[39]),
    .Tile_X48Y2_R_t(R_t_top[40]),
    .Tile_X48Y2_R_f(R_f_top[40]),
    .Tile_X51Y2_R_t(R_t_top[41]),
    .Tile_X51Y2_R_f(R_f_top[41]),
    .Tile_X54Y2_R_t(R_t_top[42]),
    .Tile_X54Y2_R_f(R_f_top[42]),
    .Tile_X57Y2_R_t(R_t_top[43]),
    .Tile_X57Y2_R_f(R_f_top[43]),
    .Tile_X60Y2_R_t(R_t_top[44]),
    .Tile_X60Y2_R_f(R_f_top[44]),
    .Tile_X63Y2_R_t(R_t_top[45]),
    .Tile_X63Y2_R_f(R_f_top[45]),
    .Tile_X66Y2_R_t(R_t_top[46]),
    .Tile_X66Y2_R_f(R_f_top[46]),
    .Tile_X69Y2_R_t(R_t_top[47]),
    .Tile_X69Y2_R_f(R_f_top[47]),
    .Tile_X72Y2_R_t(R_t_top[48]),
    .Tile_X72Y2_R_f(R_f_top[48]),
    .Tile_X75Y2_R_t(R_t_top[49]),
    .Tile_X75Y2_R_f(R_f_top[49]),
    .Tile_X3Y3_R_t(R_t_top[50]),
    .Tile_X3Y3_R_f(R_f_top[50]),
    .Tile_X6Y3_R_t(R_t_top[51]),
    .Tile_X6Y3_R_f(R_f_top[51]),
    .Tile_X9Y3_R_t(R_t_top[52]),
    .Tile_X9Y3_R_f(R_f_top[52]),
    .Tile_X12Y3_R_t(R_t_top[53]),
    .Tile_X12Y3_R_f(R_f_top[53]),
    .Tile_X15Y3_R_t(R_t_top[54]),
    .Tile_X15Y3_R_f(R_f_top[54]),
    .Tile_X18Y3_R_t(R_t_top[55]),
    .Tile_X18Y3_R_f(R_f_top[55]),
    .Tile_X21Y3_R_t(R_t_top[56]),
    .Tile_X21Y3_R_f(R_f_top[56]),
    .Tile_X24Y3_R_t(R_t_top[57]),
    .Tile_X24Y3_R_f(R_f_top[57]),
    .Tile_X27Y3_R_t(R_t_top[58]),
    .Tile_X27Y3_R_f(R_f_top[58]),
    .Tile_X30Y3_R_t(R_t_top[59]),
    .Tile_X30Y3_R_f(R_f_top[59]),
    .Tile_X33Y3_R_t(R_t_top[60]),
    .Tile_X33Y3_R_f(R_f_top[60]),
    .Tile_X36Y3_R_t(R_t_top[61]),
    .Tile_X36Y3_R_f(R_f_top[61]),
    .Tile_X39Y3_R_t(R_t_top[62]),
    .Tile_X39Y3_R_f(R_f_top[62]),
    .Tile_X42Y3_R_t(R_t_top[63]),
    .Tile_X42Y3_R_f(R_f_top[63]),
    .Tile_X45Y3_R_t(R_t_top[64]),
    .Tile_X45Y3_R_f(R_f_top[64]),
    .Tile_X48Y3_R_t(R_t_top[65]),
    .Tile_X48Y3_R_f(R_f_top[65]),
    .Tile_X51Y3_R_t(R_t_top[66]),
    .Tile_X51Y3_R_f(R_f_top[66]),
    .Tile_X54Y3_R_t(R_t_top[67]),
    .Tile_X54Y3_R_f(R_f_top[67]),
    .Tile_X57Y3_R_t(R_t_top[68]),
    .Tile_X57Y3_R_f(R_f_top[68]),
    .Tile_X60Y3_R_t(R_t_top[69]),
    .Tile_X60Y3_R_f(R_f_top[69]),
    .Tile_X63Y3_R_t(R_t_top[70]),
    .Tile_X63Y3_R_f(R_f_top[70]),
    .Tile_X66Y3_R_t(R_t_top[71]),
    .Tile_X66Y3_R_f(R_f_top[71]),
    .Tile_X69Y3_R_t(R_t_top[72]),
    .Tile_X69Y3_R_f(R_f_top[72]),
    .Tile_X72Y3_R_t(R_t_top[73]),
    .Tile_X72Y3_R_f(R_f_top[73]),
    .Tile_X75Y3_R_t(R_t_top[74]),
    .Tile_X75Y3_R_f(R_f_top[74]),
    .Tile_X3Y4_R_t(R_t_top[75]),
    .Tile_X3Y4_R_f(R_f_top[75]),
    .Tile_X6Y4_R_t(R_t_top[76]),
    .Tile_X6Y4_R_f(R_f_top[76]),
    .Tile_X9Y4_R_t(R_t_top[77]),
    .Tile_X9Y4_R_f(R_f_top[77]),
    .Tile_X12Y4_R_t(R_t_top[78]),
    .Tile_X12Y4_R_f(R_f_top[78]),
    .Tile_X15Y4_R_t(R_t_top[79]),
    .Tile_X15Y4_R_f(R_f_top[79]),
    .Tile_X18Y4_R_t(R_t_top[80]),
    .Tile_X18Y4_R_f(R_f_top[80]),
    .Tile_X21Y4_R_t(R_t_top[81]),
    .Tile_X21Y4_R_f(R_f_top[81]),
    .Tile_X24Y4_R_t(R_t_top[82]),
    .Tile_X24Y4_R_f(R_f_top[82]),
    .Tile_X27Y4_R_t(R_t_top[83]),
    .Tile_X27Y4_R_f(R_f_top[83]),
    .Tile_X30Y4_R_t(R_t_top[84]),
    .Tile_X30Y4_R_f(R_f_top[84]),
    .Tile_X33Y4_R_t(R_t_top[85]),
    .Tile_X33Y4_R_f(R_f_top[85]),
    .Tile_X36Y4_R_t(R_t_top[86]),
    .Tile_X36Y4_R_f(R_f_top[86]),
    .Tile_X39Y4_R_t(R_t_top[87]),
    .Tile_X39Y4_R_f(R_f_top[87]),
    .Tile_X42Y4_R_t(R_t_top[88]),
    .Tile_X42Y4_R_f(R_f_top[88]),
    .Tile_X45Y4_R_t(R_t_top[89]),
    .Tile_X45Y4_R_f(R_f_top[89]),
    .Tile_X48Y4_R_t(R_t_top[90]),
    .Tile_X48Y4_R_f(R_f_top[90]),
    .Tile_X51Y4_R_t(R_t_top[91]),
    .Tile_X51Y4_R_f(R_f_top[91]),
    .Tile_X54Y4_R_t(R_t_top[92]),
    .Tile_X54Y4_R_f(R_f_top[92]),
    .Tile_X57Y4_R_t(R_t_top[93]),
    .Tile_X57Y4_R_f(R_f_top[93]),
    .Tile_X60Y4_R_t(R_t_top[94]),
    .Tile_X60Y4_R_f(R_f_top[94]),
    .Tile_X63Y4_R_t(R_t_top[95]),
    .Tile_X63Y4_R_f(R_f_top[95]),
    .Tile_X66Y4_R_t(R_t_top[96]),
    .Tile_X66Y4_R_f(R_f_top[96]),
    .Tile_X69Y4_R_t(R_t_top[97]),
    .Tile_X69Y4_R_f(R_f_top[97]),
    .Tile_X72Y4_R_t(R_t_top[98]),
    .Tile_X72Y4_R_f(R_f_top[98]),
    .Tile_X75Y4_R_t(R_t_top[99]),
    .Tile_X75Y4_R_f(R_f_top[99]),
    .Tile_X3Y5_R_t(R_t_top[100]),
    .Tile_X3Y5_R_f(R_f_top[100]),
    .Tile_X6Y5_R_t(R_t_top[101]),
    .Tile_X6Y5_R_f(R_f_top[101]),
    .Tile_X9Y5_R_t(R_t_top[102]),
    .Tile_X9Y5_R_f(R_f_top[102]),
    .Tile_X12Y5_R_t(R_t_top[103]),
    .Tile_X12Y5_R_f(R_f_top[103]),
    .Tile_X15Y5_R_t(R_t_top[104]),
    .Tile_X15Y5_R_f(R_f_top[104]),
    .Tile_X18Y5_R_t(R_t_top[105]),
    .Tile_X18Y5_R_f(R_f_top[105]),
    .Tile_X21Y5_R_t(R_t_top[106]),
    .Tile_X21Y5_R_f(R_f_top[106]),
    .Tile_X24Y5_R_t(R_t_top[107]),
    .Tile_X24Y5_R_f(R_f_top[107]),
    .Tile_X27Y5_R_t(R_t_top[108]),
    .Tile_X27Y5_R_f(R_f_top[108]),
    .Tile_X30Y5_R_t(R_t_top[109]),
    .Tile_X30Y5_R_f(R_f_top[109]),
    .Tile_X33Y5_R_t(R_t_top[110]),
    .Tile_X33Y5_R_f(R_f_top[110]),
    .Tile_X36Y5_R_t(R_t_top[111]),
    .Tile_X36Y5_R_f(R_f_top[111]),
    .Tile_X39Y5_R_t(R_t_top[112]),
    .Tile_X39Y5_R_f(R_f_top[112]),
    .Tile_X42Y5_R_t(R_t_top[113]),
    .Tile_X42Y5_R_f(R_f_top[113]),
    .Tile_X45Y5_R_t(R_t_top[114]),
    .Tile_X45Y5_R_f(R_f_top[114]),
    .Tile_X48Y5_R_t(R_t_top[115]),
    .Tile_X48Y5_R_f(R_f_top[115]),
    .Tile_X51Y5_R_t(R_t_top[116]),
    .Tile_X51Y5_R_f(R_f_top[116]),
    .Tile_X54Y5_R_t(R_t_top[117]),
    .Tile_X54Y5_R_f(R_f_top[117]),
    .Tile_X57Y5_R_t(R_t_top[118]),
    .Tile_X57Y5_R_f(R_f_top[118]),
    .Tile_X60Y5_R_t(R_t_top[119]),
    .Tile_X60Y5_R_f(R_f_top[119]),
    .Tile_X63Y5_R_t(R_t_top[120]),
    .Tile_X63Y5_R_f(R_f_top[120]),
    .Tile_X66Y5_R_t(R_t_top[121]),
    .Tile_X66Y5_R_f(R_f_top[121]),
    .Tile_X69Y5_R_t(R_t_top[122]),
    .Tile_X69Y5_R_f(R_f_top[122]),
    .Tile_X72Y5_R_t(R_t_top[123]),
    .Tile_X72Y5_R_f(R_f_top[123]),
    .Tile_X75Y5_R_t(R_t_top[124]),
    .Tile_X75Y5_R_f(R_f_top[124]),
    .Tile_X3Y6_R_t(R_t_top[125]),
    .Tile_X3Y6_R_f(R_f_top[125]),
    .Tile_X6Y6_R_t(R_t_top[126]),
    .Tile_X6Y6_R_f(R_f_top[126]),
    .Tile_X9Y6_R_t(R_t_top[127]),
    .Tile_X9Y6_R_f(R_f_top[127]),
    .Tile_X12Y6_R_t(R_t_top[128]),
    .Tile_X12Y6_R_f(R_f_top[128]),
    .Tile_X15Y6_R_t(R_t_top[129]),
    .Tile_X15Y6_R_f(R_f_top[129]),
    .Tile_X18Y6_R_t(R_t_top[130]),
    .Tile_X18Y6_R_f(R_f_top[130]),
    .Tile_X21Y6_R_t(R_t_top[131]),
    .Tile_X21Y6_R_f(R_f_top[131]),
    .Tile_X24Y6_R_t(R_t_top[132]),
    .Tile_X24Y6_R_f(R_f_top[132]),
    .Tile_X27Y6_R_t(R_t_top[133]),
    .Tile_X27Y6_R_f(R_f_top[133]),
    .Tile_X30Y6_R_t(R_t_top[134]),
    .Tile_X30Y6_R_f(R_f_top[134]),
    .Tile_X33Y6_R_t(R_t_top[135]),
    .Tile_X33Y6_R_f(R_f_top[135]),
    .Tile_X36Y6_R_t(R_t_top[136]),
    .Tile_X36Y6_R_f(R_f_top[136]),
    .Tile_X39Y6_R_t(R_t_top[137]),
    .Tile_X39Y6_R_f(R_f_top[137]),
    .Tile_X42Y6_R_t(R_t_top[138]),
    .Tile_X42Y6_R_f(R_f_top[138]),
    .Tile_X45Y6_R_t(R_t_top[139]),
    .Tile_X45Y6_R_f(R_f_top[139]),
    .Tile_X48Y6_R_t(R_t_top[140]),
    .Tile_X48Y6_R_f(R_f_top[140]),
    .Tile_X51Y6_R_t(R_t_top[141]),
    .Tile_X51Y6_R_f(R_f_top[141]),
    .Tile_X54Y6_R_t(R_t_top[142]),
    .Tile_X54Y6_R_f(R_f_top[142]),
    .Tile_X57Y6_R_t(R_t_top[143]),
    .Tile_X57Y6_R_f(R_f_top[143]),
    .Tile_X60Y6_R_t(R_t_top[144]),
    .Tile_X60Y6_R_f(R_f_top[144]),
    .Tile_X63Y6_R_t(R_t_top[145]),
    .Tile_X63Y6_R_f(R_f_top[145]),
    .Tile_X66Y6_R_t(R_t_top[146]),
    .Tile_X66Y6_R_f(R_f_top[146]),
    .Tile_X69Y6_R_t(R_t_top[147]),
    .Tile_X69Y6_R_f(R_f_top[147]),
    .Tile_X72Y6_R_t(R_t_top[148]),
    .Tile_X72Y6_R_f(R_f_top[148]),
    .Tile_X75Y6_R_t(R_t_top[149]),
    .Tile_X75Y6_R_f(R_f_top[149]),
    .Tile_X3Y7_R_t(R_t_top[150]),
    .Tile_X3Y7_R_f(R_f_top[150]),
    .Tile_X6Y7_R_t(R_t_top[151]),
    .Tile_X6Y7_R_f(R_f_top[151]),
    .Tile_X9Y7_R_t(R_t_top[152]),
    .Tile_X9Y7_R_f(R_f_top[152]),
    .Tile_X12Y7_R_t(R_t_top[153]),
    .Tile_X12Y7_R_f(R_f_top[153]),
    .Tile_X15Y7_R_t(R_t_top[154]),
    .Tile_X15Y7_R_f(R_f_top[154]),
    .Tile_X18Y7_R_t(R_t_top[155]),
    .Tile_X18Y7_R_f(R_f_top[155]),
    .Tile_X21Y7_R_t(R_t_top[156]),
    .Tile_X21Y7_R_f(R_f_top[156]),
    .Tile_X24Y7_R_t(R_t_top[157]),
    .Tile_X24Y7_R_f(R_f_top[157]),
    .Tile_X27Y7_R_t(R_t_top[158]),
    .Tile_X27Y7_R_f(R_f_top[158]),
    .Tile_X30Y7_R_t(R_t_top[159]),
    .Tile_X30Y7_R_f(R_f_top[159]),
    .Tile_X33Y7_R_t(R_t_top[160]),
    .Tile_X33Y7_R_f(R_f_top[160]),
    .Tile_X36Y7_R_t(R_t_top[161]),
    .Tile_X36Y7_R_f(R_f_top[161]),
    .Tile_X39Y7_R_t(R_t_top[162]),
    .Tile_X39Y7_R_f(R_f_top[162]),
    .Tile_X42Y7_R_t(R_t_top[163]),
    .Tile_X42Y7_R_f(R_f_top[163]),
    .Tile_X45Y7_R_t(R_t_top[164]),
    .Tile_X45Y7_R_f(R_f_top[164]),
    .Tile_X48Y7_R_t(R_t_top[165]),
    .Tile_X48Y7_R_f(R_f_top[165]),
    .Tile_X51Y7_R_t(R_t_top[166]),
    .Tile_X51Y7_R_f(R_f_top[166]),
    .Tile_X54Y7_R_t(R_t_top[167]),
    .Tile_X54Y7_R_f(R_f_top[167]),
    .Tile_X57Y7_R_t(R_t_top[168]),
    .Tile_X57Y7_R_f(R_f_top[168]),
    .Tile_X60Y7_R_t(R_t_top[169]),
    .Tile_X60Y7_R_f(R_f_top[169]),
    .Tile_X63Y7_R_t(R_t_top[170]),
    .Tile_X63Y7_R_f(R_f_top[170]),
    .Tile_X66Y7_R_t(R_t_top[171]),
    .Tile_X66Y7_R_f(R_f_top[171]),
    .Tile_X69Y7_R_t(R_t_top[172]),
    .Tile_X69Y7_R_f(R_f_top[172]),
    .Tile_X72Y7_R_t(R_t_top[173]),
    .Tile_X72Y7_R_f(R_f_top[173]),
    .Tile_X75Y7_R_t(R_t_top[174]),
    .Tile_X75Y7_R_f(R_f_top[174]),
    .Tile_X3Y8_R_t(R_t_top[175]),
    .Tile_X3Y8_R_f(R_f_top[175]),
    .Tile_X6Y8_R_t(R_t_top[176]),
    .Tile_X6Y8_R_f(R_f_top[176]),
    .Tile_X9Y8_R_t(R_t_top[177]),
    .Tile_X9Y8_R_f(R_f_top[177]),
    .Tile_X12Y8_R_t(R_t_top[178]),
    .Tile_X12Y8_R_f(R_f_top[178]),
    .Tile_X15Y8_R_t(R_t_top[179]),
    .Tile_X15Y8_R_f(R_f_top[179]),
    .Tile_X18Y8_R_t(R_t_top[180]),
    .Tile_X18Y8_R_f(R_f_top[180]),
    .Tile_X21Y8_R_t(R_t_top[181]),
    .Tile_X21Y8_R_f(R_f_top[181]),
    .Tile_X24Y8_R_t(R_t_top[182]),
    .Tile_X24Y8_R_f(R_f_top[182]),
    .Tile_X27Y8_R_t(R_t_top[183]),
    .Tile_X27Y8_R_f(R_f_top[183]),
    .Tile_X30Y8_R_t(R_t_top[184]),
    .Tile_X30Y8_R_f(R_f_top[184]),
    .Tile_X33Y8_R_t(R_t_top[185]),
    .Tile_X33Y8_R_f(R_f_top[185]),
    .Tile_X36Y8_R_t(R_t_top[186]),
    .Tile_X36Y8_R_f(R_f_top[186]),
    .Tile_X39Y8_R_t(R_t_top[187]),
    .Tile_X39Y8_R_f(R_f_top[187]),
    .Tile_X42Y8_R_t(R_t_top[188]),
    .Tile_X42Y8_R_f(R_f_top[188]),
    .Tile_X45Y8_R_t(R_t_top[189]),
    .Tile_X45Y8_R_f(R_f_top[189]),
    .Tile_X48Y8_R_t(R_t_top[190]),
    .Tile_X48Y8_R_f(R_f_top[190]),
    .Tile_X51Y8_R_t(R_t_top[191]),
    .Tile_X51Y8_R_f(R_f_top[191]),
    .Tile_X54Y8_R_t(R_t_top[192]),
    .Tile_X54Y8_R_f(R_f_top[192]),
    .Tile_X57Y8_R_t(R_t_top[193]),
    .Tile_X57Y8_R_f(R_f_top[193]),
    .Tile_X60Y8_R_t(R_t_top[194]),
    .Tile_X60Y8_R_f(R_f_top[194]),
    .Tile_X63Y8_R_t(R_t_top[195]),
    .Tile_X63Y8_R_f(R_f_top[195]),
    .Tile_X66Y8_R_t(R_t_top[196]),
    .Tile_X66Y8_R_f(R_f_top[196]),
    .Tile_X69Y8_R_t(R_t_top[197]),
    .Tile_X69Y8_R_f(R_f_top[197]),
    .Tile_X72Y8_R_t(R_t_top[198]),
    .Tile_X72Y8_R_f(R_f_top[198]),
    .Tile_X75Y8_R_t(R_t_top[199]),
    .Tile_X75Y8_R_f(R_f_top[199]),
    .Tile_X3Y9_R_t(R_t_top[200]),
    .Tile_X3Y9_R_f(R_f_top[200]),
    .Tile_X6Y9_R_t(R_t_top[201]),
    .Tile_X6Y9_R_f(R_f_top[201]),
    .Tile_X9Y9_R_t(R_t_top[202]),
    .Tile_X9Y9_R_f(R_f_top[202]),
    .Tile_X12Y9_R_t(R_t_top[203]),
    .Tile_X12Y9_R_f(R_f_top[203]),
    .Tile_X15Y9_R_t(R_t_top[204]),
    .Tile_X15Y9_R_f(R_f_top[204]),
    .Tile_X18Y9_R_t(R_t_top[205]),
    .Tile_X18Y9_R_f(R_f_top[205]),
    .Tile_X21Y9_R_t(R_t_top[206]),
    .Tile_X21Y9_R_f(R_f_top[206]),
    .Tile_X24Y9_R_t(R_t_top[207]),
    .Tile_X24Y9_R_f(R_f_top[207]),
    .Tile_X27Y9_R_t(R_t_top[208]),
    .Tile_X27Y9_R_f(R_f_top[208]),
    .Tile_X30Y9_R_t(R_t_top[209]),
    .Tile_X30Y9_R_f(R_f_top[209]),
    .Tile_X33Y9_R_t(R_t_top[210]),
    .Tile_X33Y9_R_f(R_f_top[210]),
    .Tile_X36Y9_R_t(R_t_top[211]),
    .Tile_X36Y9_R_f(R_f_top[211]),
    .Tile_X39Y9_R_t(R_t_top[212]),
    .Tile_X39Y9_R_f(R_f_top[212]),
    .Tile_X42Y9_R_t(R_t_top[213]),
    .Tile_X42Y9_R_f(R_f_top[213]),
    .Tile_X45Y9_R_t(R_t_top[214]),
    .Tile_X45Y9_R_f(R_f_top[214]),
    .Tile_X48Y9_R_t(R_t_top[215]),
    .Tile_X48Y9_R_f(R_f_top[215]),
    .Tile_X51Y9_R_t(R_t_top[216]),
    .Tile_X51Y9_R_f(R_f_top[216]),
    .Tile_X54Y9_R_t(R_t_top[217]),
    .Tile_X54Y9_R_f(R_f_top[217]),
    .Tile_X57Y9_R_t(R_t_top[218]),
    .Tile_X57Y9_R_f(R_f_top[218]),
    .Tile_X60Y9_R_t(R_t_top[219]),
    .Tile_X60Y9_R_f(R_f_top[219]),
    .Tile_X63Y9_R_t(R_t_top[220]),
    .Tile_X63Y9_R_f(R_f_top[220]),
    .Tile_X66Y9_R_t(R_t_top[221]),
    .Tile_X66Y9_R_f(R_f_top[221]),
    .Tile_X69Y9_R_t(R_t_top[222]),
    .Tile_X69Y9_R_f(R_f_top[222]),
    .Tile_X72Y9_R_t(R_t_top[223]),
    .Tile_X72Y9_R_f(R_f_top[223]),
    .Tile_X75Y9_R_t(R_t_top[224]),
    .Tile_X75Y9_R_f(R_f_top[224]),
    .Tile_X3Y10_R_t(R_t_top[225]),
    .Tile_X3Y10_R_f(R_f_top[225]),
    .Tile_X6Y10_R_t(R_t_top[226]),
    .Tile_X6Y10_R_f(R_f_top[226]),
    .Tile_X9Y10_R_t(R_t_top[227]),
    .Tile_X9Y10_R_f(R_f_top[227]),
    .Tile_X12Y10_R_t(R_t_top[228]),
    .Tile_X12Y10_R_f(R_f_top[228]),
    .Tile_X15Y10_R_t(R_t_top[229]),
    .Tile_X15Y10_R_f(R_f_top[229]),
    .Tile_X18Y10_R_t(R_t_top[230]),
    .Tile_X18Y10_R_f(R_f_top[230]),
    .Tile_X21Y10_R_t(R_t_top[231]),
    .Tile_X21Y10_R_f(R_f_top[231]),
    .Tile_X24Y10_R_t(R_t_top[232]),
    .Tile_X24Y10_R_f(R_f_top[232]),
    .Tile_X27Y10_R_t(R_t_top[233]),
    .Tile_X27Y10_R_f(R_f_top[233]),
    .Tile_X30Y10_R_t(R_t_top[234]),
    .Tile_X30Y10_R_f(R_f_top[234]),
    .Tile_X33Y10_R_t(R_t_top[235]),
    .Tile_X33Y10_R_f(R_f_top[235]),
    .Tile_X36Y10_R_t(R_t_top[236]),
    .Tile_X36Y10_R_f(R_f_top[236]),
    .Tile_X39Y10_R_t(R_t_top[237]),
    .Tile_X39Y10_R_f(R_f_top[237]),
    .Tile_X42Y10_R_t(R_t_top[238]),
    .Tile_X42Y10_R_f(R_f_top[238]),
    .Tile_X45Y10_R_t(R_t_top[239]),
    .Tile_X45Y10_R_f(R_f_top[239]),
    .Tile_X48Y10_R_t(R_t_top[240]),
    .Tile_X48Y10_R_f(R_f_top[240]),
    .Tile_X51Y10_R_t(R_t_top[241]),
    .Tile_X51Y10_R_f(R_f_top[241]),
    .Tile_X54Y10_R_t(R_t_top[242]),
    .Tile_X54Y10_R_f(R_f_top[242]),
    .Tile_X57Y10_R_t(R_t_top[243]),
    .Tile_X57Y10_R_f(R_f_top[243]),
    .Tile_X60Y10_R_t(R_t_top[244]),
    .Tile_X60Y10_R_f(R_f_top[244]),
    .Tile_X63Y10_R_t(R_t_top[245]),
    .Tile_X63Y10_R_f(R_f_top[245]),
    .Tile_X66Y10_R_t(R_t_top[246]),
    .Tile_X66Y10_R_f(R_f_top[246]),
    .Tile_X69Y10_R_t(R_t_top[247]),
    .Tile_X69Y10_R_f(R_f_top[247]),
    .Tile_X72Y10_R_t(R_t_top[248]),
    .Tile_X72Y10_R_f(R_f_top[248]),
    .Tile_X75Y10_R_t(R_t_top[249]),
    .Tile_X75Y10_R_f(R_f_top[249]),
    .Tile_X3Y11_R_t(R_t_top[250]),
    .Tile_X3Y11_R_f(R_f_top[250]),
    .Tile_X6Y11_R_t(R_t_top[251]),
    .Tile_X6Y11_R_f(R_f_top[251]),
    .Tile_X9Y11_R_t(R_t_top[252]),
    .Tile_X9Y11_R_f(R_f_top[252]),
    .Tile_X12Y11_R_t(R_t_top[253]),
    .Tile_X12Y11_R_f(R_f_top[253]),
    .Tile_X15Y11_R_t(R_t_top[254]),
    .Tile_X15Y11_R_f(R_f_top[254]),
    .Tile_X18Y11_R_t(R_t_top[255]),
    .Tile_X18Y11_R_f(R_f_top[255]),
    .Tile_X21Y11_R_t(R_t_top[256]),
    .Tile_X21Y11_R_f(R_f_top[256]),
    .Tile_X24Y11_R_t(R_t_top[257]),
    .Tile_X24Y11_R_f(R_f_top[257]),
    .Tile_X27Y11_R_t(R_t_top[258]),
    .Tile_X27Y11_R_f(R_f_top[258]),
    .Tile_X30Y11_R_t(R_t_top[259]),
    .Tile_X30Y11_R_f(R_f_top[259]),
    .Tile_X33Y11_R_t(R_t_top[260]),
    .Tile_X33Y11_R_f(R_f_top[260]),
    .Tile_X36Y11_R_t(R_t_top[261]),
    .Tile_X36Y11_R_f(R_f_top[261]),
    .Tile_X39Y11_R_t(R_t_top[262]),
    .Tile_X39Y11_R_f(R_f_top[262]),
    .Tile_X42Y11_R_t(R_t_top[263]),
    .Tile_X42Y11_R_f(R_f_top[263]),
    .Tile_X45Y11_R_t(R_t_top[264]),
    .Tile_X45Y11_R_f(R_f_top[264]),
    .Tile_X48Y11_R_t(R_t_top[265]),
    .Tile_X48Y11_R_f(R_f_top[265]),
    .Tile_X51Y11_R_t(R_t_top[266]),
    .Tile_X51Y11_R_f(R_f_top[266]),
    .Tile_X54Y11_R_t(R_t_top[267]),
    .Tile_X54Y11_R_f(R_f_top[267]),
    .Tile_X57Y11_R_t(R_t_top[268]),
    .Tile_X57Y11_R_f(R_f_top[268]),
    .Tile_X60Y11_R_t(R_t_top[269]),
    .Tile_X60Y11_R_f(R_f_top[269]),
    .Tile_X63Y11_R_t(R_t_top[270]),
    .Tile_X63Y11_R_f(R_f_top[270]),
    .Tile_X66Y11_R_t(R_t_top[271]),
    .Tile_X66Y11_R_f(R_f_top[271]),
    .Tile_X69Y11_R_t(R_t_top[272]),
    .Tile_X69Y11_R_f(R_f_top[272]),
    .Tile_X72Y11_R_t(R_t_top[273]),
    .Tile_X72Y11_R_f(R_f_top[273]),
    .Tile_X75Y11_R_t(R_t_top[274]),
    .Tile_X75Y11_R_f(R_f_top[274]),
    .Tile_X3Y12_R_t(R_t_top[275]),
    .Tile_X3Y12_R_f(R_f_top[275]),
    .Tile_X6Y12_R_t(R_t_top[276]),
    .Tile_X6Y12_R_f(R_f_top[276]),
    .Tile_X9Y12_R_t(R_t_top[277]),
    .Tile_X9Y12_R_f(R_f_top[277]),
    .Tile_X12Y12_R_t(R_t_top[278]),
    .Tile_X12Y12_R_f(R_f_top[278]),
    .Tile_X15Y12_R_t(R_t_top[279]),
    .Tile_X15Y12_R_f(R_f_top[279]),
    .Tile_X18Y12_R_t(R_t_top[280]),
    .Tile_X18Y12_R_f(R_f_top[280]),
    .Tile_X21Y12_R_t(R_t_top[281]),
    .Tile_X21Y12_R_f(R_f_top[281]),
    .Tile_X24Y12_R_t(R_t_top[282]),
    .Tile_X24Y12_R_f(R_f_top[282]),
    .Tile_X27Y12_R_t(R_t_top[283]),
    .Tile_X27Y12_R_f(R_f_top[283]),
    .Tile_X30Y12_R_t(R_t_top[284]),
    .Tile_X30Y12_R_f(R_f_top[284]),
    .Tile_X33Y12_R_t(R_t_top[285]),
    .Tile_X33Y12_R_f(R_f_top[285]),
    .Tile_X36Y12_R_t(R_t_top[286]),
    .Tile_X36Y12_R_f(R_f_top[286]),
    .Tile_X39Y12_R_t(R_t_top[287]),
    .Tile_X39Y12_R_f(R_f_top[287]),
    .Tile_X42Y12_R_t(R_t_top[288]),
    .Tile_X42Y12_R_f(R_f_top[288]),
    .Tile_X45Y12_R_t(R_t_top[289]),
    .Tile_X45Y12_R_f(R_f_top[289]),
    .Tile_X48Y12_R_t(R_t_top[290]),
    .Tile_X48Y12_R_f(R_f_top[290]),
    .Tile_X51Y12_R_t(R_t_top[291]),
    .Tile_X51Y12_R_f(R_f_top[291]),
    .Tile_X54Y12_R_t(R_t_top[292]),
    .Tile_X54Y12_R_f(R_f_top[292]),
    .Tile_X57Y12_R_t(R_t_top[293]),
    .Tile_X57Y12_R_f(R_f_top[293]),
    .Tile_X60Y12_R_t(R_t_top[294]),
    .Tile_X60Y12_R_f(R_f_top[294]),
    .Tile_X63Y12_R_t(R_t_top[295]),
    .Tile_X63Y12_R_f(R_f_top[295]),
    .Tile_X66Y12_R_t(R_t_top[296]),
    .Tile_X66Y12_R_f(R_f_top[296]),
    .Tile_X69Y12_R_t(R_t_top[297]),
    .Tile_X69Y12_R_f(R_f_top[297]),
    .Tile_X72Y12_R_t(R_t_top[298]),
    .Tile_X72Y12_R_f(R_f_top[298]),
    .Tile_X75Y12_R_t(R_t_top[299]),
    .Tile_X75Y12_R_f(R_f_top[299]),
    .Tile_X3Y13_R_t(R_t_top[300]),
    .Tile_X3Y13_R_f(R_f_top[300]),
    .Tile_X6Y13_R_t(R_t_top[301]),
    .Tile_X6Y13_R_f(R_f_top[301]),
    .Tile_X9Y13_R_t(R_t_top[302]),
    .Tile_X9Y13_R_f(R_f_top[302]),
    .Tile_X12Y13_R_t(R_t_top[303]),
    .Tile_X12Y13_R_f(R_f_top[303]),
    .Tile_X15Y13_R_t(R_t_top[304]),
    .Tile_X15Y13_R_f(R_f_top[304]),
    .Tile_X18Y13_R_t(R_t_top[305]),
    .Tile_X18Y13_R_f(R_f_top[305]),
    .Tile_X21Y13_R_t(R_t_top[306]),
    .Tile_X21Y13_R_f(R_f_top[306]),
    .Tile_X24Y13_R_t(R_t_top[307]),
    .Tile_X24Y13_R_f(R_f_top[307]),
    .Tile_X27Y13_R_t(R_t_top[308]),
    .Tile_X27Y13_R_f(R_f_top[308]),
    .Tile_X30Y13_R_t(R_t_top[309]),
    .Tile_X30Y13_R_f(R_f_top[309]),
    .Tile_X33Y13_R_t(R_t_top[310]),
    .Tile_X33Y13_R_f(R_f_top[310]),
    .Tile_X36Y13_R_t(R_t_top[311]),
    .Tile_X36Y13_R_f(R_f_top[311]),
    .Tile_X39Y13_R_t(R_t_top[312]),
    .Tile_X39Y13_R_f(R_f_top[312]),
    .Tile_X42Y13_R_t(R_t_top[313]),
    .Tile_X42Y13_R_f(R_f_top[313]),
    .Tile_X45Y13_R_t(R_t_top[314]),
    .Tile_X45Y13_R_f(R_f_top[314]),
    .Tile_X48Y13_R_t(R_t_top[315]),
    .Tile_X48Y13_R_f(R_f_top[315]),
    .Tile_X51Y13_R_t(R_t_top[316]),
    .Tile_X51Y13_R_f(R_f_top[316]),
    .Tile_X54Y13_R_t(R_t_top[317]),
    .Tile_X54Y13_R_f(R_f_top[317]),
    .Tile_X57Y13_R_t(R_t_top[318]),
    .Tile_X57Y13_R_f(R_f_top[318]),
    .Tile_X60Y13_R_t(R_t_top[319]),
    .Tile_X60Y13_R_f(R_f_top[319]),
    .Tile_X63Y13_R_t(R_t_top[320]),
    .Tile_X63Y13_R_f(R_f_top[320]),
    .Tile_X66Y13_R_t(R_t_top[321]),
    .Tile_X66Y13_R_f(R_f_top[321]),
    .Tile_X69Y13_R_t(R_t_top[322]),
    .Tile_X69Y13_R_f(R_f_top[322]),
    .Tile_X72Y13_R_t(R_t_top[323]),
    .Tile_X72Y13_R_f(R_f_top[323]),
    .Tile_X75Y13_R_t(R_t_top[324]),
    .Tile_X75Y13_R_f(R_f_top[324]),
    .Tile_X3Y14_R_t(R_t_top[325]),
    .Tile_X3Y14_R_f(R_f_top[325]),
    .Tile_X6Y14_R_t(R_t_top[326]),
    .Tile_X6Y14_R_f(R_f_top[326]),
    .Tile_X9Y14_R_t(R_t_top[327]),
    .Tile_X9Y14_R_f(R_f_top[327]),
    .Tile_X12Y14_R_t(R_t_top[328]),
    .Tile_X12Y14_R_f(R_f_top[328]),
    .Tile_X15Y14_R_t(R_t_top[329]),
    .Tile_X15Y14_R_f(R_f_top[329]),
    .Tile_X18Y14_R_t(R_t_top[330]),
    .Tile_X18Y14_R_f(R_f_top[330]),
    .Tile_X21Y14_R_t(R_t_top[331]),
    .Tile_X21Y14_R_f(R_f_top[331]),
    .Tile_X24Y14_R_t(R_t_top[332]),
    .Tile_X24Y14_R_f(R_f_top[332]),
    .Tile_X27Y14_R_t(R_t_top[333]),
    .Tile_X27Y14_R_f(R_f_top[333]),
    .Tile_X30Y14_R_t(R_t_top[334]),
    .Tile_X30Y14_R_f(R_f_top[334]),
    .Tile_X33Y14_R_t(R_t_top[335]),
    .Tile_X33Y14_R_f(R_f_top[335]),
    .Tile_X36Y14_R_t(R_t_top[336]),
    .Tile_X36Y14_R_f(R_f_top[336]),
    .Tile_X39Y14_R_t(R_t_top[337]),
    .Tile_X39Y14_R_f(R_f_top[337]),
    .Tile_X42Y14_R_t(R_t_top[338]),
    .Tile_X42Y14_R_f(R_f_top[338]),
    .Tile_X45Y14_R_t(R_t_top[339]),
    .Tile_X45Y14_R_f(R_f_top[339]),
    .Tile_X48Y14_R_t(R_t_top[340]),
    .Tile_X48Y14_R_f(R_f_top[340]),
    .Tile_X51Y14_R_t(R_t_top[341]),
    .Tile_X51Y14_R_f(R_f_top[341]),
    .Tile_X54Y14_R_t(R_t_top[342]),
    .Tile_X54Y14_R_f(R_f_top[342]),
    .Tile_X57Y14_R_t(R_t_top[343]),
    .Tile_X57Y14_R_f(R_f_top[343]),
    .Tile_X60Y14_R_t(R_t_top[344]),
    .Tile_X60Y14_R_f(R_f_top[344]),
    .Tile_X63Y14_R_t(R_t_top[345]),
    .Tile_X63Y14_R_f(R_f_top[345]),
    .Tile_X66Y14_R_t(R_t_top[346]),
    .Tile_X66Y14_R_f(R_f_top[346]),
    .Tile_X69Y14_R_t(R_t_top[347]),
    .Tile_X69Y14_R_f(R_f_top[347]),
    .Tile_X72Y14_R_t(R_t_top[348]),
    .Tile_X72Y14_R_f(R_f_top[348]),
    .Tile_X75Y14_R_t(R_t_top[349]),
    .Tile_X75Y14_R_f(R_f_top[349]),
    .Tile_X3Y15_R_t(R_t_top[350]),
    .Tile_X3Y15_R_f(R_f_top[350]),
    .Tile_X6Y15_R_t(R_t_top[351]),
    .Tile_X6Y15_R_f(R_f_top[351]),
    .Tile_X9Y15_R_t(R_t_top[352]),
    .Tile_X9Y15_R_f(R_f_top[352]),
    .Tile_X12Y15_R_t(R_t_top[353]),
    .Tile_X12Y15_R_f(R_f_top[353]),
    .Tile_X15Y15_R_t(R_t_top[354]),
    .Tile_X15Y15_R_f(R_f_top[354]),
    .Tile_X18Y15_R_t(R_t_top[355]),
    .Tile_X18Y15_R_f(R_f_top[355]),
    .Tile_X21Y15_R_t(R_t_top[356]),
    .Tile_X21Y15_R_f(R_f_top[356]),
    .Tile_X24Y15_R_t(R_t_top[357]),
    .Tile_X24Y15_R_f(R_f_top[357]),
    .Tile_X27Y15_R_t(R_t_top[358]),
    .Tile_X27Y15_R_f(R_f_top[358]),
    .Tile_X30Y15_R_t(R_t_top[359]),
    .Tile_X30Y15_R_f(R_f_top[359]),
    .Tile_X33Y15_R_t(R_t_top[360]),
    .Tile_X33Y15_R_f(R_f_top[360]),
    .Tile_X36Y15_R_t(R_t_top[361]),
    .Tile_X36Y15_R_f(R_f_top[361]),
    .Tile_X39Y15_R_t(R_t_top[362]),
    .Tile_X39Y15_R_f(R_f_top[362]),
    .Tile_X42Y15_R_t(R_t_top[363]),
    .Tile_X42Y15_R_f(R_f_top[363]),
    .Tile_X45Y15_R_t(R_t_top[364]),
    .Tile_X45Y15_R_f(R_f_top[364]),
    .Tile_X48Y15_R_t(R_t_top[365]),
    .Tile_X48Y15_R_f(R_f_top[365]),
    .Tile_X51Y15_R_t(R_t_top[366]),
    .Tile_X51Y15_R_f(R_f_top[366]),
    .Tile_X54Y15_R_t(R_t_top[367]),
    .Tile_X54Y15_R_f(R_f_top[367]),
    .Tile_X57Y15_R_t(R_t_top[368]),
    .Tile_X57Y15_R_f(R_f_top[368]),
    .Tile_X60Y15_R_t(R_t_top[369]),
    .Tile_X60Y15_R_f(R_f_top[369]),
    .Tile_X63Y15_R_t(R_t_top[370]),
    .Tile_X63Y15_R_f(R_f_top[370]),
    .Tile_X66Y15_R_t(R_t_top[371]),
    .Tile_X66Y15_R_f(R_f_top[371]),
    .Tile_X69Y15_R_t(R_t_top[372]),
    .Tile_X69Y15_R_f(R_f_top[372]),
    .Tile_X72Y15_R_t(R_t_top[373]),
    .Tile_X72Y15_R_f(R_f_top[373]),
    .Tile_X75Y15_R_t(R_t_top[374]),
    .Tile_X75Y15_R_f(R_f_top[374]),
    .Tile_X3Y16_R_t(R_t_top[375]),
    .Tile_X3Y16_R_f(R_f_top[375]),
    .Tile_X6Y16_R_t(R_t_top[376]),
    .Tile_X6Y16_R_f(R_f_top[376]),
    .Tile_X9Y16_R_t(R_t_top[377]),
    .Tile_X9Y16_R_f(R_f_top[377]),
    .Tile_X12Y16_R_t(R_t_top[378]),
    .Tile_X12Y16_R_f(R_f_top[378]),
    .Tile_X15Y16_R_t(R_t_top[379]),
    .Tile_X15Y16_R_f(R_f_top[379]),
    .Tile_X18Y16_R_t(R_t_top[380]),
    .Tile_X18Y16_R_f(R_f_top[380]),
    .Tile_X21Y16_R_t(R_t_top[381]),
    .Tile_X21Y16_R_f(R_f_top[381]),
    .Tile_X24Y16_R_t(R_t_top[382]),
    .Tile_X24Y16_R_f(R_f_top[382]),
    .Tile_X27Y16_R_t(R_t_top[383]),
    .Tile_X27Y16_R_f(R_f_top[383]),
    .Tile_X30Y16_R_t(R_t_top[384]),
    .Tile_X30Y16_R_f(R_f_top[384]),
    .Tile_X33Y16_R_t(R_t_top[385]),
    .Tile_X33Y16_R_f(R_f_top[385]),
    .Tile_X36Y16_R_t(R_t_top[386]),
    .Tile_X36Y16_R_f(R_f_top[386]),
    .Tile_X39Y16_R_t(R_t_top[387]),
    .Tile_X39Y16_R_f(R_f_top[387]),
    .Tile_X42Y16_R_t(R_t_top[388]),
    .Tile_X42Y16_R_f(R_f_top[388]),
    .Tile_X45Y16_R_t(R_t_top[389]),
    .Tile_X45Y16_R_f(R_f_top[389]),
    .Tile_X48Y16_R_t(R_t_top[390]),
    .Tile_X48Y16_R_f(R_f_top[390]),
    .Tile_X51Y16_R_t(R_t_top[391]),
    .Tile_X51Y16_R_f(R_f_top[391]),
    .Tile_X54Y16_R_t(R_t_top[392]),
    .Tile_X54Y16_R_f(R_f_top[392]),
    .Tile_X57Y16_R_t(R_t_top[393]),
    .Tile_X57Y16_R_f(R_f_top[393]),
    .Tile_X60Y16_R_t(R_t_top[394]),
    .Tile_X60Y16_R_f(R_f_top[394]),
    .Tile_X63Y16_R_t(R_t_top[395]),
    .Tile_X63Y16_R_f(R_f_top[395]),
    .Tile_X66Y16_R_t(R_t_top[396]),
    .Tile_X66Y16_R_f(R_f_top[396]),
    .Tile_X69Y16_R_t(R_t_top[397]),
    .Tile_X69Y16_R_f(R_f_top[397]),
    .Tile_X72Y16_R_t(R_t_top[398]),
    .Tile_X72Y16_R_f(R_f_top[398]),
    .Tile_X75Y16_R_t(R_t_top[399]),
    .Tile_X75Y16_R_f(R_f_top[399]),
    .Tile_X3Y17_R_t(R_t_top[400]),
    .Tile_X3Y17_R_f(R_f_top[400]),
    .Tile_X6Y17_R_t(R_t_top[401]),
    .Tile_X6Y17_R_f(R_f_top[401]),
    .Tile_X9Y17_R_t(R_t_top[402]),
    .Tile_X9Y17_R_f(R_f_top[402]),
    .Tile_X12Y17_R_t(R_t_top[403]),
    .Tile_X12Y17_R_f(R_f_top[403]),
    .Tile_X15Y17_R_t(R_t_top[404]),
    .Tile_X15Y17_R_f(R_f_top[404]),
    .Tile_X18Y17_R_t(R_t_top[405]),
    .Tile_X18Y17_R_f(R_f_top[405]),
    .Tile_X21Y17_R_t(R_t_top[406]),
    .Tile_X21Y17_R_f(R_f_top[406]),
    .Tile_X24Y17_R_t(R_t_top[407]),
    .Tile_X24Y17_R_f(R_f_top[407]),
    .Tile_X27Y17_R_t(R_t_top[408]),
    .Tile_X27Y17_R_f(R_f_top[408]),
    .Tile_X30Y17_R_t(R_t_top[409]),
    .Tile_X30Y17_R_f(R_f_top[409]),
    .Tile_X33Y17_R_t(R_t_top[410]),
    .Tile_X33Y17_R_f(R_f_top[410]),
    .Tile_X36Y17_R_t(R_t_top[411]),
    .Tile_X36Y17_R_f(R_f_top[411]),
    .Tile_X39Y17_R_t(R_t_top[412]),
    .Tile_X39Y17_R_f(R_f_top[412]),
    .Tile_X42Y17_R_t(R_t_top[413]),
    .Tile_X42Y17_R_f(R_f_top[413]),
    .Tile_X45Y17_R_t(R_t_top[414]),
    .Tile_X45Y17_R_f(R_f_top[414]),
    .Tile_X48Y17_R_t(R_t_top[415]),
    .Tile_X48Y17_R_f(R_f_top[415]),
    .Tile_X51Y17_R_t(R_t_top[416]),
    .Tile_X51Y17_R_f(R_f_top[416]),
    .Tile_X54Y17_R_t(R_t_top[417]),
    .Tile_X54Y17_R_f(R_f_top[417]),
    .Tile_X57Y17_R_t(R_t_top[418]),
    .Tile_X57Y17_R_f(R_f_top[418]),
    .Tile_X60Y17_R_t(R_t_top[419]),
    .Tile_X60Y17_R_f(R_f_top[419]),
    .Tile_X63Y17_R_t(R_t_top[420]),
    .Tile_X63Y17_R_f(R_f_top[420]),
    .Tile_X66Y17_R_t(R_t_top[421]),
    .Tile_X66Y17_R_f(R_f_top[421]),
    .Tile_X69Y17_R_t(R_t_top[422]),
    .Tile_X69Y17_R_f(R_f_top[422]),
    .Tile_X72Y17_R_t(R_t_top[423]),
    .Tile_X72Y17_R_f(R_f_top[423]),
    .Tile_X75Y17_R_t(R_t_top[424]),
    .Tile_X75Y17_R_f(R_f_top[424]),
    .Tile_X3Y18_R_t(R_t_top[425]),
    .Tile_X3Y18_R_f(R_f_top[425]),
    .Tile_X6Y18_R_t(R_t_top[426]),
    .Tile_X6Y18_R_f(R_f_top[426]),
    .Tile_X9Y18_R_t(R_t_top[427]),
    .Tile_X9Y18_R_f(R_f_top[427]),
    .Tile_X12Y18_R_t(R_t_top[428]),
    .Tile_X12Y18_R_f(R_f_top[428]),
    .Tile_X15Y18_R_t(R_t_top[429]),
    .Tile_X15Y18_R_f(R_f_top[429]),
    .Tile_X18Y18_R_t(R_t_top[430]),
    .Tile_X18Y18_R_f(R_f_top[430]),
    .Tile_X21Y18_R_t(R_t_top[431]),
    .Tile_X21Y18_R_f(R_f_top[431]),
    .Tile_X24Y18_R_t(R_t_top[432]),
    .Tile_X24Y18_R_f(R_f_top[432]),
    .Tile_X27Y18_R_t(R_t_top[433]),
    .Tile_X27Y18_R_f(R_f_top[433]),
    .Tile_X30Y18_R_t(R_t_top[434]),
    .Tile_X30Y18_R_f(R_f_top[434]),
    .Tile_X33Y18_R_t(R_t_top[435]),
    .Tile_X33Y18_R_f(R_f_top[435]),
    .Tile_X36Y18_R_t(R_t_top[436]),
    .Tile_X36Y18_R_f(R_f_top[436]),
    .Tile_X39Y18_R_t(R_t_top[437]),
    .Tile_X39Y18_R_f(R_f_top[437]),
    .Tile_X42Y18_R_t(R_t_top[438]),
    .Tile_X42Y18_R_f(R_f_top[438]),
    .Tile_X45Y18_R_t(R_t_top[439]),
    .Tile_X45Y18_R_f(R_f_top[439]),
    .Tile_X48Y18_R_t(R_t_top[440]),
    .Tile_X48Y18_R_f(R_f_top[440]),
    .Tile_X51Y18_R_t(R_t_top[441]),
    .Tile_X51Y18_R_f(R_f_top[441]),
    .Tile_X54Y18_R_t(R_t_top[442]),
    .Tile_X54Y18_R_f(R_f_top[442]),
    .Tile_X57Y18_R_t(R_t_top[443]),
    .Tile_X57Y18_R_f(R_f_top[443]),
    .Tile_X60Y18_R_t(R_t_top[444]),
    .Tile_X60Y18_R_f(R_f_top[444]),
    .Tile_X63Y18_R_t(R_t_top[445]),
    .Tile_X63Y18_R_f(R_f_top[445]),
    .Tile_X66Y18_R_t(R_t_top[446]),
    .Tile_X66Y18_R_f(R_f_top[446]),
    .Tile_X69Y18_R_t(R_t_top[447]),
    .Tile_X69Y18_R_f(R_f_top[447]),
    .Tile_X72Y18_R_t(R_t_top[448]),
    .Tile_X72Y18_R_f(R_f_top[448]),
    .Tile_X75Y18_R_t(R_t_top[449]),
    .Tile_X75Y18_R_f(R_f_top[449]),
    .Tile_X3Y19_R_t(R_t_top[450]),
    .Tile_X3Y19_R_f(R_f_top[450]),
    .Tile_X6Y19_R_t(R_t_top[451]),
    .Tile_X6Y19_R_f(R_f_top[451]),
    .Tile_X9Y19_R_t(R_t_top[452]),
    .Tile_X9Y19_R_f(R_f_top[452]),
    .Tile_X12Y19_R_t(R_t_top[453]),
    .Tile_X12Y19_R_f(R_f_top[453]),
    .Tile_X15Y19_R_t(R_t_top[454]),
    .Tile_X15Y19_R_f(R_f_top[454]),
    .Tile_X18Y19_R_t(R_t_top[455]),
    .Tile_X18Y19_R_f(R_f_top[455]),
    .Tile_X21Y19_R_t(R_t_top[456]),
    .Tile_X21Y19_R_f(R_f_top[456]),
    .Tile_X24Y19_R_t(R_t_top[457]),
    .Tile_X24Y19_R_f(R_f_top[457]),
    .Tile_X27Y19_R_t(R_t_top[458]),
    .Tile_X27Y19_R_f(R_f_top[458]),
    .Tile_X30Y19_R_t(R_t_top[459]),
    .Tile_X30Y19_R_f(R_f_top[459]),
    .Tile_X33Y19_R_t(R_t_top[460]),
    .Tile_X33Y19_R_f(R_f_top[460]),
    .Tile_X36Y19_R_t(R_t_top[461]),
    .Tile_X36Y19_R_f(R_f_top[461]),
    .Tile_X39Y19_R_t(R_t_top[462]),
    .Tile_X39Y19_R_f(R_f_top[462]),
    .Tile_X42Y19_R_t(R_t_top[463]),
    .Tile_X42Y19_R_f(R_f_top[463]),
    .Tile_X45Y19_R_t(R_t_top[464]),
    .Tile_X45Y19_R_f(R_f_top[464]),
    .Tile_X48Y19_R_t(R_t_top[465]),
    .Tile_X48Y19_R_f(R_f_top[465]),
    .Tile_X51Y19_R_t(R_t_top[466]),
    .Tile_X51Y19_R_f(R_f_top[466]),
    .Tile_X54Y19_R_t(R_t_top[467]),
    .Tile_X54Y19_R_f(R_f_top[467]),
    .Tile_X57Y19_R_t(R_t_top[468]),
    .Tile_X57Y19_R_f(R_f_top[468]),
    .Tile_X60Y19_R_t(R_t_top[469]),
    .Tile_X60Y19_R_f(R_f_top[469]),
    .Tile_X63Y19_R_t(R_t_top[470]),
    .Tile_X63Y19_R_f(R_f_top[470]),
    .Tile_X66Y19_R_t(R_t_top[471]),
    .Tile_X66Y19_R_f(R_f_top[471]),
    .Tile_X69Y19_R_t(R_t_top[472]),
    .Tile_X69Y19_R_f(R_f_top[472]),
    .Tile_X72Y19_R_t(R_t_top[473]),
    .Tile_X72Y19_R_f(R_f_top[473]),
    .Tile_X75Y19_R_t(R_t_top[474]),
    .Tile_X75Y19_R_f(R_f_top[474]),
    .Tile_X3Y20_R_t(R_t_top[475]),
    .Tile_X3Y20_R_f(R_f_top[475]),
    .Tile_X6Y20_R_t(R_t_top[476]),
    .Tile_X6Y20_R_f(R_f_top[476]),
    .Tile_X9Y20_R_t(R_t_top[477]),
    .Tile_X9Y20_R_f(R_f_top[477]),
    .Tile_X12Y20_R_t(R_t_top[478]),
    .Tile_X12Y20_R_f(R_f_top[478]),
    .Tile_X15Y20_R_t(R_t_top[479]),
    .Tile_X15Y20_R_f(R_f_top[479]),
    .Tile_X18Y20_R_t(R_t_top[480]),
    .Tile_X18Y20_R_f(R_f_top[480]),
    .Tile_X21Y20_R_t(R_t_top[481]),
    .Tile_X21Y20_R_f(R_f_top[481]),
    .Tile_X24Y20_R_t(R_t_top[482]),
    .Tile_X24Y20_R_f(R_f_top[482]),
    .Tile_X27Y20_R_t(R_t_top[483]),
    .Tile_X27Y20_R_f(R_f_top[483]),
    .Tile_X30Y20_R_t(R_t_top[484]),
    .Tile_X30Y20_R_f(R_f_top[484]),
    .Tile_X33Y20_R_t(R_t_top[485]),
    .Tile_X33Y20_R_f(R_f_top[485]),
    .Tile_X36Y20_R_t(R_t_top[486]),
    .Tile_X36Y20_R_f(R_f_top[486]),
    .Tile_X39Y20_R_t(R_t_top[487]),
    .Tile_X39Y20_R_f(R_f_top[487]),
    .Tile_X42Y20_R_t(R_t_top[488]),
    .Tile_X42Y20_R_f(R_f_top[488]),
    .Tile_X45Y20_R_t(R_t_top[489]),
    .Tile_X45Y20_R_f(R_f_top[489]),
    .Tile_X48Y20_R_t(R_t_top[490]),
    .Tile_X48Y20_R_f(R_f_top[490]),
    .Tile_X51Y20_R_t(R_t_top[491]),
    .Tile_X51Y20_R_f(R_f_top[491]),
    .Tile_X54Y20_R_t(R_t_top[492]),
    .Tile_X54Y20_R_f(R_f_top[492]),
    .Tile_X57Y20_R_t(R_t_top[493]),
    .Tile_X57Y20_R_f(R_f_top[493]),
    .Tile_X60Y20_R_t(R_t_top[494]),
    .Tile_X60Y20_R_f(R_f_top[494]),
    .Tile_X63Y20_R_t(R_t_top[495]),
    .Tile_X63Y20_R_f(R_f_top[495]),
    .Tile_X66Y20_R_t(R_t_top[496]),
    .Tile_X66Y20_R_f(R_f_top[496]),
    .Tile_X69Y20_R_t(R_t_top[497]),
    .Tile_X69Y20_R_f(R_f_top[497]),
    .Tile_X72Y20_R_t(R_t_top[498]),
    .Tile_X72Y20_R_f(R_f_top[498]),
    .Tile_X75Y20_R_t(R_t_top[499]),
    .Tile_X75Y20_R_f(R_f_top[499]),
    .Tile_X3Y21_R_t(R_t_top[500]),
    .Tile_X3Y21_R_f(R_f_top[500]),
    .Tile_X6Y21_R_t(R_t_top[501]),
    .Tile_X6Y21_R_f(R_f_top[501]),
    .Tile_X9Y21_R_t(R_t_top[502]),
    .Tile_X9Y21_R_f(R_f_top[502]),
    .Tile_X12Y21_R_t(R_t_top[503]),
    .Tile_X12Y21_R_f(R_f_top[503]),
    .Tile_X15Y21_R_t(R_t_top[504]),
    .Tile_X15Y21_R_f(R_f_top[504]),
    .Tile_X18Y21_R_t(R_t_top[505]),
    .Tile_X18Y21_R_f(R_f_top[505]),
    .Tile_X21Y21_R_t(R_t_top[506]),
    .Tile_X21Y21_R_f(R_f_top[506]),
    .Tile_X24Y21_R_t(R_t_top[507]),
    .Tile_X24Y21_R_f(R_f_top[507]),
    .Tile_X27Y21_R_t(R_t_top[508]),
    .Tile_X27Y21_R_f(R_f_top[508]),
    .Tile_X30Y21_R_t(R_t_top[509]),
    .Tile_X30Y21_R_f(R_f_top[509]),
    .Tile_X33Y21_R_t(R_t_top[510]),
    .Tile_X33Y21_R_f(R_f_top[510]),
    .Tile_X36Y21_R_t(R_t_top[511]),
    .Tile_X36Y21_R_f(R_f_top[511]),
    .Tile_X39Y21_R_t(R_t_top[512]),
    .Tile_X39Y21_R_f(R_f_top[512]),
    .Tile_X42Y21_R_t(R_t_top[513]),
    .Tile_X42Y21_R_f(R_f_top[513]),
    .Tile_X45Y21_R_t(R_t_top[514]),
    .Tile_X45Y21_R_f(R_f_top[514]),
    .Tile_X48Y21_R_t(R_t_top[515]),
    .Tile_X48Y21_R_f(R_f_top[515]),
    .Tile_X51Y21_R_t(R_t_top[516]),
    .Tile_X51Y21_R_f(R_f_top[516]),
    .Tile_X54Y21_R_t(R_t_top[517]),
    .Tile_X54Y21_R_f(R_f_top[517]),
    .Tile_X57Y21_R_t(R_t_top[518]),
    .Tile_X57Y21_R_f(R_f_top[518]),
    .Tile_X60Y21_R_t(R_t_top[519]),
    .Tile_X60Y21_R_f(R_f_top[519]),
    .Tile_X63Y21_R_t(R_t_top[520]),
    .Tile_X63Y21_R_f(R_f_top[520]),
    .Tile_X66Y21_R_t(R_t_top[521]),
    .Tile_X66Y21_R_f(R_f_top[521]),
    .Tile_X69Y21_R_t(R_t_top[522]),
    .Tile_X69Y21_R_f(R_f_top[522]),
    .Tile_X72Y21_R_t(R_t_top[523]),
    .Tile_X72Y21_R_f(R_f_top[523]),
    .Tile_X75Y21_R_t(R_t_top[524]),
    .Tile_X75Y21_R_f(R_f_top[524]),
    .Tile_X3Y22_R_t(R_t_top[525]),
    .Tile_X3Y22_R_f(R_f_top[525]),
    .Tile_X6Y22_R_t(R_t_top[526]),
    .Tile_X6Y22_R_f(R_f_top[526]),
    .Tile_X9Y22_R_t(R_t_top[527]),
    .Tile_X9Y22_R_f(R_f_top[527]),
    .Tile_X12Y22_R_t(R_t_top[528]),
    .Tile_X12Y22_R_f(R_f_top[528]),
    .Tile_X15Y22_R_t(R_t_top[529]),
    .Tile_X15Y22_R_f(R_f_top[529]),
    .Tile_X18Y22_R_t(R_t_top[530]),
    .Tile_X18Y22_R_f(R_f_top[530]),
    .Tile_X21Y22_R_t(R_t_top[531]),
    .Tile_X21Y22_R_f(R_f_top[531]),
    .Tile_X24Y22_R_t(R_t_top[532]),
    .Tile_X24Y22_R_f(R_f_top[532]),
    .Tile_X27Y22_R_t(R_t_top[533]),
    .Tile_X27Y22_R_f(R_f_top[533]),
    .Tile_X30Y22_R_t(R_t_top[534]),
    .Tile_X30Y22_R_f(R_f_top[534]),
    .Tile_X33Y22_R_t(R_t_top[535]),
    .Tile_X33Y22_R_f(R_f_top[535]),
    .Tile_X36Y22_R_t(R_t_top[536]),
    .Tile_X36Y22_R_f(R_f_top[536]),
    .Tile_X39Y22_R_t(R_t_top[537]),
    .Tile_X39Y22_R_f(R_f_top[537]),
    .Tile_X42Y22_R_t(R_t_top[538]),
    .Tile_X42Y22_R_f(R_f_top[538]),
    .Tile_X45Y22_R_t(R_t_top[539]),
    .Tile_X45Y22_R_f(R_f_top[539]),
    .Tile_X48Y22_R_t(R_t_top[540]),
    .Tile_X48Y22_R_f(R_f_top[540]),
    .Tile_X51Y22_R_t(R_t_top[541]),
    .Tile_X51Y22_R_f(R_f_top[541]),
    .Tile_X54Y22_R_t(R_t_top[542]),
    .Tile_X54Y22_R_f(R_f_top[542]),
    .Tile_X57Y22_R_t(R_t_top[543]),
    .Tile_X57Y22_R_f(R_f_top[543]),
    .Tile_X60Y22_R_t(R_t_top[544]),
    .Tile_X60Y22_R_f(R_f_top[544]),
    .Tile_X63Y22_R_t(R_t_top[545]),
    .Tile_X63Y22_R_f(R_f_top[545]),
    .Tile_X66Y22_R_t(R_t_top[546]),
    .Tile_X66Y22_R_f(R_f_top[546]),
    .Tile_X69Y22_R_t(R_t_top[547]),
    .Tile_X69Y22_R_f(R_f_top[547]),
    .Tile_X72Y22_R_t(R_t_top[548]),
    .Tile_X72Y22_R_f(R_f_top[548]),
    .Tile_X75Y22_R_t(R_t_top[549]),
    .Tile_X75Y22_R_f(R_f_top[549]),
    .Tile_X3Y23_R_t(R_t_top[550]),
    .Tile_X3Y23_R_f(R_f_top[550]),
    .Tile_X6Y23_R_t(R_t_top[551]),
    .Tile_X6Y23_R_f(R_f_top[551]),
    .Tile_X9Y23_R_t(R_t_top[552]),
    .Tile_X9Y23_R_f(R_f_top[552]),
    .Tile_X12Y23_R_t(R_t_top[553]),
    .Tile_X12Y23_R_f(R_f_top[553]),
    .Tile_X15Y23_R_t(R_t_top[554]),
    .Tile_X15Y23_R_f(R_f_top[554]),
    .Tile_X18Y23_R_t(R_t_top[555]),
    .Tile_X18Y23_R_f(R_f_top[555]),
    .Tile_X21Y23_R_t(R_t_top[556]),
    .Tile_X21Y23_R_f(R_f_top[556]),
    .Tile_X24Y23_R_t(R_t_top[557]),
    .Tile_X24Y23_R_f(R_f_top[557]),
    .Tile_X27Y23_R_t(R_t_top[558]),
    .Tile_X27Y23_R_f(R_f_top[558]),
    .Tile_X30Y23_R_t(R_t_top[559]),
    .Tile_X30Y23_R_f(R_f_top[559]),
    .Tile_X33Y23_R_t(R_t_top[560]),
    .Tile_X33Y23_R_f(R_f_top[560]),
    .Tile_X36Y23_R_t(R_t_top[561]),
    .Tile_X36Y23_R_f(R_f_top[561]),
    .Tile_X39Y23_R_t(R_t_top[562]),
    .Tile_X39Y23_R_f(R_f_top[562]),
    .Tile_X42Y23_R_t(R_t_top[563]),
    .Tile_X42Y23_R_f(R_f_top[563]),
    .Tile_X45Y23_R_t(R_t_top[564]),
    .Tile_X45Y23_R_f(R_f_top[564]),
    .Tile_X48Y23_R_t(R_t_top[565]),
    .Tile_X48Y23_R_f(R_f_top[565]),
    .Tile_X51Y23_R_t(R_t_top[566]),
    .Tile_X51Y23_R_f(R_f_top[566]),
    .Tile_X54Y23_R_t(R_t_top[567]),
    .Tile_X54Y23_R_f(R_f_top[567]),
    .Tile_X57Y23_R_t(R_t_top[568]),
    .Tile_X57Y23_R_f(R_f_top[568]),
    .Tile_X60Y23_R_t(R_t_top[569]),
    .Tile_X60Y23_R_f(R_f_top[569]),
    .Tile_X63Y23_R_t(R_t_top[570]),
    .Tile_X63Y23_R_f(R_f_top[570]),
    .Tile_X66Y23_R_t(R_t_top[571]),
    .Tile_X66Y23_R_f(R_f_top[571]),
    .Tile_X69Y23_R_t(R_t_top[572]),
    .Tile_X69Y23_R_f(R_f_top[572]),
    .Tile_X72Y23_R_t(R_t_top[573]),
    .Tile_X72Y23_R_f(R_f_top[573]),
    .Tile_X75Y23_R_t(R_t_top[574]),
    .Tile_X75Y23_R_f(R_f_top[574]),
    .Tile_X0Y1_A_F_masked1(F_masked1_top[0]),
    .Tile_X0Y1_A_F_masked2(F_masked2_top[0]),
    .Tile_X0Y2_A_F_masked1(F_masked1_top[1]),
    .Tile_X0Y2_A_F_masked2(F_masked2_top[1]),
    .Tile_X0Y3_A_F_masked1(F_masked1_top[2]),
    .Tile_X0Y3_A_F_masked2(F_masked2_top[2]),
    .Tile_X0Y4_A_F_masked1(F_masked1_top[3]),
    .Tile_X0Y4_A_F_masked2(F_masked2_top[3]),
    .Tile_X0Y5_A_F_masked1(F_masked1_top[4]),
    .Tile_X0Y5_A_F_masked2(F_masked2_top[4]),
    .Tile_X0Y6_A_F_masked1(F_masked1_top[5]),
    .Tile_X0Y6_A_F_masked2(F_masked2_top[5]),
    .Tile_X0Y7_A_F_masked1(F_masked1_top[6]),
    .Tile_X0Y7_A_F_masked2(F_masked2_top[6]),
    .Tile_X0Y8_A_F_masked1(F_masked1_top[7]),
    .Tile_X0Y8_A_F_masked2(F_masked2_top[7]),
    .Tile_X0Y9_A_F_masked1(F_masked1_top[8]),
    .Tile_X0Y9_A_F_masked2(F_masked2_top[8]),
    .Tile_X0Y10_A_F_masked1(F_masked1_top[9]),
    .Tile_X0Y10_A_F_masked2(F_masked2_top[9]),
    .Tile_X0Y11_A_F_masked1(F_masked1_top[10]),
    .Tile_X0Y11_A_F_masked2(F_masked2_top[10]),
    .Tile_X0Y12_A_F_masked1(F_masked1_top[11]),
    .Tile_X0Y12_A_F_masked2(F_masked2_top[11]),
    .Tile_X0Y13_A_F_masked1(F_masked1_top[12]),
    .Tile_X0Y13_A_F_masked2(F_masked2_top[12]),
    .Tile_X0Y14_A_F_masked1(F_masked1_top[13]),
    .Tile_X0Y14_A_F_masked2(F_masked2_top[13]),
    .Tile_X0Y15_A_F_masked1(F_masked1_top[14]),
    .Tile_X0Y15_A_F_masked2(F_masked2_top[14]),
    .Tile_X0Y16_A_F_masked1(F_masked1_top[15]),
    .Tile_X0Y16_A_F_masked2(F_masked2_top[15]),
    .Tile_X0Y17_A_F_masked1(F_masked1_top[16]),
    .Tile_X0Y17_A_F_masked2(F_masked2_top[16]),
    .Tile_X0Y18_A_F_masked1(F_masked1_top[17]),
    .Tile_X0Y18_A_F_masked2(F_masked2_top[17]),
    .Tile_X0Y19_A_F_masked1(F_masked1_top[18]),
    .Tile_X0Y19_A_F_masked2(F_masked2_top[18]),
    .Tile_X0Y20_A_F_masked1(F_masked1_top[19]),
    .Tile_X0Y20_A_F_masked2(F_masked2_top[19]),
    .Tile_X0Y21_A_F_masked1(F_masked1_top[20]),
    .Tile_X0Y21_A_F_masked2(F_masked2_top[20]),
    .Tile_X0Y22_A_F_masked1(F_masked1_top[21]),
    .Tile_X0Y22_A_F_masked2(F_masked2_top[21]),
    .Tile_X0Y23_A_F_masked1(F_masked1_top[22]),
    .Tile_X0Y23_A_F_masked2(F_masked2_top[22]),
    .Tile_X10Y1_A_F_ctrl(F_ctrl_top[0]),
    .Tile_X10Y2_A_F_ctrl(F_ctrl_top[1]),
    .Tile_X10Y3_A_F_ctrl(F_ctrl_top[2]),
    .Tile_X10Y4_A_F_ctrl(F_ctrl_top[3]),
    .Tile_X10Y5_A_F_ctrl(F_ctrl_top[4]),
    .Tile_X10Y6_A_F_ctrl(F_ctrl_top[5]),
    .Tile_X10Y7_A_F_ctrl(F_ctrl_top[6]),
    .Tile_X10Y8_A_F_ctrl(F_ctrl_top[7]),
    .Tile_X10Y9_A_F_ctrl(F_ctrl_top[8]),
    .Tile_X10Y10_A_F_ctrl(F_ctrl_top[9]),
    .Tile_X10Y11_A_F_ctrl(F_ctrl_top[10]),
    .Tile_X10Y12_A_F_ctrl(F_ctrl_top[11]),
    .Tile_X10Y13_A_F_ctrl(F_ctrl_top[12]),
    .Tile_X10Y14_A_F_ctrl(F_ctrl_top[13]),
    .Tile_X10Y15_A_F_ctrl(F_ctrl_top[14]),
    .Tile_X10Y16_A_F_ctrl(F_ctrl_top[15]),
    .Tile_X10Y17_A_F_ctrl(F_ctrl_top[16]),
    .Tile_X10Y18_A_F_ctrl(F_ctrl_top[17]),
    .Tile_X10Y19_A_F_ctrl(F_ctrl_top[18]),
    .Tile_X10Y20_A_F_ctrl(F_ctrl_top[19]),
    .Tile_X10Y21_A_F_ctrl(F_ctrl_top[20]),
    .Tile_X10Y22_A_F_ctrl(F_ctrl_top[21]),
    .Tile_X10Y23_A_F_ctrl(F_ctrl_top[22]),
    .Tile_X0Y1_A_prech1(prech1),
    .Tile_X0Y1_A_prech2(prech2),
    .Tile_X10Y1_A_prech2(prech2),
    .Tile_X0Y2_A_prech1(prech1),
    .Tile_X0Y2_A_prech2(prech2),
    .Tile_X10Y2_A_prech2(prech2),
    .Tile_X0Y3_A_prech1(prech1),
    .Tile_X0Y3_A_prech2(prech2),
    .Tile_X10Y3_A_prech2(prech2),
    .Tile_X0Y4_A_prech1(prech1),
    .Tile_X0Y4_A_prech2(prech2),
    .Tile_X10Y4_A_prech2(prech2),
    .Tile_X0Y5_A_prech1(prech1),
    .Tile_X0Y5_A_prech2(prech2),
    .Tile_X10Y5_A_prech2(prech2),
    .Tile_X0Y6_A_prech1(prech1),
    .Tile_X0Y6_A_prech2(prech2),
    .Tile_X10Y6_A_prech2(prech2),
    .Tile_X0Y7_A_prech1(prech1),
    .Tile_X0Y7_A_prech2(prech2),
    .Tile_X10Y7_A_prech2(prech2),
    .Tile_X0Y8_A_prech1(prech1),
    .Tile_X0Y8_A_prech2(prech2),
    .Tile_X10Y8_A_prech2(prech2),
    .Tile_X0Y9_A_prech1(prech1),
    .Tile_X0Y9_A_prech2(prech2),
    .Tile_X10Y9_A_prech2(prech2),
    .Tile_X0Y10_A_prech1(prech1),
    .Tile_X0Y10_A_prech2(prech2),
    .Tile_X10Y10_A_prech2(prech2),
    .Tile_X0Y11_A_prech1(prech1),
    .Tile_X0Y11_A_prech2(prech2),
    .Tile_X10Y11_A_prech2(prech2),
    .Tile_X0Y12_A_prech1(prech1),
    .Tile_X0Y12_A_prech2(prech2),
    .Tile_X10Y12_A_prech2(prech2),
    .Tile_X0Y13_A_prech1(prech1),
    .Tile_X0Y13_A_prech2(prech2),
    .Tile_X10Y13_A_prech2(prech2),
    .Tile_X0Y14_A_prech1(prech1),
    .Tile_X0Y14_A_prech2(prech2),
    .Tile_X10Y14_A_prech2(prech2),
    .Tile_X0Y15_A_prech1(prech1),
    .Tile_X0Y15_A_prech2(prech2),
    .Tile_X10Y15_A_prech2(prech2),
    .Tile_X0Y16_A_prech1(prech1),
    .Tile_X0Y16_A_prech2(prech2),
    .Tile_X10Y16_A_prech2(prech2),
    .Tile_X0Y17_A_prech1(prech1),
    .Tile_X0Y17_A_prech2(prech2),
    .Tile_X10Y17_A_prech2(prech2),
    .Tile_X0Y18_A_prech1(prech1),
    .Tile_X0Y18_A_prech2(prech2),
    .Tile_X10Y18_A_prech2(prech2),
    .Tile_X0Y19_A_prech1(prech1),
    .Tile_X0Y19_A_prech2(prech2),
    .Tile_X10Y19_A_prech2(prech2),
    .Tile_X0Y20_A_prech1(prech1),
    .Tile_X0Y20_A_prech2(prech2),
    .Tile_X10Y20_A_prech2(prech2),
    .Tile_X0Y21_A_prech1(prech1),
    .Tile_X0Y21_A_prech2(prech2),
    .Tile_X10Y21_A_prech2(prech2),
    .Tile_X0Y22_A_prech1(prech1),
    .Tile_X0Y22_A_prech2(prech2),
    .Tile_X10Y22_A_prech2(prech2),
    .Tile_X0Y23_A_prech1(prech1),
    .Tile_X0Y23_A_prech2(prech2),
    .Tile_X10Y23_A_prech2(prech2),
    .Tile_X0Y1_A_I_top_0_t(I_top_0_t[0]),
    .Tile_X0Y1_A_I_top_0_f(I_top_0_f[0]),
    .Tile_X0Y1_A_I_top_1_t(I_top_1_t[0]),
    .Tile_X0Y1_A_I_top_1_f(I_top_1_f[0]),
    .Tile_X0Y2_A_I_top_0_t(I_top_0_t[1]),
    .Tile_X0Y2_A_I_top_0_f(I_top_0_f[1]),
    .Tile_X0Y2_A_I_top_1_t(I_top_1_t[1]),
    .Tile_X0Y2_A_I_top_1_f(I_top_1_f[1]),
    .Tile_X0Y3_A_I_top_0_t(I_top_0_t[2]),
    .Tile_X0Y3_A_I_top_0_f(I_top_0_f[2]),
    .Tile_X0Y3_A_I_top_1_t(I_top_1_t[2]),
    .Tile_X0Y3_A_I_top_1_f(I_top_1_f[2]),
    .Tile_X0Y4_A_I_top_0_t(I_top_0_t[3]),
    .Tile_X0Y4_A_I_top_0_f(I_top_0_f[3]),
    .Tile_X0Y4_A_I_top_1_t(I_top_1_t[3]),
    .Tile_X0Y4_A_I_top_1_f(I_top_1_f[3]),
    .Tile_X0Y5_A_I_top_0_t(I_top_0_t[4]),
    .Tile_X0Y5_A_I_top_0_f(I_top_0_f[4]),
    .Tile_X0Y5_A_I_top_1_t(I_top_1_t[4]),
    .Tile_X0Y5_A_I_top_1_f(I_top_1_f[4]),
    .Tile_X0Y6_A_I_top_0_t(I_top_0_t[5]),
    .Tile_X0Y6_A_I_top_0_f(I_top_0_f[5]),
    .Tile_X0Y6_A_I_top_1_t(I_top_1_t[5]),
    .Tile_X0Y6_A_I_top_1_f(I_top_1_f[5]),
    .Tile_X0Y7_A_I_top_0_t(I_top_0_t[6]),
    .Tile_X0Y7_A_I_top_0_f(I_top_0_f[6]),
    .Tile_X0Y7_A_I_top_1_t(I_top_1_t[6]),
    .Tile_X0Y7_A_I_top_1_f(I_top_1_f[6]),
    .Tile_X0Y8_A_I_top_0_t(I_top_0_t[7]),
    .Tile_X0Y8_A_I_top_0_f(I_top_0_f[7]),
    .Tile_X0Y8_A_I_top_1_t(I_top_1_t[7]),
    .Tile_X0Y8_A_I_top_1_f(I_top_1_f[7]),
    .Tile_X0Y9_A_I_top_0_t(I_top_0_t[8]),
    .Tile_X0Y9_A_I_top_0_f(I_top_0_f[8]),
    .Tile_X0Y9_A_I_top_1_t(I_top_1_t[8]),
    .Tile_X0Y9_A_I_top_1_f(I_top_1_f[8]),
    .Tile_X0Y10_A_I_top_0_t(I_top_0_t[9]),
    .Tile_X0Y10_A_I_top_0_f(I_top_0_f[9]),
    .Tile_X0Y10_A_I_top_1_t(I_top_1_t[9]),
    .Tile_X0Y10_A_I_top_1_f(I_top_1_f[9]),
    .Tile_X0Y11_A_I_top_0_t(I_top_0_t[10]),
    .Tile_X0Y11_A_I_top_0_f(I_top_0_f[10]),
    .Tile_X0Y11_A_I_top_1_t(I_top_1_t[10]),
    .Tile_X0Y11_A_I_top_1_f(I_top_1_f[10]),
    .Tile_X0Y12_A_I_top_0_t(I_top_0_t[11]),
    .Tile_X0Y12_A_I_top_0_f(I_top_0_f[11]),
    .Tile_X0Y12_A_I_top_1_t(I_top_1_t[11]),
    .Tile_X0Y12_A_I_top_1_f(I_top_1_f[11]),
    .Tile_X0Y13_A_I_top_0_t(I_top_0_t[12]),
    .Tile_X0Y13_A_I_top_0_f(I_top_0_f[12]),
    .Tile_X0Y13_A_I_top_1_t(I_top_1_t[12]),
    .Tile_X0Y13_A_I_top_1_f(I_top_1_f[12]),
    .Tile_X0Y14_A_I_top_0_t(I_top_0_t[13]),
    .Tile_X0Y14_A_I_top_0_f(I_top_0_f[13]),
    .Tile_X0Y14_A_I_top_1_t(I_top_1_t[13]),
    .Tile_X0Y14_A_I_top_1_f(I_top_1_f[13]),
    .Tile_X0Y15_A_I_top_0_t(I_top_0_t[14]),
    .Tile_X0Y15_A_I_top_0_f(I_top_0_f[14]),
    .Tile_X0Y15_A_I_top_1_t(I_top_1_t[14]),
    .Tile_X0Y15_A_I_top_1_f(I_top_1_f[14]),
    .Tile_X0Y16_A_I_top_0_t(I_top_0_t[15]),
    .Tile_X0Y16_A_I_top_0_f(I_top_0_f[15]),
    .Tile_X0Y16_A_I_top_1_t(I_top_1_t[15]),
    .Tile_X0Y16_A_I_top_1_f(I_top_1_f[15]),
    .Tile_X0Y17_A_I_top_0_t(I_top_0_t[16]),
    .Tile_X0Y17_A_I_top_0_f(I_top_0_f[16]),
    .Tile_X0Y17_A_I_top_1_t(I_top_1_t[16]),
    .Tile_X0Y17_A_I_top_1_f(I_top_1_f[16]),
    .Tile_X0Y18_A_I_top_0_t(I_top_0_t[17]),
    .Tile_X0Y18_A_I_top_0_f(I_top_0_f[17]),
    .Tile_X0Y18_A_I_top_1_t(I_top_1_t[17]),
    .Tile_X0Y18_A_I_top_1_f(I_top_1_f[17]),
    .Tile_X0Y19_A_I_top_0_t(I_top_0_t[18]),
    .Tile_X0Y19_A_I_top_0_f(I_top_0_f[18]),
    .Tile_X0Y19_A_I_top_1_t(I_top_1_t[18]),
    .Tile_X0Y19_A_I_top_1_f(I_top_1_f[18]),
    .Tile_X0Y20_A_I_top_0_t(I_top_0_t[19]),
    .Tile_X0Y20_A_I_top_0_f(I_top_0_f[19]),
    .Tile_X0Y20_A_I_top_1_t(I_top_1_t[19]),
    .Tile_X0Y20_A_I_top_1_f(I_top_1_f[19]),
    .Tile_X0Y21_A_I_top_0_t(I_top_0_t[20]),
    .Tile_X0Y21_A_I_top_0_f(I_top_0_f[20]),
    .Tile_X0Y21_A_I_top_1_t(I_top_1_t[20]),
    .Tile_X0Y21_A_I_top_1_f(I_top_1_f[20]),
    .Tile_X0Y22_A_I_top_0_t(I_top_0_t[21]),
    .Tile_X0Y22_A_I_top_0_f(I_top_0_f[21]),
    .Tile_X0Y22_A_I_top_1_t(I_top_1_t[21]),
    .Tile_X0Y22_A_I_top_1_f(I_top_1_f[21]),
    .Tile_X0Y23_A_I_top_0_t(I_top_0_t[22]),
    .Tile_X0Y23_A_I_top_0_f(I_top_0_f[22]),
    .Tile_X0Y23_A_I_top_1_t(I_top_1_t[22]),
    .Tile_X0Y23_A_I_top_1_f(I_top_1_f[22]),
    .Tile_X0Y1_A_T_top(T_top[0]),
    .Tile_X0Y2_A_T_top(T_top[1]),
    .Tile_X0Y3_A_T_top(T_top[2]),
    .Tile_X0Y4_A_T_top(T_top[3]),
    .Tile_X0Y5_A_T_top(T_top[4]),
    .Tile_X0Y6_A_T_top(T_top[5]),
    .Tile_X0Y7_A_T_top(T_top[6]),
    .Tile_X0Y8_A_T_top(T_top[7]),
    .Tile_X0Y9_A_T_top(T_top[8]),
    .Tile_X0Y10_A_T_top(T_top[9]),
    .Tile_X0Y11_A_T_top(T_top[10]),
    .Tile_X0Y12_A_T_top(T_top[11]),
    .Tile_X0Y13_A_T_top(T_top[12]),
    .Tile_X0Y14_A_T_top(T_top[13]),
    .Tile_X0Y15_A_T_top(T_top[14]),
    .Tile_X0Y16_A_T_top(T_top[15]),
    .Tile_X0Y17_A_T_top(T_top[16]),
    .Tile_X0Y18_A_T_top(T_top[17]),
    .Tile_X0Y19_A_T_top(T_top[18]),
    .Tile_X0Y20_A_T_top(T_top[19]),
    .Tile_X0Y21_A_T_top(T_top[20]),
    .Tile_X0Y22_A_T_top(T_top[21]),
    .Tile_X0Y23_A_T_top(T_top[22]),
    .Tile_X0Y1_A_O_top_0_t(O_top_0_t[0]),
    .Tile_X0Y1_A_O_top_0_f(O_top_0_f[0]),
    .Tile_X0Y1_A_O_top_1_t(O_top_1_t[0]),
    .Tile_X0Y1_A_O_top_1_f(O_top_1_f[0]),
    .Tile_X0Y2_A_O_top_0_t(O_top_0_t[1]),
    .Tile_X0Y2_A_O_top_0_f(O_top_0_f[1]),
    .Tile_X0Y2_A_O_top_1_t(O_top_1_t[1]),
    .Tile_X0Y2_A_O_top_1_f(O_top_1_f[1]),
    .Tile_X0Y3_A_O_top_0_t(O_top_0_t[2]),
    .Tile_X0Y3_A_O_top_0_f(O_top_0_f[2]),
    .Tile_X0Y3_A_O_top_1_t(O_top_1_t[2]),
    .Tile_X0Y3_A_O_top_1_f(O_top_1_f[2]),
    .Tile_X0Y4_A_O_top_0_t(O_top_0_t[3]),
    .Tile_X0Y4_A_O_top_0_f(O_top_0_f[3]),
    .Tile_X0Y4_A_O_top_1_t(O_top_1_t[3]),
    .Tile_X0Y4_A_O_top_1_f(O_top_1_f[3]),
    .Tile_X0Y5_A_O_top_0_t(O_top_0_t[4]),
    .Tile_X0Y5_A_O_top_0_f(O_top_0_f[4]),
    .Tile_X0Y5_A_O_top_1_t(O_top_1_t[4]),
    .Tile_X0Y5_A_O_top_1_f(O_top_1_f[4]),
    .Tile_X0Y6_A_O_top_0_t(O_top_0_t[5]),
    .Tile_X0Y6_A_O_top_0_f(O_top_0_f[5]),
    .Tile_X0Y6_A_O_top_1_t(O_top_1_t[5]),
    .Tile_X0Y6_A_O_top_1_f(O_top_1_f[5]),
    .Tile_X0Y7_A_O_top_0_t(O_top_0_t[6]),
    .Tile_X0Y7_A_O_top_0_f(O_top_0_f[6]),
    .Tile_X0Y7_A_O_top_1_t(O_top_1_t[6]),
    .Tile_X0Y7_A_O_top_1_f(O_top_1_f[6]),
    .Tile_X0Y8_A_O_top_0_t(O_top_0_t[7]),
    .Tile_X0Y8_A_O_top_0_f(O_top_0_f[7]),
    .Tile_X0Y8_A_O_top_1_t(O_top_1_t[7]),
    .Tile_X0Y8_A_O_top_1_f(O_top_1_f[7]),
    .Tile_X0Y9_A_O_top_0_t(O_top_0_t[8]),
    .Tile_X0Y9_A_O_top_0_f(O_top_0_f[8]),
    .Tile_X0Y9_A_O_top_1_t(O_top_1_t[8]),
    .Tile_X0Y9_A_O_top_1_f(O_top_1_f[8]),
    .Tile_X0Y10_A_O_top_0_t(O_top_0_t[9]),
    .Tile_X0Y10_A_O_top_0_f(O_top_0_f[9]),
    .Tile_X0Y10_A_O_top_1_t(O_top_1_t[9]),
    .Tile_X0Y10_A_O_top_1_f(O_top_1_f[9]),
    .Tile_X0Y11_A_O_top_0_t(O_top_0_t[10]),
    .Tile_X0Y11_A_O_top_0_f(O_top_0_f[10]),
    .Tile_X0Y11_A_O_top_1_t(O_top_1_t[10]),
    .Tile_X0Y11_A_O_top_1_f(O_top_1_f[10]),
    .Tile_X0Y12_A_O_top_0_t(O_top_0_t[11]),
    .Tile_X0Y12_A_O_top_0_f(O_top_0_f[11]),
    .Tile_X0Y12_A_O_top_1_t(O_top_1_t[11]),
    .Tile_X0Y12_A_O_top_1_f(O_top_1_f[11]),
    .Tile_X0Y13_A_O_top_0_t(O_top_0_t[12]),
    .Tile_X0Y13_A_O_top_0_f(O_top_0_f[12]),
    .Tile_X0Y13_A_O_top_1_t(O_top_1_t[12]),
    .Tile_X0Y13_A_O_top_1_f(O_top_1_f[12]),
    .Tile_X0Y14_A_O_top_0_t(O_top_0_t[13]),
    .Tile_X0Y14_A_O_top_0_f(O_top_0_f[13]),
    .Tile_X0Y14_A_O_top_1_t(O_top_1_t[13]),
    .Tile_X0Y14_A_O_top_1_f(O_top_1_f[13]),
    .Tile_X0Y15_A_O_top_0_t(O_top_0_t[14]),
    .Tile_X0Y15_A_O_top_0_f(O_top_0_f[14]),
    .Tile_X0Y15_A_O_top_1_t(O_top_1_t[14]),
    .Tile_X0Y15_A_O_top_1_f(O_top_1_f[14]),
    .Tile_X0Y16_A_O_top_0_t(O_top_0_t[15]),
    .Tile_X0Y16_A_O_top_0_f(O_top_0_f[15]),
    .Tile_X0Y16_A_O_top_1_t(O_top_1_t[15]),
    .Tile_X0Y16_A_O_top_1_f(O_top_1_f[15]),
    .Tile_X0Y17_A_O_top_0_t(O_top_0_t[16]),
    .Tile_X0Y17_A_O_top_0_f(O_top_0_f[16]),
    .Tile_X0Y17_A_O_top_1_t(O_top_1_t[16]),
    .Tile_X0Y17_A_O_top_1_f(O_top_1_f[16]),
    .Tile_X0Y18_A_O_top_0_t(O_top_0_t[17]),
    .Tile_X0Y18_A_O_top_0_f(O_top_0_f[17]),
    .Tile_X0Y18_A_O_top_1_t(O_top_1_t[17]),
    .Tile_X0Y18_A_O_top_1_f(O_top_1_f[17]),
    .Tile_X0Y19_A_O_top_0_t(O_top_0_t[18]),
    .Tile_X0Y19_A_O_top_0_f(O_top_0_f[18]),
    .Tile_X0Y19_A_O_top_1_t(O_top_1_t[18]),
    .Tile_X0Y19_A_O_top_1_f(O_top_1_f[18]),
    .Tile_X0Y20_A_O_top_0_t(O_top_0_t[19]),
    .Tile_X0Y20_A_O_top_0_f(O_top_0_f[19]),
    .Tile_X0Y20_A_O_top_1_t(O_top_1_t[19]),
    .Tile_X0Y20_A_O_top_1_f(O_top_1_f[19]),
    .Tile_X0Y21_A_O_top_0_t(O_top_0_t[20]),
    .Tile_X0Y21_A_O_top_0_f(O_top_0_f[20]),
    .Tile_X0Y21_A_O_top_1_t(O_top_1_t[20]),
    .Tile_X0Y21_A_O_top_1_f(O_top_1_f[20]),
    .Tile_X0Y22_A_O_top_0_t(O_top_0_t[21]),
    .Tile_X0Y22_A_O_top_0_f(O_top_0_f[21]),
    .Tile_X0Y22_A_O_top_1_t(O_top_1_t[21]),
    .Tile_X0Y22_A_O_top_1_f(O_top_1_f[21]),
    .Tile_X0Y23_A_O_top_0_t(O_top_0_t[22]),
    .Tile_X0Y23_A_O_top_0_f(O_top_0_f[22]),
    .Tile_X0Y23_A_O_top_1_t(O_top_1_t[22]),
    .Tile_X0Y23_A_O_top_1_f(O_top_1_f[22]),
    .Tile_X10Y1_A_I_top_0_t(ctrl_I_top_0_t[0]),
    .Tile_X10Y1_A_I_top_0_f(ctrl_I_top_0_f[0]),
    .Tile_X10Y1_A_T_top(ctrl_T_top[0]),
    .Tile_X10Y1_A_O_top_0_t(ctrl_O_top_0_t[0]),
    .Tile_X10Y1_A_O_top_0_f(ctrl_O_top_0_f[0]),
    .Tile_X10Y2_A_I_top_0_t(ctrl_I_top_0_t[1]),
    .Tile_X10Y2_A_I_top_0_f(ctrl_I_top_0_f[1]),
    .Tile_X10Y2_A_T_top(ctrl_T_top[1]),
    .Tile_X10Y2_A_O_top_0_t(ctrl_O_top_0_t[1]),
    .Tile_X10Y2_A_O_top_0_f(ctrl_O_top_0_f[1]),
    .Tile_X10Y3_A_I_top_0_t(ctrl_I_top_0_t[2]),
    .Tile_X10Y3_A_I_top_0_f(ctrl_I_top_0_f[2]),
    .Tile_X10Y3_A_T_top(ctrl_T_top[2]),
    .Tile_X10Y3_A_O_top_0_t(ctrl_O_top_0_t[2]),
    .Tile_X10Y3_A_O_top_0_f(ctrl_O_top_0_f[2]),
    .Tile_X10Y4_A_I_top_0_t(ctrl_I_top_0_t[3]),
    .Tile_X10Y4_A_I_top_0_f(ctrl_I_top_0_f[3]),
    .Tile_X10Y4_A_T_top(ctrl_T_top[3]),
    .Tile_X10Y4_A_O_top_0_t(ctrl_O_top_0_t[3]),
    .Tile_X10Y4_A_O_top_0_f(ctrl_O_top_0_f[3]),
    .Tile_X10Y5_A_I_top_0_t(ctrl_I_top_0_t[4]),
    .Tile_X10Y5_A_I_top_0_f(ctrl_I_top_0_f[4]),
    .Tile_X10Y5_A_T_top(ctrl_T_top[4]),
    .Tile_X10Y5_A_O_top_0_t(ctrl_O_top_0_t[4]),
    .Tile_X10Y5_A_O_top_0_f(ctrl_O_top_0_f[4]),
    .Tile_X10Y6_A_I_top_0_t(ctrl_I_top_0_t[5]),
    .Tile_X10Y6_A_I_top_0_f(ctrl_I_top_0_f[5]),
    .Tile_X10Y6_A_T_top(ctrl_T_top[5]),
    .Tile_X10Y6_A_O_top_0_t(ctrl_O_top_0_t[5]),
    .Tile_X10Y6_A_O_top_0_f(ctrl_O_top_0_f[5]),
    .Tile_X10Y7_A_I_top_0_t(ctrl_I_top_0_t[6]),
    .Tile_X10Y7_A_I_top_0_f(ctrl_I_top_0_f[6]),
    .Tile_X10Y7_A_T_top(ctrl_T_top[6]),
    .Tile_X10Y7_A_O_top_0_t(ctrl_O_top_0_t[6]),
    .Tile_X10Y7_A_O_top_0_f(ctrl_O_top_0_f[6]),
    .Tile_X10Y8_A_I_top_0_t(ctrl_I_top_0_t[7]),
    .Tile_X10Y8_A_I_top_0_f(ctrl_I_top_0_f[7]),
    .Tile_X10Y8_A_T_top(ctrl_T_top[7]),
    .Tile_X10Y8_A_O_top_0_t(ctrl_O_top_0_t[7]),
    .Tile_X10Y8_A_O_top_0_f(ctrl_O_top_0_f[7]),
    .Tile_X10Y9_A_I_top_0_t(ctrl_I_top_0_t[8]),
    .Tile_X10Y9_A_I_top_0_f(ctrl_I_top_0_f[8]),
    .Tile_X10Y9_A_T_top(ctrl_T_top[8]),
    .Tile_X10Y9_A_O_top_0_t(ctrl_O_top_0_t[8]),
    .Tile_X10Y9_A_O_top_0_f(ctrl_O_top_0_f[8]),
    .Tile_X10Y10_A_I_top_0_t(ctrl_I_top_0_t[9]),
    .Tile_X10Y10_A_I_top_0_f(ctrl_I_top_0_f[9]),
    .Tile_X10Y10_A_T_top(ctrl_T_top[9]),
    .Tile_X10Y10_A_O_top_0_t(ctrl_O_top_0_t[9]),
    .Tile_X10Y10_A_O_top_0_f(ctrl_O_top_0_f[9]),
    .Tile_X10Y11_A_I_top_0_t(ctrl_I_top_0_t[10]),
    .Tile_X10Y11_A_I_top_0_f(ctrl_I_top_0_f[10]),
    .Tile_X10Y11_A_T_top(ctrl_T_top[10]),
    .Tile_X10Y11_A_O_top_0_t(ctrl_O_top_0_t[10]),
    .Tile_X10Y11_A_O_top_0_f(ctrl_O_top_0_f[10]),
    .Tile_X10Y12_A_I_top_0_t(ctrl_I_top_0_t[11]),
    .Tile_X10Y12_A_I_top_0_f(ctrl_I_top_0_f[11]),
    .Tile_X10Y12_A_T_top(ctrl_T_top[11]),
    .Tile_X10Y12_A_O_top_0_t(ctrl_O_top_0_t[11]),
    .Tile_X10Y12_A_O_top_0_f(ctrl_O_top_0_f[11]),
    .Tile_X10Y13_A_I_top_0_t(ctrl_I_top_0_t[12]),
    .Tile_X10Y13_A_I_top_0_f(ctrl_I_top_0_f[12]),
    .Tile_X10Y13_A_T_top(ctrl_T_top[12]),
    .Tile_X10Y13_A_O_top_0_t(ctrl_O_top_0_t[12]),
    .Tile_X10Y13_A_O_top_0_f(ctrl_O_top_0_f[12]),
    .Tile_X10Y14_A_I_top_0_t(ctrl_I_top_0_t[13]),
    .Tile_X10Y14_A_I_top_0_f(ctrl_I_top_0_f[13]),
    .Tile_X10Y14_A_T_top(ctrl_T_top[13]),
    .Tile_X10Y14_A_O_top_0_t(ctrl_O_top_0_t[13]),
    .Tile_X10Y14_A_O_top_0_f(ctrl_O_top_0_f[13]),
    .Tile_X10Y15_A_I_top_0_t(ctrl_I_top_0_t[14]),
    .Tile_X10Y15_A_I_top_0_f(ctrl_I_top_0_f[14]),
    .Tile_X10Y15_A_T_top(ctrl_T_top[14]),
    .Tile_X10Y15_A_O_top_0_t(ctrl_O_top_0_t[14]),
    .Tile_X10Y15_A_O_top_0_f(ctrl_O_top_0_f[14]),
    .Tile_X10Y16_A_I_top_0_t(ctrl_I_top_0_t[15]),
    .Tile_X10Y16_A_I_top_0_f(ctrl_I_top_0_f[15]),
    .Tile_X10Y16_A_T_top(ctrl_T_top[15]),
    .Tile_X10Y16_A_O_top_0_t(ctrl_O_top_0_t[15]),
    .Tile_X10Y16_A_O_top_0_f(ctrl_O_top_0_f[15]),
    .Tile_X10Y17_A_I_top_0_t(ctrl_I_top_0_t[16]),
    .Tile_X10Y17_A_I_top_0_f(ctrl_I_top_0_f[16]),
    .Tile_X10Y17_A_T_top(ctrl_T_top[16]),
    .Tile_X10Y17_A_O_top_0_t(ctrl_O_top_0_t[16]),
    .Tile_X10Y17_A_O_top_0_f(ctrl_O_top_0_f[16]),
    .Tile_X10Y18_A_I_top_0_t(ctrl_I_top_0_t[17]),
    .Tile_X10Y18_A_I_top_0_f(ctrl_I_top_0_f[17]),
    .Tile_X10Y18_A_T_top(ctrl_T_top[17]),
    .Tile_X10Y18_A_O_top_0_t(ctrl_O_top_0_t[17]),
    .Tile_X10Y18_A_O_top_0_f(ctrl_O_top_0_f[17]),
    .Tile_X10Y19_A_I_top_0_t(ctrl_I_top_0_t[18]),
    .Tile_X10Y19_A_I_top_0_f(ctrl_I_top_0_f[18]),
    .Tile_X10Y19_A_T_top(ctrl_T_top[18]),
    .Tile_X10Y19_A_O_top_0_t(ctrl_O_top_0_t[18]),
    .Tile_X10Y19_A_O_top_0_f(ctrl_O_top_0_f[18]),
    .Tile_X10Y20_A_I_top_0_t(ctrl_I_top_0_t[19]),
    .Tile_X10Y20_A_I_top_0_f(ctrl_I_top_0_f[19]),
    .Tile_X10Y20_A_T_top(ctrl_T_top[19]),
    .Tile_X10Y20_A_O_top_0_t(ctrl_O_top_0_t[19]),
    .Tile_X10Y20_A_O_top_0_f(ctrl_O_top_0_f[19]),
    .Tile_X10Y21_A_I_top_0_t(ctrl_I_top_0_t[20]),
    .Tile_X10Y21_A_I_top_0_f(ctrl_I_top_0_f[20]),
    .Tile_X10Y21_A_T_top(ctrl_T_top[20]),
    .Tile_X10Y21_A_O_top_0_t(ctrl_O_top_0_t[20]),
    .Tile_X10Y21_A_O_top_0_f(ctrl_O_top_0_f[20]),
    .Tile_X10Y22_A_I_top_0_t(ctrl_I_top_0_t[21]),
    .Tile_X10Y22_A_I_top_0_f(ctrl_I_top_0_f[21]),
    .Tile_X10Y22_A_T_top(ctrl_T_top[21]),
    .Tile_X10Y22_A_O_top_0_t(ctrl_O_top_0_t[21]),
    .Tile_X10Y22_A_O_top_0_f(ctrl_O_top_0_f[21]),
    .Tile_X10Y23_A_I_top_0_t(ctrl_I_top_0_t[22]),
    .Tile_X10Y23_A_I_top_0_f(ctrl_I_top_0_f[22]),
    .Tile_X10Y23_A_T_top(ctrl_T_top[22]),
    .Tile_X10Y23_A_O_top_0_t(ctrl_O_top_0_t[22]),
    .Tile_X10Y23_A_O_top_0_f(ctrl_O_top_0_f[22]),
    .rst(rst),
    .Tile_X0Y1_A_config_C_bit0(A_config_C[91]),
    .Tile_X0Y1_A_config_C_bit1(A_config_C[90]),
    .Tile_X0Y1_A_config_C_bit2(A_config_C[89]),
    .Tile_X0Y1_A_config_C_bit3(A_config_C[88]),
    .Tile_X0Y2_A_config_C_bit0(A_config_C[87]),
    .Tile_X0Y2_A_config_C_bit1(A_config_C[86]),
    .Tile_X0Y2_A_config_C_bit2(A_config_C[85]),
    .Tile_X0Y2_A_config_C_bit3(A_config_C[84]),
    .Tile_X0Y3_A_config_C_bit0(A_config_C[83]),
    .Tile_X0Y3_A_config_C_bit1(A_config_C[82]),
    .Tile_X0Y3_A_config_C_bit2(A_config_C[81]),
    .Tile_X0Y3_A_config_C_bit3(A_config_C[80]),
    .Tile_X0Y4_A_config_C_bit0(A_config_C[79]),
    .Tile_X0Y4_A_config_C_bit1(A_config_C[78]),
    .Tile_X0Y4_A_config_C_bit2(A_config_C[77]),
    .Tile_X0Y4_A_config_C_bit3(A_config_C[76]),
    .Tile_X0Y5_A_config_C_bit0(A_config_C[75]),
    .Tile_X0Y5_A_config_C_bit1(A_config_C[74]),
    .Tile_X0Y5_A_config_C_bit2(A_config_C[73]),
    .Tile_X0Y5_A_config_C_bit3(A_config_C[72]),
    .Tile_X0Y6_A_config_C_bit0(A_config_C[71]),
    .Tile_X0Y6_A_config_C_bit1(A_config_C[70]),
    .Tile_X0Y6_A_config_C_bit2(A_config_C[69]),
    .Tile_X0Y6_A_config_C_bit3(A_config_C[68]),
    .Tile_X0Y7_A_config_C_bit0(A_config_C[67]),
    .Tile_X0Y7_A_config_C_bit1(A_config_C[66]),
    .Tile_X0Y7_A_config_C_bit2(A_config_C[65]),
    .Tile_X0Y7_A_config_C_bit3(A_config_C[64]),
    .Tile_X0Y8_A_config_C_bit0(A_config_C[63]),
    .Tile_X0Y8_A_config_C_bit1(A_config_C[62]),
    .Tile_X0Y8_A_config_C_bit2(A_config_C[61]),
    .Tile_X0Y8_A_config_C_bit3(A_config_C[60]),
    .Tile_X0Y9_A_config_C_bit0(A_config_C[59]),
    .Tile_X0Y9_A_config_C_bit1(A_config_C[58]),
    .Tile_X0Y9_A_config_C_bit2(A_config_C[57]),
    .Tile_X0Y9_A_config_C_bit3(A_config_C[56]),
    .Tile_X0Y10_A_config_C_bit0(A_config_C[55]),
    .Tile_X0Y10_A_config_C_bit1(A_config_C[54]),
    .Tile_X0Y10_A_config_C_bit2(A_config_C[53]),
    .Tile_X0Y10_A_config_C_bit3(A_config_C[52]),
    .Tile_X0Y11_A_config_C_bit0(A_config_C[51]),
    .Tile_X0Y11_A_config_C_bit1(A_config_C[50]),
    .Tile_X0Y11_A_config_C_bit2(A_config_C[49]),
    .Tile_X0Y11_A_config_C_bit3(A_config_C[48]),
    .Tile_X0Y12_A_config_C_bit0(A_config_C[47]),
    .Tile_X0Y12_A_config_C_bit1(A_config_C[46]),
    .Tile_X0Y12_A_config_C_bit2(A_config_C[45]),
    .Tile_X0Y12_A_config_C_bit3(A_config_C[44]),
    .Tile_X0Y13_A_config_C_bit0(A_config_C[43]),
    .Tile_X0Y13_A_config_C_bit1(A_config_C[42]),
    .Tile_X0Y13_A_config_C_bit2(A_config_C[41]),
    .Tile_X0Y13_A_config_C_bit3(A_config_C[40]),
    .Tile_X0Y14_A_config_C_bit0(A_config_C[39]),
    .Tile_X0Y14_A_config_C_bit1(A_config_C[38]),
    .Tile_X0Y14_A_config_C_bit2(A_config_C[37]),
    .Tile_X0Y14_A_config_C_bit3(A_config_C[36]),
    .Tile_X0Y15_A_config_C_bit0(A_config_C[35]),
    .Tile_X0Y15_A_config_C_bit1(A_config_C[34]),
    .Tile_X0Y15_A_config_C_bit2(A_config_C[33]),
    .Tile_X0Y15_A_config_C_bit3(A_config_C[32]),
    .Tile_X0Y16_A_config_C_bit0(A_config_C[31]),
    .Tile_X0Y16_A_config_C_bit1(A_config_C[30]),
    .Tile_X0Y16_A_config_C_bit2(A_config_C[29]),
    .Tile_X0Y16_A_config_C_bit3(A_config_C[28]),
    .Tile_X0Y17_A_config_C_bit0(A_config_C[27]),
    .Tile_X0Y17_A_config_C_bit1(A_config_C[26]),
    .Tile_X0Y17_A_config_C_bit2(A_config_C[25]),
    .Tile_X0Y17_A_config_C_bit3(A_config_C[24]),
    .Tile_X0Y18_A_config_C_bit0(A_config_C[23]),
    .Tile_X0Y18_A_config_C_bit1(A_config_C[22]),
    .Tile_X0Y18_A_config_C_bit2(A_config_C[21]),
    .Tile_X0Y18_A_config_C_bit3(A_config_C[20]),
    .Tile_X0Y19_A_config_C_bit0(A_config_C[19]),
    .Tile_X0Y19_A_config_C_bit1(A_config_C[18]),
    .Tile_X0Y19_A_config_C_bit2(A_config_C[17]),
    .Tile_X0Y19_A_config_C_bit3(A_config_C[16]),
    .Tile_X0Y20_A_config_C_bit0(A_config_C[15]),
    .Tile_X0Y20_A_config_C_bit1(A_config_C[14]),
    .Tile_X0Y20_A_config_C_bit2(A_config_C[13]),
    .Tile_X0Y20_A_config_C_bit3(A_config_C[12]),
    .Tile_X0Y21_A_config_C_bit0(A_config_C[11]),
    .Tile_X0Y21_A_config_C_bit1(A_config_C[10]),
    .Tile_X0Y21_A_config_C_bit2(A_config_C[9]),
    .Tile_X0Y21_A_config_C_bit3(A_config_C[8]),
    .Tile_X0Y22_A_config_C_bit0(A_config_C[7]),
    .Tile_X0Y22_A_config_C_bit1(A_config_C[6]),
    .Tile_X0Y22_A_config_C_bit2(A_config_C[5]),
    .Tile_X0Y22_A_config_C_bit3(A_config_C[4]),
    .Tile_X0Y23_A_config_C_bit0(A_config_C[3]),
    .Tile_X0Y23_A_config_C_bit1(A_config_C[2]),
    .Tile_X0Y23_A_config_C_bit2(A_config_C[1]),
    .Tile_X0Y23_A_config_C_bit3(A_config_C[0]),
    .Tile_X0Y1_B_config_C_bit0(B_config_C[91]),
    .Tile_X0Y1_B_config_C_bit1(B_config_C[90]),
    .Tile_X0Y1_B_config_C_bit2(B_config_C[89]),
    .Tile_X0Y1_B_config_C_bit3(B_config_C[88]),
    .Tile_X0Y2_B_config_C_bit0(B_config_C[87]),
    .Tile_X0Y2_B_config_C_bit1(B_config_C[86]),
    .Tile_X0Y2_B_config_C_bit2(B_config_C[85]),
    .Tile_X0Y2_B_config_C_bit3(B_config_C[84]),
    .Tile_X0Y3_B_config_C_bit0(B_config_C[83]),
    .Tile_X0Y3_B_config_C_bit1(B_config_C[82]),
    .Tile_X0Y3_B_config_C_bit2(B_config_C[81]),
    .Tile_X0Y3_B_config_C_bit3(B_config_C[80]),
    .Tile_X0Y4_B_config_C_bit0(B_config_C[79]),
    .Tile_X0Y4_B_config_C_bit1(B_config_C[78]),
    .Tile_X0Y4_B_config_C_bit2(B_config_C[77]),
    .Tile_X0Y4_B_config_C_bit3(B_config_C[76]),
    .Tile_X0Y5_B_config_C_bit0(B_config_C[75]),
    .Tile_X0Y5_B_config_C_bit1(B_config_C[74]),
    .Tile_X0Y5_B_config_C_bit2(B_config_C[73]),
    .Tile_X0Y5_B_config_C_bit3(B_config_C[72]),
    .Tile_X0Y6_B_config_C_bit0(B_config_C[71]),
    .Tile_X0Y6_B_config_C_bit1(B_config_C[70]),
    .Tile_X0Y6_B_config_C_bit2(B_config_C[69]),
    .Tile_X0Y6_B_config_C_bit3(B_config_C[68]),
    .Tile_X0Y7_B_config_C_bit0(B_config_C[67]),
    .Tile_X0Y7_B_config_C_bit1(B_config_C[66]),
    .Tile_X0Y7_B_config_C_bit2(B_config_C[65]),
    .Tile_X0Y7_B_config_C_bit3(B_config_C[64]),
    .Tile_X0Y8_B_config_C_bit0(B_config_C[63]),
    .Tile_X0Y8_B_config_C_bit1(B_config_C[62]),
    .Tile_X0Y8_B_config_C_bit2(B_config_C[61]),
    .Tile_X0Y8_B_config_C_bit3(B_config_C[60]),
    .Tile_X0Y9_B_config_C_bit0(B_config_C[59]),
    .Tile_X0Y9_B_config_C_bit1(B_config_C[58]),
    .Tile_X0Y9_B_config_C_bit2(B_config_C[57]),
    .Tile_X0Y9_B_config_C_bit3(B_config_C[56]),
    .Tile_X0Y10_B_config_C_bit0(B_config_C[55]),
    .Tile_X0Y10_B_config_C_bit1(B_config_C[54]),
    .Tile_X0Y10_B_config_C_bit2(B_config_C[53]),
    .Tile_X0Y10_B_config_C_bit3(B_config_C[52]),
    .Tile_X0Y11_B_config_C_bit0(B_config_C[51]),
    .Tile_X0Y11_B_config_C_bit1(B_config_C[50]),
    .Tile_X0Y11_B_config_C_bit2(B_config_C[49]),
    .Tile_X0Y11_B_config_C_bit3(B_config_C[48]),
    .Tile_X0Y12_B_config_C_bit0(B_config_C[47]),
    .Tile_X0Y12_B_config_C_bit1(B_config_C[46]),
    .Tile_X0Y12_B_config_C_bit2(B_config_C[45]),
    .Tile_X0Y12_B_config_C_bit3(B_config_C[44]),
    .Tile_X0Y13_B_config_C_bit0(B_config_C[43]),
    .Tile_X0Y13_B_config_C_bit1(B_config_C[42]),
    .Tile_X0Y13_B_config_C_bit2(B_config_C[41]),
    .Tile_X0Y13_B_config_C_bit3(B_config_C[40]),
    .Tile_X0Y14_B_config_C_bit0(B_config_C[39]),
    .Tile_X0Y14_B_config_C_bit1(B_config_C[38]),
    .Tile_X0Y14_B_config_C_bit2(B_config_C[37]),
    .Tile_X0Y14_B_config_C_bit3(B_config_C[36]),
    .Tile_X0Y15_B_config_C_bit0(B_config_C[35]),
    .Tile_X0Y15_B_config_C_bit1(B_config_C[34]),
    .Tile_X0Y15_B_config_C_bit2(B_config_C[33]),
    .Tile_X0Y15_B_config_C_bit3(B_config_C[32]),
    .Tile_X0Y16_B_config_C_bit0(B_config_C[31]),
    .Tile_X0Y16_B_config_C_bit1(B_config_C[30]),
    .Tile_X0Y16_B_config_C_bit2(B_config_C[29]),
    .Tile_X0Y16_B_config_C_bit3(B_config_C[28]),
    .Tile_X0Y17_B_config_C_bit0(B_config_C[27]),
    .Tile_X0Y17_B_config_C_bit1(B_config_C[26]),
    .Tile_X0Y17_B_config_C_bit2(B_config_C[25]),
    .Tile_X0Y17_B_config_C_bit3(B_config_C[24]),
    .Tile_X0Y18_B_config_C_bit0(B_config_C[23]),
    .Tile_X0Y18_B_config_C_bit1(B_config_C[22]),
    .Tile_X0Y18_B_config_C_bit2(B_config_C[21]),
    .Tile_X0Y18_B_config_C_bit3(B_config_C[20]),
    .Tile_X0Y19_B_config_C_bit0(B_config_C[19]),
    .Tile_X0Y19_B_config_C_bit1(B_config_C[18]),
    .Tile_X0Y19_B_config_C_bit2(B_config_C[17]),
    .Tile_X0Y19_B_config_C_bit3(B_config_C[16]),
    .Tile_X0Y20_B_config_C_bit0(B_config_C[15]),
    .Tile_X0Y20_B_config_C_bit1(B_config_C[14]),
    .Tile_X0Y20_B_config_C_bit2(B_config_C[13]),
    .Tile_X0Y20_B_config_C_bit3(B_config_C[12]),
    .Tile_X0Y21_B_config_C_bit0(B_config_C[11]),
    .Tile_X0Y21_B_config_C_bit1(B_config_C[10]),
    .Tile_X0Y21_B_config_C_bit2(B_config_C[9]),
    .Tile_X0Y21_B_config_C_bit3(B_config_C[8]),
    .Tile_X0Y22_B_config_C_bit0(B_config_C[7]),
    .Tile_X0Y22_B_config_C_bit1(B_config_C[6]),
    .Tile_X0Y22_B_config_C_bit2(B_config_C[5]),
    .Tile_X0Y22_B_config_C_bit3(B_config_C[4]),
    .Tile_X0Y23_B_config_C_bit0(B_config_C[3]),
    .Tile_X0Y23_B_config_C_bit1(B_config_C[2]),
    .Tile_X0Y23_B_config_C_bit2(B_config_C[1]),
    .Tile_X0Y23_B_config_C_bit3(B_config_C[0]),
    .UserCLK(CLK),
    .FrameData(FrameData),
    .FrameStrobe(FrameSelect)
);


fault_detector  #(.Nm1(22), .Nm2(22), .Nctrl(22)) DR_check (
    .CLK(CLK),
    .rst(rst),
    .prech1(prech1),
    .prech2(prech2),
    .f_m1(F_masked1_top),
    .f_m2(F_masked2_top),
    .f_ctrl(F_ctrl_top),
    .f_detected(f_detected)
);

prech_signal_module prech_signal_module_i (
    .rst(rst),
    .CLK(CLK),
    .prech1(prech1),
    .prech2(prech2)
);

Trivium_DRP  #(.output_bits(575)) Trivium_DRP_i (
    .clk(CLK),
    .rst(prng_rst),
    .prech1(prech1),
    .key_t(key_t),
    .key_f(key_f),
    .iv_t(iv_t),
    .iv_f(iv_f),
    .stream_out_t(R_t_top),
    .stream_out_f(R_f_top)
);

assign FrameData = {32'h12345678,FrameRegister,32'h12345678};
endmodule