/* modified netlist. Source: module Cipher in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/10_CRAFT_round_based_encryption_PortParallel/4-AGEMA/Cipher.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module Cipher_SAUBER_Pipeline_d1 (Input, Key, rst, Output, done);
    input [63:0] Input ;
    input [127:0] Key ;
    input rst ;
    output [63:0] Output ;
    output done ;
    wire RoundConstant_4_ ;
    wire RoundConstant_0 ;
    wire InputMUX_MUXInst_0_U1_Y ;
    wire InputMUX_MUXInst_0_U1_X ;
    wire InputMUX_MUXInst_1_U1_Y ;
    wire InputMUX_MUXInst_1_U1_X ;
    wire InputMUX_MUXInst_2_U1_Y ;
    wire InputMUX_MUXInst_2_U1_X ;
    wire InputMUX_MUXInst_3_U1_Y ;
    wire InputMUX_MUXInst_3_U1_X ;
    wire InputMUX_MUXInst_4_U1_Y ;
    wire InputMUX_MUXInst_4_U1_X ;
    wire InputMUX_MUXInst_5_U1_Y ;
    wire InputMUX_MUXInst_5_U1_X ;
    wire InputMUX_MUXInst_6_U1_Y ;
    wire InputMUX_MUXInst_6_U1_X ;
    wire InputMUX_MUXInst_7_U1_Y ;
    wire InputMUX_MUXInst_7_U1_X ;
    wire InputMUX_MUXInst_8_U1_Y ;
    wire InputMUX_MUXInst_8_U1_X ;
    wire InputMUX_MUXInst_9_U1_Y ;
    wire InputMUX_MUXInst_9_U1_X ;
    wire InputMUX_MUXInst_10_U1_Y ;
    wire InputMUX_MUXInst_10_U1_X ;
    wire InputMUX_MUXInst_11_U1_Y ;
    wire InputMUX_MUXInst_11_U1_X ;
    wire InputMUX_MUXInst_12_U1_Y ;
    wire InputMUX_MUXInst_12_U1_X ;
    wire InputMUX_MUXInst_13_U1_Y ;
    wire InputMUX_MUXInst_13_U1_X ;
    wire InputMUX_MUXInst_14_U1_Y ;
    wire InputMUX_MUXInst_14_U1_X ;
    wire InputMUX_MUXInst_15_U1_Y ;
    wire InputMUX_MUXInst_15_U1_X ;
    wire InputMUX_MUXInst_16_U1_Y ;
    wire InputMUX_MUXInst_16_U1_X ;
    wire InputMUX_MUXInst_17_U1_Y ;
    wire InputMUX_MUXInst_17_U1_X ;
    wire InputMUX_MUXInst_18_U1_Y ;
    wire InputMUX_MUXInst_18_U1_X ;
    wire InputMUX_MUXInst_19_U1_Y ;
    wire InputMUX_MUXInst_19_U1_X ;
    wire InputMUX_MUXInst_20_U1_Y ;
    wire InputMUX_MUXInst_20_U1_X ;
    wire InputMUX_MUXInst_21_U1_Y ;
    wire InputMUX_MUXInst_21_U1_X ;
    wire InputMUX_MUXInst_22_U1_Y ;
    wire InputMUX_MUXInst_22_U1_X ;
    wire InputMUX_MUXInst_23_U1_Y ;
    wire InputMUX_MUXInst_23_U1_X ;
    wire InputMUX_MUXInst_24_U1_Y ;
    wire InputMUX_MUXInst_24_U1_X ;
    wire InputMUX_MUXInst_25_U1_Y ;
    wire InputMUX_MUXInst_25_U1_X ;
    wire InputMUX_MUXInst_26_U1_Y ;
    wire InputMUX_MUXInst_26_U1_X ;
    wire InputMUX_MUXInst_27_U1_Y ;
    wire InputMUX_MUXInst_27_U1_X ;
    wire InputMUX_MUXInst_28_U1_Y ;
    wire InputMUX_MUXInst_28_U1_X ;
    wire InputMUX_MUXInst_29_U1_Y ;
    wire InputMUX_MUXInst_29_U1_X ;
    wire InputMUX_MUXInst_30_U1_Y ;
    wire InputMUX_MUXInst_30_U1_X ;
    wire InputMUX_MUXInst_31_U1_Y ;
    wire InputMUX_MUXInst_31_U1_X ;
    wire InputMUX_MUXInst_32_U1_Y ;
    wire InputMUX_MUXInst_32_U1_X ;
    wire InputMUX_MUXInst_33_U1_Y ;
    wire InputMUX_MUXInst_33_U1_X ;
    wire InputMUX_MUXInst_34_U1_Y ;
    wire InputMUX_MUXInst_34_U1_X ;
    wire InputMUX_MUXInst_35_U1_Y ;
    wire InputMUX_MUXInst_35_U1_X ;
    wire InputMUX_MUXInst_36_U1_Y ;
    wire InputMUX_MUXInst_36_U1_X ;
    wire InputMUX_MUXInst_37_U1_Y ;
    wire InputMUX_MUXInst_37_U1_X ;
    wire InputMUX_MUXInst_38_U1_Y ;
    wire InputMUX_MUXInst_38_U1_X ;
    wire InputMUX_MUXInst_39_U1_Y ;
    wire InputMUX_MUXInst_39_U1_X ;
    wire InputMUX_MUXInst_40_U1_Y ;
    wire InputMUX_MUXInst_40_U1_X ;
    wire InputMUX_MUXInst_41_U1_Y ;
    wire InputMUX_MUXInst_41_U1_X ;
    wire InputMUX_MUXInst_42_U1_Y ;
    wire InputMUX_MUXInst_42_U1_X ;
    wire InputMUX_MUXInst_43_U1_Y ;
    wire InputMUX_MUXInst_43_U1_X ;
    wire InputMUX_MUXInst_44_U1_Y ;
    wire InputMUX_MUXInst_44_U1_X ;
    wire InputMUX_MUXInst_45_U1_Y ;
    wire InputMUX_MUXInst_45_U1_X ;
    wire InputMUX_MUXInst_46_U1_Y ;
    wire InputMUX_MUXInst_46_U1_X ;
    wire InputMUX_MUXInst_47_U1_Y ;
    wire InputMUX_MUXInst_47_U1_X ;
    wire InputMUX_MUXInst_48_U1_Y ;
    wire InputMUX_MUXInst_48_U1_X ;
    wire InputMUX_MUXInst_49_U1_Y ;
    wire InputMUX_MUXInst_49_U1_X ;
    wire InputMUX_MUXInst_50_U1_Y ;
    wire InputMUX_MUXInst_50_U1_X ;
    wire InputMUX_MUXInst_51_U1_Y ;
    wire InputMUX_MUXInst_51_U1_X ;
    wire InputMUX_MUXInst_52_U1_Y ;
    wire InputMUX_MUXInst_52_U1_X ;
    wire InputMUX_MUXInst_53_U1_Y ;
    wire InputMUX_MUXInst_53_U1_X ;
    wire InputMUX_MUXInst_54_U1_Y ;
    wire InputMUX_MUXInst_54_U1_X ;
    wire InputMUX_MUXInst_55_U1_Y ;
    wire InputMUX_MUXInst_55_U1_X ;
    wire InputMUX_MUXInst_56_U1_Y ;
    wire InputMUX_MUXInst_56_U1_X ;
    wire InputMUX_MUXInst_57_U1_Y ;
    wire InputMUX_MUXInst_57_U1_X ;
    wire InputMUX_MUXInst_58_U1_Y ;
    wire InputMUX_MUXInst_58_U1_X ;
    wire InputMUX_MUXInst_59_U1_Y ;
    wire InputMUX_MUXInst_59_U1_X ;
    wire InputMUX_MUXInst_60_U1_Y ;
    wire InputMUX_MUXInst_60_U1_X ;
    wire InputMUX_MUXInst_61_U1_Y ;
    wire InputMUX_MUXInst_61_U1_X ;
    wire InputMUX_MUXInst_62_U1_Y ;
    wire InputMUX_MUXInst_62_U1_X ;
    wire InputMUX_MUXInst_63_U1_Y ;
    wire InputMUX_MUXInst_63_U1_X ;
    wire MCInst_XOR_r0_Inst_0_n1 ;
    wire MCInst_XOR_r0_Inst_1_n1 ;
    wire MCInst_XOR_r0_Inst_2_n1 ;
    wire MCInst_XOR_r0_Inst_3_n1 ;
    wire MCInst_XOR_r0_Inst_4_n1 ;
    wire MCInst_XOR_r0_Inst_5_n1 ;
    wire MCInst_XOR_r0_Inst_6_n1 ;
    wire MCInst_XOR_r0_Inst_7_n1 ;
    wire MCInst_XOR_r0_Inst_8_n1 ;
    wire MCInst_XOR_r0_Inst_9_n1 ;
    wire MCInst_XOR_r0_Inst_10_n1 ;
    wire MCInst_XOR_r0_Inst_11_n1 ;
    wire MCInst_XOR_r0_Inst_12_n1 ;
    wire MCInst_XOR_r0_Inst_13_n1 ;
    wire MCInst_XOR_r0_Inst_14_n1 ;
    wire MCInst_XOR_r0_Inst_15_n1 ;
    wire AddKeyConstXOR_XORInst_0_0_n1 ;
    wire AddKeyConstXOR_XORInst_0_1_n1 ;
    wire AddKeyConstXOR_XORInst_0_2_n1 ;
    wire AddKeyConstXOR_XORInst_1_0_n1 ;
    wire AddKeyConstXOR_XORInst_1_1_n1 ;
    wire AddKeyConstXOR_XORInst_1_2_n1 ;
    wire AddKeyConstXOR_XORInst_1_3_n1 ;
    wire SubCellInst_SboxInst_0_n15 ;
    wire SubCellInst_SboxInst_0_n14 ;
    wire SubCellInst_SboxInst_0_n13 ;
    wire SubCellInst_SboxInst_0_n11 ;
    wire SubCellInst_SboxInst_0_n10 ;
    wire SubCellInst_SboxInst_0_n9 ;
    wire SubCellInst_SboxInst_0_n7 ;
    wire SubCellInst_SboxInst_0_n6 ;
    wire SubCellInst_SboxInst_0_n5 ;
    wire SubCellInst_SboxInst_0_n4 ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_n1 ;
    wire SubCellInst_SboxInst_1_n15 ;
    wire SubCellInst_SboxInst_1_n14 ;
    wire SubCellInst_SboxInst_1_n13 ;
    wire SubCellInst_SboxInst_1_n11 ;
    wire SubCellInst_SboxInst_1_n10 ;
    wire SubCellInst_SboxInst_1_n9 ;
    wire SubCellInst_SboxInst_1_n7 ;
    wire SubCellInst_SboxInst_1_n6 ;
    wire SubCellInst_SboxInst_1_n5 ;
    wire SubCellInst_SboxInst_1_n4 ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_n1 ;
    wire SubCellInst_SboxInst_2_n15 ;
    wire SubCellInst_SboxInst_2_n14 ;
    wire SubCellInst_SboxInst_2_n13 ;
    wire SubCellInst_SboxInst_2_n11 ;
    wire SubCellInst_SboxInst_2_n10 ;
    wire SubCellInst_SboxInst_2_n9 ;
    wire SubCellInst_SboxInst_2_n7 ;
    wire SubCellInst_SboxInst_2_n6 ;
    wire SubCellInst_SboxInst_2_n5 ;
    wire SubCellInst_SboxInst_2_n4 ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_n1 ;
    wire SubCellInst_SboxInst_3_n15 ;
    wire SubCellInst_SboxInst_3_n14 ;
    wire SubCellInst_SboxInst_3_n13 ;
    wire SubCellInst_SboxInst_3_n11 ;
    wire SubCellInst_SboxInst_3_n10 ;
    wire SubCellInst_SboxInst_3_n9 ;
    wire SubCellInst_SboxInst_3_n7 ;
    wire SubCellInst_SboxInst_3_n6 ;
    wire SubCellInst_SboxInst_3_n5 ;
    wire SubCellInst_SboxInst_3_n4 ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_n1 ;
    wire SubCellInst_SboxInst_4_n15 ;
    wire SubCellInst_SboxInst_4_n14 ;
    wire SubCellInst_SboxInst_4_n13 ;
    wire SubCellInst_SboxInst_4_n10 ;
    wire SubCellInst_SboxInst_4_n9 ;
    wire SubCellInst_SboxInst_4_n8 ;
    wire SubCellInst_SboxInst_4_n7 ;
    wire SubCellInst_SboxInst_4_n6 ;
    wire SubCellInst_SboxInst_4_n5 ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_n2 ;
    wire SubCellInst_SboxInst_4_n1 ;
    wire SubCellInst_SboxInst_5_n15 ;
    wire SubCellInst_SboxInst_5_n14 ;
    wire SubCellInst_SboxInst_5_n13 ;
    wire SubCellInst_SboxInst_5_n10 ;
    wire SubCellInst_SboxInst_5_n9 ;
    wire SubCellInst_SboxInst_5_n8 ;
    wire SubCellInst_SboxInst_5_n7 ;
    wire SubCellInst_SboxInst_5_n6 ;
    wire SubCellInst_SboxInst_5_n5 ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_n2 ;
    wire SubCellInst_SboxInst_5_n1 ;
    wire SubCellInst_SboxInst_6_n15 ;
    wire SubCellInst_SboxInst_6_n14 ;
    wire SubCellInst_SboxInst_6_n13 ;
    wire SubCellInst_SboxInst_6_n10 ;
    wire SubCellInst_SboxInst_6_n9 ;
    wire SubCellInst_SboxInst_6_n8 ;
    wire SubCellInst_SboxInst_6_n7 ;
    wire SubCellInst_SboxInst_6_n6 ;
    wire SubCellInst_SboxInst_6_n5 ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_n2 ;
    wire SubCellInst_SboxInst_6_n1 ;
    wire SubCellInst_SboxInst_7_n15 ;
    wire SubCellInst_SboxInst_7_n14 ;
    wire SubCellInst_SboxInst_7_n13 ;
    wire SubCellInst_SboxInst_7_n10 ;
    wire SubCellInst_SboxInst_7_n9 ;
    wire SubCellInst_SboxInst_7_n8 ;
    wire SubCellInst_SboxInst_7_n7 ;
    wire SubCellInst_SboxInst_7_n6 ;
    wire SubCellInst_SboxInst_7_n5 ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_n2 ;
    wire SubCellInst_SboxInst_7_n1 ;
    wire SubCellInst_SboxInst_8_n15 ;
    wire SubCellInst_SboxInst_8_n14 ;
    wire SubCellInst_SboxInst_8_n13 ;
    wire SubCellInst_SboxInst_8_n10 ;
    wire SubCellInst_SboxInst_8_n9 ;
    wire SubCellInst_SboxInst_8_n8 ;
    wire SubCellInst_SboxInst_8_n7 ;
    wire SubCellInst_SboxInst_8_n6 ;
    wire SubCellInst_SboxInst_8_n5 ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_n2 ;
    wire SubCellInst_SboxInst_8_n1 ;
    wire SubCellInst_SboxInst_9_n15 ;
    wire SubCellInst_SboxInst_9_n14 ;
    wire SubCellInst_SboxInst_9_n13 ;
    wire SubCellInst_SboxInst_9_n10 ;
    wire SubCellInst_SboxInst_9_n9 ;
    wire SubCellInst_SboxInst_9_n8 ;
    wire SubCellInst_SboxInst_9_n7 ;
    wire SubCellInst_SboxInst_9_n6 ;
    wire SubCellInst_SboxInst_9_n5 ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_n2 ;
    wire SubCellInst_SboxInst_9_n1 ;
    wire SubCellInst_SboxInst_10_n15 ;
    wire SubCellInst_SboxInst_10_n14 ;
    wire SubCellInst_SboxInst_10_n13 ;
    wire SubCellInst_SboxInst_10_n10 ;
    wire SubCellInst_SboxInst_10_n9 ;
    wire SubCellInst_SboxInst_10_n8 ;
    wire SubCellInst_SboxInst_10_n7 ;
    wire SubCellInst_SboxInst_10_n6 ;
    wire SubCellInst_SboxInst_10_n5 ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_n2 ;
    wire SubCellInst_SboxInst_10_n1 ;
    wire SubCellInst_SboxInst_11_n15 ;
    wire SubCellInst_SboxInst_11_n14 ;
    wire SubCellInst_SboxInst_11_n13 ;
    wire SubCellInst_SboxInst_11_n10 ;
    wire SubCellInst_SboxInst_11_n9 ;
    wire SubCellInst_SboxInst_11_n8 ;
    wire SubCellInst_SboxInst_11_n7 ;
    wire SubCellInst_SboxInst_11_n6 ;
    wire SubCellInst_SboxInst_11_n5 ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_n2 ;
    wire SubCellInst_SboxInst_11_n1 ;
    wire SubCellInst_SboxInst_12_n15 ;
    wire SubCellInst_SboxInst_12_n14 ;
    wire SubCellInst_SboxInst_12_n13 ;
    wire SubCellInst_SboxInst_12_n10 ;
    wire SubCellInst_SboxInst_12_n9 ;
    wire SubCellInst_SboxInst_12_n8 ;
    wire SubCellInst_SboxInst_12_n7 ;
    wire SubCellInst_SboxInst_12_n6 ;
    wire SubCellInst_SboxInst_12_n5 ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_n2 ;
    wire SubCellInst_SboxInst_12_n1 ;
    wire SubCellInst_SboxInst_13_n15 ;
    wire SubCellInst_SboxInst_13_n14 ;
    wire SubCellInst_SboxInst_13_n13 ;
    wire SubCellInst_SboxInst_13_n10 ;
    wire SubCellInst_SboxInst_13_n9 ;
    wire SubCellInst_SboxInst_13_n8 ;
    wire SubCellInst_SboxInst_13_n7 ;
    wire SubCellInst_SboxInst_13_n6 ;
    wire SubCellInst_SboxInst_13_n5 ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_n2 ;
    wire SubCellInst_SboxInst_13_n1 ;
    wire SubCellInst_SboxInst_14_n15 ;
    wire SubCellInst_SboxInst_14_n14 ;
    wire SubCellInst_SboxInst_14_n13 ;
    wire SubCellInst_SboxInst_14_n10 ;
    wire SubCellInst_SboxInst_14_n9 ;
    wire SubCellInst_SboxInst_14_n8 ;
    wire SubCellInst_SboxInst_14_n7 ;
    wire SubCellInst_SboxInst_14_n6 ;
    wire SubCellInst_SboxInst_14_n5 ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_n2 ;
    wire SubCellInst_SboxInst_14_n1 ;
    wire SubCellInst_SboxInst_15_n15 ;
    wire SubCellInst_SboxInst_15_n14 ;
    wire SubCellInst_SboxInst_15_n13 ;
    wire SubCellInst_SboxInst_15_n10 ;
    wire SubCellInst_SboxInst_15_n9 ;
    wire SubCellInst_SboxInst_15_n8 ;
    wire SubCellInst_SboxInst_15_n7 ;
    wire SubCellInst_SboxInst_15_n6 ;
    wire SubCellInst_SboxInst_15_n5 ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_n2 ;
    wire SubCellInst_SboxInst_15_n1 ;
    wire KeyMUX_MUXInst_0_U1_Y ;
    wire KeyMUX_MUXInst_0_U1_X ;
    wire KeyMUX_MUXInst_1_U1_Y ;
    wire KeyMUX_MUXInst_1_U1_X ;
    wire KeyMUX_MUXInst_2_U1_Y ;
    wire KeyMUX_MUXInst_2_U1_X ;
    wire KeyMUX_MUXInst_3_U1_Y ;
    wire KeyMUX_MUXInst_3_U1_X ;
    wire KeyMUX_MUXInst_4_U1_Y ;
    wire KeyMUX_MUXInst_4_U1_X ;
    wire KeyMUX_MUXInst_5_U1_Y ;
    wire KeyMUX_MUXInst_5_U1_X ;
    wire KeyMUX_MUXInst_6_U1_Y ;
    wire KeyMUX_MUXInst_6_U1_X ;
    wire KeyMUX_MUXInst_7_U1_Y ;
    wire KeyMUX_MUXInst_7_U1_X ;
    wire KeyMUX_MUXInst_8_U1_Y ;
    wire KeyMUX_MUXInst_8_U1_X ;
    wire KeyMUX_MUXInst_9_U1_Y ;
    wire KeyMUX_MUXInst_9_U1_X ;
    wire KeyMUX_MUXInst_10_U1_Y ;
    wire KeyMUX_MUXInst_10_U1_X ;
    wire KeyMUX_MUXInst_11_U1_Y ;
    wire KeyMUX_MUXInst_11_U1_X ;
    wire KeyMUX_MUXInst_12_U1_Y ;
    wire KeyMUX_MUXInst_12_U1_X ;
    wire KeyMUX_MUXInst_13_U1_Y ;
    wire KeyMUX_MUXInst_13_U1_X ;
    wire KeyMUX_MUXInst_14_U1_Y ;
    wire KeyMUX_MUXInst_14_U1_X ;
    wire KeyMUX_MUXInst_15_U1_Y ;
    wire KeyMUX_MUXInst_15_U1_X ;
    wire KeyMUX_MUXInst_16_U1_Y ;
    wire KeyMUX_MUXInst_16_U1_X ;
    wire KeyMUX_MUXInst_17_U1_Y ;
    wire KeyMUX_MUXInst_17_U1_X ;
    wire KeyMUX_MUXInst_18_U1_Y ;
    wire KeyMUX_MUXInst_18_U1_X ;
    wire KeyMUX_MUXInst_19_U1_Y ;
    wire KeyMUX_MUXInst_19_U1_X ;
    wire KeyMUX_MUXInst_20_U1_Y ;
    wire KeyMUX_MUXInst_20_U1_X ;
    wire KeyMUX_MUXInst_21_U1_Y ;
    wire KeyMUX_MUXInst_21_U1_X ;
    wire KeyMUX_MUXInst_22_U1_Y ;
    wire KeyMUX_MUXInst_22_U1_X ;
    wire KeyMUX_MUXInst_23_U1_Y ;
    wire KeyMUX_MUXInst_23_U1_X ;
    wire KeyMUX_MUXInst_24_U1_Y ;
    wire KeyMUX_MUXInst_24_U1_X ;
    wire KeyMUX_MUXInst_25_U1_Y ;
    wire KeyMUX_MUXInst_25_U1_X ;
    wire KeyMUX_MUXInst_26_U1_Y ;
    wire KeyMUX_MUXInst_26_U1_X ;
    wire KeyMUX_MUXInst_27_U1_Y ;
    wire KeyMUX_MUXInst_27_U1_X ;
    wire KeyMUX_MUXInst_28_U1_Y ;
    wire KeyMUX_MUXInst_28_U1_X ;
    wire KeyMUX_MUXInst_29_U1_Y ;
    wire KeyMUX_MUXInst_29_U1_X ;
    wire KeyMUX_MUXInst_30_U1_Y ;
    wire KeyMUX_MUXInst_30_U1_X ;
    wire KeyMUX_MUXInst_31_U1_Y ;
    wire KeyMUX_MUXInst_31_U1_X ;
    wire KeyMUX_MUXInst_32_U1_Y ;
    wire KeyMUX_MUXInst_32_U1_X ;
    wire KeyMUX_MUXInst_33_U1_Y ;
    wire KeyMUX_MUXInst_33_U1_X ;
    wire KeyMUX_MUXInst_34_U1_Y ;
    wire KeyMUX_MUXInst_34_U1_X ;
    wire KeyMUX_MUXInst_35_U1_Y ;
    wire KeyMUX_MUXInst_35_U1_X ;
    wire KeyMUX_MUXInst_36_U1_Y ;
    wire KeyMUX_MUXInst_36_U1_X ;
    wire KeyMUX_MUXInst_37_U1_Y ;
    wire KeyMUX_MUXInst_37_U1_X ;
    wire KeyMUX_MUXInst_38_U1_Y ;
    wire KeyMUX_MUXInst_38_U1_X ;
    wire KeyMUX_MUXInst_39_U1_Y ;
    wire KeyMUX_MUXInst_39_U1_X ;
    wire KeyMUX_MUXInst_40_U1_Y ;
    wire KeyMUX_MUXInst_40_U1_X ;
    wire KeyMUX_MUXInst_41_U1_Y ;
    wire KeyMUX_MUXInst_41_U1_X ;
    wire KeyMUX_MUXInst_42_U1_Y ;
    wire KeyMUX_MUXInst_42_U1_X ;
    wire KeyMUX_MUXInst_43_U1_Y ;
    wire KeyMUX_MUXInst_43_U1_X ;
    wire KeyMUX_MUXInst_44_U1_Y ;
    wire KeyMUX_MUXInst_44_U1_X ;
    wire KeyMUX_MUXInst_45_U1_Y ;
    wire KeyMUX_MUXInst_45_U1_X ;
    wire KeyMUX_MUXInst_46_U1_Y ;
    wire KeyMUX_MUXInst_46_U1_X ;
    wire KeyMUX_MUXInst_47_U1_Y ;
    wire KeyMUX_MUXInst_47_U1_X ;
    wire KeyMUX_MUXInst_48_U1_Y ;
    wire KeyMUX_MUXInst_48_U1_X ;
    wire KeyMUX_MUXInst_49_U1_Y ;
    wire KeyMUX_MUXInst_49_U1_X ;
    wire KeyMUX_MUXInst_50_U1_Y ;
    wire KeyMUX_MUXInst_50_U1_X ;
    wire KeyMUX_MUXInst_51_U1_Y ;
    wire KeyMUX_MUXInst_51_U1_X ;
    wire KeyMUX_MUXInst_52_U1_Y ;
    wire KeyMUX_MUXInst_52_U1_X ;
    wire KeyMUX_MUXInst_53_U1_Y ;
    wire KeyMUX_MUXInst_53_U1_X ;
    wire KeyMUX_MUXInst_54_U1_Y ;
    wire KeyMUX_MUXInst_54_U1_X ;
    wire KeyMUX_MUXInst_55_U1_Y ;
    wire KeyMUX_MUXInst_55_U1_X ;
    wire KeyMUX_MUXInst_56_U1_Y ;
    wire KeyMUX_MUXInst_56_U1_X ;
    wire KeyMUX_MUXInst_57_U1_Y ;
    wire KeyMUX_MUXInst_57_U1_X ;
    wire KeyMUX_MUXInst_58_U1_Y ;
    wire KeyMUX_MUXInst_58_U1_X ;
    wire KeyMUX_MUXInst_59_U1_Y ;
    wire KeyMUX_MUXInst_59_U1_X ;
    wire KeyMUX_MUXInst_60_U1_Y ;
    wire KeyMUX_MUXInst_60_U1_X ;
    wire KeyMUX_MUXInst_61_U1_Y ;
    wire KeyMUX_MUXInst_61_U1_X ;
    wire KeyMUX_MUXInst_62_U1_Y ;
    wire KeyMUX_MUXInst_62_U1_X ;
    wire KeyMUX_MUXInst_63_U1_Y ;
    wire KeyMUX_MUXInst_63_U1_X ;
    wire FSMSignalsInst_n5 ;
    wire FSMSignalsInst_n4 ;
    wire FSMSignalsInst_n3 ;
    wire FSMSignalsInst_n2 ;
    wire FSMSignalsInst_n1 ;
    wire [63:0] Feedback ;
    wire [63:32] MCInput ;
    wire [63:0] MCOutput ;
    wire [63:0] SelectedKey ;
    wire [1:0] selects ;
    wire [6:0] FSMReg ;
    wire [5:0] FSMUpdate ;
    wire [1:0] selectsReg ;

    /* cells in depth 0 */
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_0_U1_XOR1_U1 ( .A0_t (Feedback[0]), .B0_t (Input[0]), .Z0_t (InputMUX_MUXInst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_0_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_0_U1_X), .Z0_t (InputMUX_MUXInst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_0_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_0_U1_Y), .B0_t (Feedback[0]), .Z0_t (MCOutput[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_1_U1_XOR1_U1 ( .A0_t (Feedback[1]), .B0_t (Input[1]), .Z0_t (InputMUX_MUXInst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_1_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_1_U1_X), .Z0_t (InputMUX_MUXInst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_1_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_1_U1_Y), .B0_t (Feedback[1]), .Z0_t (MCOutput[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_2_U1_XOR1_U1 ( .A0_t (Feedback[2]), .B0_t (Input[2]), .Z0_t (InputMUX_MUXInst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_2_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_2_U1_X), .Z0_t (InputMUX_MUXInst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_2_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_2_U1_Y), .B0_t (Feedback[2]), .Z0_t (MCOutput[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_3_U1_XOR1_U1 ( .A0_t (Feedback[3]), .B0_t (Input[3]), .Z0_t (InputMUX_MUXInst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_3_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_3_U1_X), .Z0_t (InputMUX_MUXInst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_3_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_3_U1_Y), .B0_t (Feedback[3]), .Z0_t (MCOutput[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_4_U1_XOR1_U1 ( .A0_t (Feedback[4]), .B0_t (Input[4]), .Z0_t (InputMUX_MUXInst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_4_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_4_U1_X), .Z0_t (InputMUX_MUXInst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_4_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_4_U1_Y), .B0_t (Feedback[4]), .Z0_t (MCOutput[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_5_U1_XOR1_U1 ( .A0_t (Feedback[5]), .B0_t (Input[5]), .Z0_t (InputMUX_MUXInst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_5_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_5_U1_X), .Z0_t (InputMUX_MUXInst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_5_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_5_U1_Y), .B0_t (Feedback[5]), .Z0_t (MCOutput[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_6_U1_XOR1_U1 ( .A0_t (Feedback[6]), .B0_t (Input[6]), .Z0_t (InputMUX_MUXInst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_6_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_6_U1_X), .Z0_t (InputMUX_MUXInst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_6_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_6_U1_Y), .B0_t (Feedback[6]), .Z0_t (MCOutput[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_7_U1_XOR1_U1 ( .A0_t (Feedback[7]), .B0_t (Input[7]), .Z0_t (InputMUX_MUXInst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_7_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_7_U1_X), .Z0_t (InputMUX_MUXInst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_7_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_7_U1_Y), .B0_t (Feedback[7]), .Z0_t (MCOutput[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_8_U1_XOR1_U1 ( .A0_t (Feedback[8]), .B0_t (Input[8]), .Z0_t (InputMUX_MUXInst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_8_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_8_U1_X), .Z0_t (InputMUX_MUXInst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_8_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_8_U1_Y), .B0_t (Feedback[8]), .Z0_t (MCOutput[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_9_U1_XOR1_U1 ( .A0_t (Feedback[9]), .B0_t (Input[9]), .Z0_t (InputMUX_MUXInst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_9_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_9_U1_X), .Z0_t (InputMUX_MUXInst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_9_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_9_U1_Y), .B0_t (Feedback[9]), .Z0_t (MCOutput[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_10_U1_XOR1_U1 ( .A0_t (Feedback[10]), .B0_t (Input[10]), .Z0_t (InputMUX_MUXInst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_10_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_10_U1_X), .Z0_t (InputMUX_MUXInst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_10_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_10_U1_Y), .B0_t (Feedback[10]), .Z0_t (MCOutput[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_11_U1_XOR1_U1 ( .A0_t (Feedback[11]), .B0_t (Input[11]), .Z0_t (InputMUX_MUXInst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_11_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_11_U1_X), .Z0_t (InputMUX_MUXInst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_11_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_11_U1_Y), .B0_t (Feedback[11]), .Z0_t (MCOutput[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_12_U1_XOR1_U1 ( .A0_t (Feedback[12]), .B0_t (Input[12]), .Z0_t (InputMUX_MUXInst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_12_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_12_U1_X), .Z0_t (InputMUX_MUXInst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_12_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_12_U1_Y), .B0_t (Feedback[12]), .Z0_t (MCOutput[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_13_U1_XOR1_U1 ( .A0_t (Feedback[13]), .B0_t (Input[13]), .Z0_t (InputMUX_MUXInst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_13_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_13_U1_X), .Z0_t (InputMUX_MUXInst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_13_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_13_U1_Y), .B0_t (Feedback[13]), .Z0_t (MCOutput[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_14_U1_XOR1_U1 ( .A0_t (Feedback[14]), .B0_t (Input[14]), .Z0_t (InputMUX_MUXInst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_14_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_14_U1_X), .Z0_t (InputMUX_MUXInst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_14_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_14_U1_Y), .B0_t (Feedback[14]), .Z0_t (MCOutput[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_15_U1_XOR1_U1 ( .A0_t (Feedback[15]), .B0_t (Input[15]), .Z0_t (InputMUX_MUXInst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_15_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_15_U1_X), .Z0_t (InputMUX_MUXInst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_15_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_15_U1_Y), .B0_t (Feedback[15]), .Z0_t (MCOutput[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_16_U1_XOR1_U1 ( .A0_t (Feedback[16]), .B0_t (Input[16]), .Z0_t (InputMUX_MUXInst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_16_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_16_U1_X), .Z0_t (InputMUX_MUXInst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_16_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_16_U1_Y), .B0_t (Feedback[16]), .Z0_t (MCOutput[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_17_U1_XOR1_U1 ( .A0_t (Feedback[17]), .B0_t (Input[17]), .Z0_t (InputMUX_MUXInst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_17_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_17_U1_X), .Z0_t (InputMUX_MUXInst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_17_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_17_U1_Y), .B0_t (Feedback[17]), .Z0_t (MCOutput[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_18_U1_XOR1_U1 ( .A0_t (Feedback[18]), .B0_t (Input[18]), .Z0_t (InputMUX_MUXInst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_18_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_18_U1_X), .Z0_t (InputMUX_MUXInst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_18_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_18_U1_Y), .B0_t (Feedback[18]), .Z0_t (MCOutput[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_19_U1_XOR1_U1 ( .A0_t (Feedback[19]), .B0_t (Input[19]), .Z0_t (InputMUX_MUXInst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_19_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_19_U1_X), .Z0_t (InputMUX_MUXInst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_19_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_19_U1_Y), .B0_t (Feedback[19]), .Z0_t (MCOutput[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_20_U1_XOR1_U1 ( .A0_t (Feedback[20]), .B0_t (Input[20]), .Z0_t (InputMUX_MUXInst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_20_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_20_U1_X), .Z0_t (InputMUX_MUXInst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_20_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_20_U1_Y), .B0_t (Feedback[20]), .Z0_t (MCOutput[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_21_U1_XOR1_U1 ( .A0_t (Feedback[21]), .B0_t (Input[21]), .Z0_t (InputMUX_MUXInst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_21_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_21_U1_X), .Z0_t (InputMUX_MUXInst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_21_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_21_U1_Y), .B0_t (Feedback[21]), .Z0_t (MCOutput[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_22_U1_XOR1_U1 ( .A0_t (Feedback[22]), .B0_t (Input[22]), .Z0_t (InputMUX_MUXInst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_22_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_22_U1_X), .Z0_t (InputMUX_MUXInst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_22_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_22_U1_Y), .B0_t (Feedback[22]), .Z0_t (MCOutput[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_23_U1_XOR1_U1 ( .A0_t (Feedback[23]), .B0_t (Input[23]), .Z0_t (InputMUX_MUXInst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_23_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_23_U1_X), .Z0_t (InputMUX_MUXInst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_23_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_23_U1_Y), .B0_t (Feedback[23]), .Z0_t (MCOutput[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_24_U1_XOR1_U1 ( .A0_t (Feedback[24]), .B0_t (Input[24]), .Z0_t (InputMUX_MUXInst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_24_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_24_U1_X), .Z0_t (InputMUX_MUXInst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_24_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_24_U1_Y), .B0_t (Feedback[24]), .Z0_t (MCOutput[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_25_U1_XOR1_U1 ( .A0_t (Feedback[25]), .B0_t (Input[25]), .Z0_t (InputMUX_MUXInst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_25_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_25_U1_X), .Z0_t (InputMUX_MUXInst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_25_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_25_U1_Y), .B0_t (Feedback[25]), .Z0_t (MCOutput[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_26_U1_XOR1_U1 ( .A0_t (Feedback[26]), .B0_t (Input[26]), .Z0_t (InputMUX_MUXInst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_26_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_26_U1_X), .Z0_t (InputMUX_MUXInst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_26_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_26_U1_Y), .B0_t (Feedback[26]), .Z0_t (MCOutput[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_27_U1_XOR1_U1 ( .A0_t (Feedback[27]), .B0_t (Input[27]), .Z0_t (InputMUX_MUXInst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_27_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_27_U1_X), .Z0_t (InputMUX_MUXInst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_27_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_27_U1_Y), .B0_t (Feedback[27]), .Z0_t (MCOutput[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_28_U1_XOR1_U1 ( .A0_t (Feedback[28]), .B0_t (Input[28]), .Z0_t (InputMUX_MUXInst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_28_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_28_U1_X), .Z0_t (InputMUX_MUXInst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_28_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_28_U1_Y), .B0_t (Feedback[28]), .Z0_t (MCOutput[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_29_U1_XOR1_U1 ( .A0_t (Feedback[29]), .B0_t (Input[29]), .Z0_t (InputMUX_MUXInst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_29_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_29_U1_X), .Z0_t (InputMUX_MUXInst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_29_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_29_U1_Y), .B0_t (Feedback[29]), .Z0_t (MCOutput[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_30_U1_XOR1_U1 ( .A0_t (Feedback[30]), .B0_t (Input[30]), .Z0_t (InputMUX_MUXInst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_30_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_30_U1_X), .Z0_t (InputMUX_MUXInst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_30_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_30_U1_Y), .B0_t (Feedback[30]), .Z0_t (MCOutput[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_31_U1_XOR1_U1 ( .A0_t (Feedback[31]), .B0_t (Input[31]), .Z0_t (InputMUX_MUXInst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_31_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_31_U1_X), .Z0_t (InputMUX_MUXInst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_31_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_31_U1_Y), .B0_t (Feedback[31]), .Z0_t (MCOutput[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_32_U1_XOR1_U1 ( .A0_t (Feedback[32]), .B0_t (Input[32]), .Z0_t (InputMUX_MUXInst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_32_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_32_U1_X), .Z0_t (InputMUX_MUXInst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_32_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_32_U1_Y), .B0_t (Feedback[32]), .Z0_t (MCInput[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_33_U1_XOR1_U1 ( .A0_t (Feedback[33]), .B0_t (Input[33]), .Z0_t (InputMUX_MUXInst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_33_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_33_U1_X), .Z0_t (InputMUX_MUXInst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_33_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_33_U1_Y), .B0_t (Feedback[33]), .Z0_t (MCInput[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_34_U1_XOR1_U1 ( .A0_t (Feedback[34]), .B0_t (Input[34]), .Z0_t (InputMUX_MUXInst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_34_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_34_U1_X), .Z0_t (InputMUX_MUXInst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_34_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_34_U1_Y), .B0_t (Feedback[34]), .Z0_t (MCInput[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_35_U1_XOR1_U1 ( .A0_t (Feedback[35]), .B0_t (Input[35]), .Z0_t (InputMUX_MUXInst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_35_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_35_U1_X), .Z0_t (InputMUX_MUXInst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_35_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_35_U1_Y), .B0_t (Feedback[35]), .Z0_t (MCInput[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_36_U1_XOR1_U1 ( .A0_t (Feedback[36]), .B0_t (Input[36]), .Z0_t (InputMUX_MUXInst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_36_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_36_U1_X), .Z0_t (InputMUX_MUXInst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_36_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_36_U1_Y), .B0_t (Feedback[36]), .Z0_t (MCInput[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_37_U1_XOR1_U1 ( .A0_t (Feedback[37]), .B0_t (Input[37]), .Z0_t (InputMUX_MUXInst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_37_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_37_U1_X), .Z0_t (InputMUX_MUXInst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_37_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_37_U1_Y), .B0_t (Feedback[37]), .Z0_t (MCInput[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_38_U1_XOR1_U1 ( .A0_t (Feedback[38]), .B0_t (Input[38]), .Z0_t (InputMUX_MUXInst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_38_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_38_U1_X), .Z0_t (InputMUX_MUXInst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_38_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_38_U1_Y), .B0_t (Feedback[38]), .Z0_t (MCInput[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_39_U1_XOR1_U1 ( .A0_t (Feedback[39]), .B0_t (Input[39]), .Z0_t (InputMUX_MUXInst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_39_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_39_U1_X), .Z0_t (InputMUX_MUXInst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_39_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_39_U1_Y), .B0_t (Feedback[39]), .Z0_t (MCInput[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_40_U1_XOR1_U1 ( .A0_t (Feedback[40]), .B0_t (Input[40]), .Z0_t (InputMUX_MUXInst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_40_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_40_U1_X), .Z0_t (InputMUX_MUXInst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_40_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_40_U1_Y), .B0_t (Feedback[40]), .Z0_t (MCInput[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_41_U1_XOR1_U1 ( .A0_t (Feedback[41]), .B0_t (Input[41]), .Z0_t (InputMUX_MUXInst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_41_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_41_U1_X), .Z0_t (InputMUX_MUXInst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_41_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_41_U1_Y), .B0_t (Feedback[41]), .Z0_t (MCInput[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_42_U1_XOR1_U1 ( .A0_t (Feedback[42]), .B0_t (Input[42]), .Z0_t (InputMUX_MUXInst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_42_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_42_U1_X), .Z0_t (InputMUX_MUXInst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_42_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_42_U1_Y), .B0_t (Feedback[42]), .Z0_t (MCInput[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_43_U1_XOR1_U1 ( .A0_t (Feedback[43]), .B0_t (Input[43]), .Z0_t (InputMUX_MUXInst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_43_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_43_U1_X), .Z0_t (InputMUX_MUXInst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_43_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_43_U1_Y), .B0_t (Feedback[43]), .Z0_t (MCInput[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_44_U1_XOR1_U1 ( .A0_t (Feedback[44]), .B0_t (Input[44]), .Z0_t (InputMUX_MUXInst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_44_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_44_U1_X), .Z0_t (InputMUX_MUXInst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_44_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_44_U1_Y), .B0_t (Feedback[44]), .Z0_t (MCInput[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_45_U1_XOR1_U1 ( .A0_t (Feedback[45]), .B0_t (Input[45]), .Z0_t (InputMUX_MUXInst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_45_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_45_U1_X), .Z0_t (InputMUX_MUXInst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_45_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_45_U1_Y), .B0_t (Feedback[45]), .Z0_t (MCInput[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_46_U1_XOR1_U1 ( .A0_t (Feedback[46]), .B0_t (Input[46]), .Z0_t (InputMUX_MUXInst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_46_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_46_U1_X), .Z0_t (InputMUX_MUXInst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_46_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_46_U1_Y), .B0_t (Feedback[46]), .Z0_t (MCInput[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_47_U1_XOR1_U1 ( .A0_t (Feedback[47]), .B0_t (Input[47]), .Z0_t (InputMUX_MUXInst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_47_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_47_U1_X), .Z0_t (InputMUX_MUXInst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_47_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_47_U1_Y), .B0_t (Feedback[47]), .Z0_t (MCInput[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_48_U1_XOR1_U1 ( .A0_t (Feedback[48]), .B0_t (Input[48]), .Z0_t (InputMUX_MUXInst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_48_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_48_U1_X), .Z0_t (InputMUX_MUXInst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_48_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_48_U1_Y), .B0_t (Feedback[48]), .Z0_t (MCInput[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_49_U1_XOR1_U1 ( .A0_t (Feedback[49]), .B0_t (Input[49]), .Z0_t (InputMUX_MUXInst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_49_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_49_U1_X), .Z0_t (InputMUX_MUXInst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_49_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_49_U1_Y), .B0_t (Feedback[49]), .Z0_t (MCInput[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_50_U1_XOR1_U1 ( .A0_t (Feedback[50]), .B0_t (Input[50]), .Z0_t (InputMUX_MUXInst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_50_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_50_U1_X), .Z0_t (InputMUX_MUXInst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_50_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_50_U1_Y), .B0_t (Feedback[50]), .Z0_t (MCInput[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_51_U1_XOR1_U1 ( .A0_t (Feedback[51]), .B0_t (Input[51]), .Z0_t (InputMUX_MUXInst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_51_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_51_U1_X), .Z0_t (InputMUX_MUXInst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_51_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_51_U1_Y), .B0_t (Feedback[51]), .Z0_t (MCInput[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_52_U1_XOR1_U1 ( .A0_t (Feedback[52]), .B0_t (Input[52]), .Z0_t (InputMUX_MUXInst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_52_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_52_U1_X), .Z0_t (InputMUX_MUXInst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_52_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_52_U1_Y), .B0_t (Feedback[52]), .Z0_t (MCInput[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_53_U1_XOR1_U1 ( .A0_t (Feedback[53]), .B0_t (Input[53]), .Z0_t (InputMUX_MUXInst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_53_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_53_U1_X), .Z0_t (InputMUX_MUXInst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_53_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_53_U1_Y), .B0_t (Feedback[53]), .Z0_t (MCInput[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_54_U1_XOR1_U1 ( .A0_t (Feedback[54]), .B0_t (Input[54]), .Z0_t (InputMUX_MUXInst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_54_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_54_U1_X), .Z0_t (InputMUX_MUXInst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_54_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_54_U1_Y), .B0_t (Feedback[54]), .Z0_t (MCInput[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_55_U1_XOR1_U1 ( .A0_t (Feedback[55]), .B0_t (Input[55]), .Z0_t (InputMUX_MUXInst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_55_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_55_U1_X), .Z0_t (InputMUX_MUXInst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_55_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_55_U1_Y), .B0_t (Feedback[55]), .Z0_t (MCInput[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_56_U1_XOR1_U1 ( .A0_t (Feedback[56]), .B0_t (Input[56]), .Z0_t (InputMUX_MUXInst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_56_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_56_U1_X), .Z0_t (InputMUX_MUXInst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_56_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_56_U1_Y), .B0_t (Feedback[56]), .Z0_t (MCInput[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_57_U1_XOR1_U1 ( .A0_t (Feedback[57]), .B0_t (Input[57]), .Z0_t (InputMUX_MUXInst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_57_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_57_U1_X), .Z0_t (InputMUX_MUXInst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_57_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_57_U1_Y), .B0_t (Feedback[57]), .Z0_t (MCInput[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_58_U1_XOR1_U1 ( .A0_t (Feedback[58]), .B0_t (Input[58]), .Z0_t (InputMUX_MUXInst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_58_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_58_U1_X), .Z0_t (InputMUX_MUXInst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_58_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_58_U1_Y), .B0_t (Feedback[58]), .Z0_t (MCInput[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_59_U1_XOR1_U1 ( .A0_t (Feedback[59]), .B0_t (Input[59]), .Z0_t (InputMUX_MUXInst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_59_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_59_U1_X), .Z0_t (InputMUX_MUXInst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_59_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_59_U1_Y), .B0_t (Feedback[59]), .Z0_t (MCInput[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_60_U1_XOR1_U1 ( .A0_t (Feedback[60]), .B0_t (Input[60]), .Z0_t (InputMUX_MUXInst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_60_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_60_U1_X), .Z0_t (InputMUX_MUXInst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_60_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_60_U1_Y), .B0_t (Feedback[60]), .Z0_t (MCInput[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_61_U1_XOR1_U1 ( .A0_t (Feedback[61]), .B0_t (Input[61]), .Z0_t (InputMUX_MUXInst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_61_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_61_U1_X), .Z0_t (InputMUX_MUXInst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_61_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_61_U1_Y), .B0_t (Feedback[61]), .Z0_t (MCInput[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_62_U1_XOR1_U1 ( .A0_t (Feedback[62]), .B0_t (Input[62]), .Z0_t (InputMUX_MUXInst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_62_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_62_U1_X), .Z0_t (InputMUX_MUXInst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_62_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_62_U1_Y), .B0_t (Feedback[62]), .Z0_t (MCInput[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_63_U1_XOR1_U1 ( .A0_t (Feedback[63]), .B0_t (Input[63]), .Z0_t (InputMUX_MUXInst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_63_U1_AND1_U1 ( .A0_t (rst), .B0_t (InputMUX_MUXInst_63_U1_X), .Z0_t (InputMUX_MUXInst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_63_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_63_U1_Y), .B0_t (Feedback[63]), .Z0_t (MCInput[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_0_U2 ( .A0_t (MCInst_XOR_r0_Inst_0_n1), .B0_t (MCOutput[0]), .Z0_t (MCOutput[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_0_U1 ( .A0_t (MCInput[48]), .B0_t (MCOutput[16]), .Z0_t (MCInst_XOR_r0_Inst_0_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_0_U1 ( .A0_t (MCInput[32]), .B0_t (MCOutput[0]), .Z0_t (MCOutput[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_1_U2 ( .A0_t (MCInst_XOR_r0_Inst_1_n1), .B0_t (MCOutput[1]), .Z0_t (MCOutput[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_1_U1 ( .A0_t (MCInput[49]), .B0_t (MCOutput[17]), .Z0_t (MCInst_XOR_r0_Inst_1_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_1_U1 ( .A0_t (MCInput[33]), .B0_t (MCOutput[1]), .Z0_t (MCOutput[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_2_U2 ( .A0_t (MCInst_XOR_r0_Inst_2_n1), .B0_t (MCOutput[2]), .Z0_t (MCOutput[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_2_U1 ( .A0_t (MCInput[50]), .B0_t (MCOutput[18]), .Z0_t (MCInst_XOR_r0_Inst_2_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_2_U1 ( .A0_t (MCInput[34]), .B0_t (MCOutput[2]), .Z0_t (MCOutput[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_3_U2 ( .A0_t (MCInst_XOR_r0_Inst_3_n1), .B0_t (MCOutput[3]), .Z0_t (MCOutput[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_3_U1 ( .A0_t (MCInput[51]), .B0_t (MCOutput[19]), .Z0_t (MCInst_XOR_r0_Inst_3_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_3_U1 ( .A0_t (MCInput[35]), .B0_t (MCOutput[3]), .Z0_t (MCOutput[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_4_U2 ( .A0_t (MCInst_XOR_r0_Inst_4_n1), .B0_t (MCOutput[4]), .Z0_t (MCOutput[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_4_U1 ( .A0_t (MCInput[52]), .B0_t (MCOutput[20]), .Z0_t (MCInst_XOR_r0_Inst_4_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_4_U1 ( .A0_t (MCInput[36]), .B0_t (MCOutput[4]), .Z0_t (MCOutput[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_5_U2 ( .A0_t (MCInst_XOR_r0_Inst_5_n1), .B0_t (MCOutput[5]), .Z0_t (MCOutput[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_5_U1 ( .A0_t (MCInput[53]), .B0_t (MCOutput[21]), .Z0_t (MCInst_XOR_r0_Inst_5_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_5_U1 ( .A0_t (MCInput[37]), .B0_t (MCOutput[5]), .Z0_t (MCOutput[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_6_U2 ( .A0_t (MCInst_XOR_r0_Inst_6_n1), .B0_t (MCOutput[6]), .Z0_t (MCOutput[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_6_U1 ( .A0_t (MCInput[54]), .B0_t (MCOutput[22]), .Z0_t (MCInst_XOR_r0_Inst_6_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_6_U1 ( .A0_t (MCInput[38]), .B0_t (MCOutput[6]), .Z0_t (MCOutput[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_7_U2 ( .A0_t (MCInst_XOR_r0_Inst_7_n1), .B0_t (MCOutput[7]), .Z0_t (MCOutput[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_7_U1 ( .A0_t (MCInput[55]), .B0_t (MCOutput[23]), .Z0_t (MCInst_XOR_r0_Inst_7_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_7_U1 ( .A0_t (MCInput[39]), .B0_t (MCOutput[7]), .Z0_t (MCOutput[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_8_U2 ( .A0_t (MCInst_XOR_r0_Inst_8_n1), .B0_t (MCOutput[8]), .Z0_t (MCOutput[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_8_U1 ( .A0_t (MCInput[56]), .B0_t (MCOutput[24]), .Z0_t (MCInst_XOR_r0_Inst_8_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_8_U1 ( .A0_t (MCInput[40]), .B0_t (MCOutput[8]), .Z0_t (MCOutput[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_9_U2 ( .A0_t (MCInst_XOR_r0_Inst_9_n1), .B0_t (MCOutput[9]), .Z0_t (MCOutput[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_9_U1 ( .A0_t (MCInput[57]), .B0_t (MCOutput[25]), .Z0_t (MCInst_XOR_r0_Inst_9_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_9_U1 ( .A0_t (MCInput[41]), .B0_t (MCOutput[9]), .Z0_t (MCOutput[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_10_U2 ( .A0_t (MCInst_XOR_r0_Inst_10_n1), .B0_t (MCOutput[10]), .Z0_t (MCOutput[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_10_U1 ( .A0_t (MCInput[58]), .B0_t (MCOutput[26]), .Z0_t (MCInst_XOR_r0_Inst_10_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_10_U1 ( .A0_t (MCInput[42]), .B0_t (MCOutput[10]), .Z0_t (MCOutput[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_11_U2 ( .A0_t (MCInst_XOR_r0_Inst_11_n1), .B0_t (MCOutput[11]), .Z0_t (MCOutput[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_11_U1 ( .A0_t (MCInput[59]), .B0_t (MCOutput[27]), .Z0_t (MCInst_XOR_r0_Inst_11_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_11_U1 ( .A0_t (MCInput[43]), .B0_t (MCOutput[11]), .Z0_t (MCOutput[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_12_U2 ( .A0_t (MCInst_XOR_r0_Inst_12_n1), .B0_t (MCOutput[12]), .Z0_t (MCOutput[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_12_U1 ( .A0_t (MCInput[60]), .B0_t (MCOutput[28]), .Z0_t (MCInst_XOR_r0_Inst_12_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_12_U1 ( .A0_t (MCInput[44]), .B0_t (MCOutput[12]), .Z0_t (MCOutput[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_13_U2 ( .A0_t (MCInst_XOR_r0_Inst_13_n1), .B0_t (MCOutput[13]), .Z0_t (MCOutput[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_13_U1 ( .A0_t (MCInput[61]), .B0_t (MCOutput[29]), .Z0_t (MCInst_XOR_r0_Inst_13_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_13_U1 ( .A0_t (MCInput[45]), .B0_t (MCOutput[13]), .Z0_t (MCOutput[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_14_U2 ( .A0_t (MCInst_XOR_r0_Inst_14_n1), .B0_t (MCOutput[14]), .Z0_t (MCOutput[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_14_U1 ( .A0_t (MCInput[62]), .B0_t (MCOutput[30]), .Z0_t (MCInst_XOR_r0_Inst_14_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_14_U1 ( .A0_t (MCInput[46]), .B0_t (MCOutput[14]), .Z0_t (MCOutput[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_15_U2 ( .A0_t (MCInst_XOR_r0_Inst_15_n1), .B0_t (MCOutput[15]), .Z0_t (MCOutput[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_15_U1 ( .A0_t (MCInput[63]), .B0_t (MCOutput[31]), .Z0_t (MCInst_XOR_r0_Inst_15_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_15_U1 ( .A0_t (MCInput[47]), .B0_t (MCOutput[15]), .Z0_t (MCOutput[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_0_0_U1 ( .A0_t (MCOutput[48]), .B0_t (SelectedKey[48]), .Z0_t (Output[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_0_1_U1 ( .A0_t (MCOutput[49]), .B0_t (SelectedKey[49]), .Z0_t (Output[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_0_2_U1 ( .A0_t (MCOutput[50]), .B0_t (SelectedKey[50]), .Z0_t (Output[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_0_3_U1 ( .A0_t (MCOutput[51]), .B0_t (SelectedKey[51]), .Z0_t (Output[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_1_0_U1 ( .A0_t (MCOutput[52]), .B0_t (SelectedKey[52]), .Z0_t (Output[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_1_1_U1 ( .A0_t (MCOutput[53]), .B0_t (SelectedKey[53]), .Z0_t (Output[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_1_2_U1 ( .A0_t (MCOutput[54]), .B0_t (SelectedKey[54]), .Z0_t (Output[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_1_3_U1 ( .A0_t (MCOutput[55]), .B0_t (SelectedKey[55]), .Z0_t (Output[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_2_0_U1 ( .A0_t (MCOutput[56]), .B0_t (SelectedKey[56]), .Z0_t (Output[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_2_1_U1 ( .A0_t (MCOutput[57]), .B0_t (SelectedKey[57]), .Z0_t (Output[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_2_2_U1 ( .A0_t (MCOutput[58]), .B0_t (SelectedKey[58]), .Z0_t (Output[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_2_3_U1 ( .A0_t (MCOutput[59]), .B0_t (SelectedKey[59]), .Z0_t (Output[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_3_0_U1 ( .A0_t (MCOutput[60]), .B0_t (SelectedKey[60]), .Z0_t (Output[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_3_1_U1 ( .A0_t (MCOutput[61]), .B0_t (SelectedKey[61]), .Z0_t (Output[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_3_2_U1 ( .A0_t (MCOutput[62]), .B0_t (SelectedKey[62]), .Z0_t (Output[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_3_3_U1 ( .A0_t (MCOutput[63]), .B0_t (SelectedKey[63]), .Z0_t (Output[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_0_0_U2 ( .A0_t (AddKeyConstXOR_XORInst_0_0_n1), .B0_t (SelectedKey[40]), .Z0_t (Output[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_0_0_U1 ( .A0_t (RoundConstant_0), .B0_t (MCOutput[40]), .Z0_t (AddKeyConstXOR_XORInst_0_0_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_0_1_U2 ( .A0_t (AddKeyConstXOR_XORInst_0_1_n1), .B0_t (SelectedKey[41]), .Z0_t (Output[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_0_1_U1 ( .A0_t (FSMUpdate[0]), .B0_t (MCOutput[41]), .Z0_t (AddKeyConstXOR_XORInst_0_1_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_0_2_U2 ( .A0_t (AddKeyConstXOR_XORInst_0_2_n1), .B0_t (SelectedKey[42]), .Z0_t (Output[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_0_2_U1 ( .A0_t (FSMUpdate[1]), .B0_t (MCOutput[42]), .Z0_t (AddKeyConstXOR_XORInst_0_2_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyConstXOR_XORInst_0_3_U1 ( .A0_t (MCOutput[43]), .B0_t (SelectedKey[43]), .Z0_t (Output[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_1_0_U2 ( .A0_t (AddKeyConstXOR_XORInst_1_0_n1), .B0_t (SelectedKey[44]), .Z0_t (Output[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_1_0_U1 ( .A0_t (RoundConstant_4_), .B0_t (MCOutput[44]), .Z0_t (AddKeyConstXOR_XORInst_1_0_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_1_1_U2 ( .A0_t (AddKeyConstXOR_XORInst_1_1_n1), .B0_t (SelectedKey[45]), .Z0_t (Output[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_1_1_U1 ( .A0_t (FSMUpdate[3]), .B0_t (MCOutput[45]), .Z0_t (AddKeyConstXOR_XORInst_1_1_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_1_2_U2 ( .A0_t (AddKeyConstXOR_XORInst_1_2_n1), .B0_t (SelectedKey[46]), .Z0_t (Output[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_1_2_U1 ( .A0_t (FSMUpdate[4]), .B0_t (MCOutput[46]), .Z0_t (AddKeyConstXOR_XORInst_1_2_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_1_3_U2 ( .A0_t (AddKeyConstXOR_XORInst_1_3_n1), .B0_t (SelectedKey[47]), .Z0_t (Output[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_1_3_U1 ( .A0_t (FSMUpdate[5]), .B0_t (MCOutput[47]), .Z0_t (AddKeyConstXOR_XORInst_1_3_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_0_0_U1 ( .A0_t (MCOutput[0]), .B0_t (SelectedKey[0]), .Z0_t (Output[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_0_1_U1 ( .A0_t (MCOutput[1]), .B0_t (SelectedKey[1]), .Z0_t (Output[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_0_2_U1 ( .A0_t (MCOutput[2]), .B0_t (SelectedKey[2]), .Z0_t (Output[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_0_3_U1 ( .A0_t (MCOutput[3]), .B0_t (SelectedKey[3]), .Z0_t (Output[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_1_0_U1 ( .A0_t (MCOutput[4]), .B0_t (SelectedKey[4]), .Z0_t (Output[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_1_1_U1 ( .A0_t (MCOutput[5]), .B0_t (SelectedKey[5]), .Z0_t (Output[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_1_2_U1 ( .A0_t (MCOutput[6]), .B0_t (SelectedKey[6]), .Z0_t (Output[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_1_3_U1 ( .A0_t (MCOutput[7]), .B0_t (SelectedKey[7]), .Z0_t (Output[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_2_0_U1 ( .A0_t (MCOutput[8]), .B0_t (SelectedKey[8]), .Z0_t (Output[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_2_1_U1 ( .A0_t (MCOutput[9]), .B0_t (SelectedKey[9]), .Z0_t (Output[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_2_2_U1 ( .A0_t (MCOutput[10]), .B0_t (SelectedKey[10]), .Z0_t (Output[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_2_3_U1 ( .A0_t (MCOutput[11]), .B0_t (SelectedKey[11]), .Z0_t (Output[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_3_0_U1 ( .A0_t (MCOutput[12]), .B0_t (SelectedKey[12]), .Z0_t (Output[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_3_1_U1 ( .A0_t (MCOutput[13]), .B0_t (SelectedKey[13]), .Z0_t (Output[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_3_2_U1 ( .A0_t (MCOutput[14]), .B0_t (SelectedKey[14]), .Z0_t (Output[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_3_3_U1 ( .A0_t (MCOutput[15]), .B0_t (SelectedKey[15]), .Z0_t (Output[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_4_0_U1 ( .A0_t (MCOutput[16]), .B0_t (SelectedKey[16]), .Z0_t (Output[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_4_1_U1 ( .A0_t (MCOutput[17]), .B0_t (SelectedKey[17]), .Z0_t (Output[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_4_2_U1 ( .A0_t (MCOutput[18]), .B0_t (SelectedKey[18]), .Z0_t (Output[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_4_3_U1 ( .A0_t (MCOutput[19]), .B0_t (SelectedKey[19]), .Z0_t (Output[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_5_0_U1 ( .A0_t (MCOutput[20]), .B0_t (SelectedKey[20]), .Z0_t (Output[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_5_1_U1 ( .A0_t (MCOutput[21]), .B0_t (SelectedKey[21]), .Z0_t (Output[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_5_2_U1 ( .A0_t (MCOutput[22]), .B0_t (SelectedKey[22]), .Z0_t (Output[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_5_3_U1 ( .A0_t (MCOutput[23]), .B0_t (SelectedKey[23]), .Z0_t (Output[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_6_0_U1 ( .A0_t (MCOutput[24]), .B0_t (SelectedKey[24]), .Z0_t (Output[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_6_1_U1 ( .A0_t (MCOutput[25]), .B0_t (SelectedKey[25]), .Z0_t (Output[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_6_2_U1 ( .A0_t (MCOutput[26]), .B0_t (SelectedKey[26]), .Z0_t (Output[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_6_3_U1 ( .A0_t (MCOutput[27]), .B0_t (SelectedKey[27]), .Z0_t (Output[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_7_0_U1 ( .A0_t (MCOutput[28]), .B0_t (SelectedKey[28]), .Z0_t (Output[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_7_1_U1 ( .A0_t (MCOutput[29]), .B0_t (SelectedKey[29]), .Z0_t (Output[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_7_2_U1 ( .A0_t (MCOutput[30]), .B0_t (SelectedKey[30]), .Z0_t (Output[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_7_3_U1 ( .A0_t (MCOutput[31]), .B0_t (SelectedKey[31]), .Z0_t (Output[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_8_0_U1 ( .A0_t (MCOutput[32]), .B0_t (SelectedKey[32]), .Z0_t (Output[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_8_1_U1 ( .A0_t (MCOutput[33]), .B0_t (SelectedKey[33]), .Z0_t (Output[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_8_2_U1 ( .A0_t (MCOutput[34]), .B0_t (SelectedKey[34]), .Z0_t (Output[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_8_3_U1 ( .A0_t (MCOutput[35]), .B0_t (SelectedKey[35]), .Z0_t (Output[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_9_0_U1 ( .A0_t (MCOutput[36]), .B0_t (SelectedKey[36]), .Z0_t (Output[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_9_1_U1 ( .A0_t (MCOutput[37]), .B0_t (SelectedKey[37]), .Z0_t (Output[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_9_2_U1 ( .A0_t (MCOutput[38]), .B0_t (SelectedKey[38]), .Z0_t (Output[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_9_3_U1 ( .A0_t (MCOutput[39]), .B0_t (SelectedKey[39]), .Z0_t (Output[39]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_U19 ( .A0_t (SubCellInst_SboxInst_0_n15), .B0_t (SubCellInst_SboxInst_0_n14), .Z0_t (Feedback[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_U18 ( .A0_t (Output[61]), .B0_t (SubCellInst_SboxInst_0_n13), .Z0_t (SubCellInst_SboxInst_0_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_U17 ( .A0_t (Output[60]), .B0_t (SubCellInst_SboxInst_0_n11), .Z0_t (SubCellInst_SboxInst_0_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_U16 ( .A0_t (Output[62]), .B0_t (Output[63]), .Z0_t (SubCellInst_SboxInst_0_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U15 ( .A0_t (SubCellInst_SboxInst_0_n10), .B0_t (SubCellInst_SboxInst_0_n9), .Z0_t (Feedback[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U14 ( .A0_t (Output[60]), .B0_t (Output[63]), .Z0_t (SubCellInst_SboxInst_0_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U13 ( .A0_t (Output[62]), .B0_t (SubCellInst_SboxInst_0_n7), .Z0_t (SubCellInst_SboxInst_0_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U12 ( .A0_t (Output[63]), .B0_t (Output[60]), .Z0_t (SubCellInst_SboxInst_0_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U11 ( .A0_t (SubCellInst_SboxInst_0_n6), .B0_t (SubCellInst_SboxInst_0_n5), .Z0_t (Feedback[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U10 ( .A0_t (SubCellInst_SboxInst_0_n4), .B0_t (Output[61]), .Z0_t (SubCellInst_SboxInst_0_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U9 ( .A0_t (SubCellInst_SboxInst_0_n3), .B0_t (Output[62]), .Z0_t (SubCellInst_SboxInst_0_n4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U8 ( .A0_t (Output[60]), .B0_t (Output[63]), .Z0_t (SubCellInst_SboxInst_0_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U7 ( .A0_t (SubCellInst_SboxInst_0_n5), .B0_t (SubCellInst_SboxInst_0_n1), .Z0_t (Feedback[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U6 ( .A0_t (Output[61]), .B0_t (SubCellInst_SboxInst_0_n14), .Z0_t (SubCellInst_SboxInst_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_U5 ( .A0_t (Output[62]), .B0_t (Output[63]), .Z0_t (SubCellInst_SboxInst_0_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U3 ( .A0_t (Output[63]), .B0_t (Output[60]), .Z0_t (SubCellInst_SboxInst_0_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_U19 ( .A0_t (SubCellInst_SboxInst_1_n15), .B0_t (SubCellInst_SboxInst_1_n14), .Z0_t (Feedback[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_U18 ( .A0_t (Output[49]), .B0_t (SubCellInst_SboxInst_1_n13), .Z0_t (SubCellInst_SboxInst_1_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_U17 ( .A0_t (Output[48]), .B0_t (SubCellInst_SboxInst_1_n11), .Z0_t (SubCellInst_SboxInst_1_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_U16 ( .A0_t (Output[50]), .B0_t (Output[51]), .Z0_t (SubCellInst_SboxInst_1_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U15 ( .A0_t (SubCellInst_SboxInst_1_n10), .B0_t (SubCellInst_SboxInst_1_n9), .Z0_t (Feedback[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U14 ( .A0_t (Output[48]), .B0_t (Output[51]), .Z0_t (SubCellInst_SboxInst_1_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U13 ( .A0_t (Output[50]), .B0_t (SubCellInst_SboxInst_1_n7), .Z0_t (SubCellInst_SboxInst_1_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U12 ( .A0_t (Output[51]), .B0_t (Output[48]), .Z0_t (SubCellInst_SboxInst_1_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U11 ( .A0_t (SubCellInst_SboxInst_1_n6), .B0_t (SubCellInst_SboxInst_1_n5), .Z0_t (Feedback[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U10 ( .A0_t (SubCellInst_SboxInst_1_n4), .B0_t (Output[49]), .Z0_t (SubCellInst_SboxInst_1_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U9 ( .A0_t (SubCellInst_SboxInst_1_n3), .B0_t (Output[50]), .Z0_t (SubCellInst_SboxInst_1_n4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U8 ( .A0_t (Output[48]), .B0_t (Output[51]), .Z0_t (SubCellInst_SboxInst_1_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U7 ( .A0_t (SubCellInst_SboxInst_1_n5), .B0_t (SubCellInst_SboxInst_1_n1), .Z0_t (Feedback[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U6 ( .A0_t (Output[49]), .B0_t (SubCellInst_SboxInst_1_n14), .Z0_t (SubCellInst_SboxInst_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_U5 ( .A0_t (Output[50]), .B0_t (Output[51]), .Z0_t (SubCellInst_SboxInst_1_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U3 ( .A0_t (Output[51]), .B0_t (Output[48]), .Z0_t (SubCellInst_SboxInst_1_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_U19 ( .A0_t (SubCellInst_SboxInst_2_n15), .B0_t (SubCellInst_SboxInst_2_n14), .Z0_t (Feedback[8]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_U18 ( .A0_t (Output[53]), .B0_t (SubCellInst_SboxInst_2_n13), .Z0_t (SubCellInst_SboxInst_2_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_U17 ( .A0_t (Output[52]), .B0_t (SubCellInst_SboxInst_2_n11), .Z0_t (SubCellInst_SboxInst_2_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_U16 ( .A0_t (Output[54]), .B0_t (Output[55]), .Z0_t (SubCellInst_SboxInst_2_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U15 ( .A0_t (SubCellInst_SboxInst_2_n10), .B0_t (SubCellInst_SboxInst_2_n9), .Z0_t (Feedback[9]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U14 ( .A0_t (Output[52]), .B0_t (Output[55]), .Z0_t (SubCellInst_SboxInst_2_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U13 ( .A0_t (Output[54]), .B0_t (SubCellInst_SboxInst_2_n7), .Z0_t (SubCellInst_SboxInst_2_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U12 ( .A0_t (Output[55]), .B0_t (Output[52]), .Z0_t (SubCellInst_SboxInst_2_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U11 ( .A0_t (SubCellInst_SboxInst_2_n6), .B0_t (SubCellInst_SboxInst_2_n5), .Z0_t (Feedback[10]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U10 ( .A0_t (SubCellInst_SboxInst_2_n4), .B0_t (Output[53]), .Z0_t (SubCellInst_SboxInst_2_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U9 ( .A0_t (SubCellInst_SboxInst_2_n3), .B0_t (Output[54]), .Z0_t (SubCellInst_SboxInst_2_n4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U8 ( .A0_t (Output[52]), .B0_t (Output[55]), .Z0_t (SubCellInst_SboxInst_2_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U7 ( .A0_t (SubCellInst_SboxInst_2_n5), .B0_t (SubCellInst_SboxInst_2_n1), .Z0_t (Feedback[11]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U6 ( .A0_t (Output[53]), .B0_t (SubCellInst_SboxInst_2_n14), .Z0_t (SubCellInst_SboxInst_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_U5 ( .A0_t (Output[54]), .B0_t (Output[55]), .Z0_t (SubCellInst_SboxInst_2_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U3 ( .A0_t (Output[55]), .B0_t (Output[52]), .Z0_t (SubCellInst_SboxInst_2_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_U19 ( .A0_t (SubCellInst_SboxInst_3_n15), .B0_t (SubCellInst_SboxInst_3_n14), .Z0_t (Feedback[12]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_U18 ( .A0_t (Output[57]), .B0_t (SubCellInst_SboxInst_3_n13), .Z0_t (SubCellInst_SboxInst_3_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_U17 ( .A0_t (Output[56]), .B0_t (SubCellInst_SboxInst_3_n11), .Z0_t (SubCellInst_SboxInst_3_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_U16 ( .A0_t (Output[58]), .B0_t (Output[59]), .Z0_t (SubCellInst_SboxInst_3_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U15 ( .A0_t (SubCellInst_SboxInst_3_n10), .B0_t (SubCellInst_SboxInst_3_n9), .Z0_t (Feedback[13]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U14 ( .A0_t (Output[56]), .B0_t (Output[59]), .Z0_t (SubCellInst_SboxInst_3_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U13 ( .A0_t (Output[58]), .B0_t (SubCellInst_SboxInst_3_n7), .Z0_t (SubCellInst_SboxInst_3_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U12 ( .A0_t (Output[59]), .B0_t (Output[56]), .Z0_t (SubCellInst_SboxInst_3_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U11 ( .A0_t (SubCellInst_SboxInst_3_n6), .B0_t (SubCellInst_SboxInst_3_n5), .Z0_t (Feedback[14]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U10 ( .A0_t (SubCellInst_SboxInst_3_n4), .B0_t (Output[57]), .Z0_t (SubCellInst_SboxInst_3_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U9 ( .A0_t (SubCellInst_SboxInst_3_n3), .B0_t (Output[58]), .Z0_t (SubCellInst_SboxInst_3_n4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U8 ( .A0_t (Output[56]), .B0_t (Output[59]), .Z0_t (SubCellInst_SboxInst_3_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U7 ( .A0_t (SubCellInst_SboxInst_3_n5), .B0_t (SubCellInst_SboxInst_3_n1), .Z0_t (Feedback[15]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U6 ( .A0_t (Output[57]), .B0_t (SubCellInst_SboxInst_3_n14), .Z0_t (SubCellInst_SboxInst_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_U5 ( .A0_t (Output[58]), .B0_t (Output[59]), .Z0_t (SubCellInst_SboxInst_3_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U3 ( .A0_t (Output[59]), .B0_t (Output[56]), .Z0_t (SubCellInst_SboxInst_3_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U19 ( .A0_t (SubCellInst_SboxInst_4_n15), .B0_t (SubCellInst_SboxInst_4_n14), .Z0_t (Feedback[17]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U18 ( .A0_t (Output[34]), .B0_t (SubCellInst_SboxInst_4_n13), .Z0_t (SubCellInst_SboxInst_4_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U17 ( .A0_t (Output[35]), .B0_t (Output[32]), .Z0_t (SubCellInst_SboxInst_4_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U16 ( .A0_t (Output[32]), .B0_t (Output[35]), .Z0_t (SubCellInst_SboxInst_4_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U15 ( .A0_t (SubCellInst_SboxInst_4_n10), .B0_t (SubCellInst_SboxInst_4_n9), .Z0_t (Feedback[19]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U14 ( .A0_t (Output[33]), .B0_t (SubCellInst_SboxInst_4_n8), .Z0_t (SubCellInst_SboxInst_4_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_U13 ( .A0_t (SubCellInst_SboxInst_4_n8), .B0_t (SubCellInst_SboxInst_4_n7), .Z0_t (Feedback[16]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_U12 ( .A0_t (Output[33]), .B0_t (SubCellInst_SboxInst_4_n6), .Z0_t (SubCellInst_SboxInst_4_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_U11 ( .A0_t (Output[32]), .B0_t (SubCellInst_SboxInst_4_n5), .Z0_t (SubCellInst_SboxInst_4_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_U10 ( .A0_t (Output[35]), .B0_t (Output[34]), .Z0_t (SubCellInst_SboxInst_4_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_U9 ( .A0_t (Output[35]), .B0_t (Output[34]), .Z0_t (SubCellInst_SboxInst_4_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U8 ( .A0_t (SubCellInst_SboxInst_4_n10), .B0_t (SubCellInst_SboxInst_4_n3), .Z0_t (Feedback[18]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U7 ( .A0_t (SubCellInst_SboxInst_4_n2), .B0_t (Output[33]), .Z0_t (SubCellInst_SboxInst_4_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U6 ( .A0_t (SubCellInst_SboxInst_4_n1), .B0_t (Output[34]), .Z0_t (SubCellInst_SboxInst_4_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U4 ( .A0_t (Output[35]), .B0_t (Output[32]), .Z0_t (SubCellInst_SboxInst_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U3 ( .A0_t (Output[32]), .B0_t (Output[35]), .Z0_t (SubCellInst_SboxInst_4_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U19 ( .A0_t (SubCellInst_SboxInst_5_n15), .B0_t (SubCellInst_SboxInst_5_n14), .Z0_t (Feedback[21]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U18 ( .A0_t (Output[46]), .B0_t (SubCellInst_SboxInst_5_n13), .Z0_t (SubCellInst_SboxInst_5_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U17 ( .A0_t (Output[47]), .B0_t (Output[44]), .Z0_t (SubCellInst_SboxInst_5_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U16 ( .A0_t (Output[44]), .B0_t (Output[47]), .Z0_t (SubCellInst_SboxInst_5_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U15 ( .A0_t (SubCellInst_SboxInst_5_n10), .B0_t (SubCellInst_SboxInst_5_n9), .Z0_t (Feedback[23]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U14 ( .A0_t (Output[45]), .B0_t (SubCellInst_SboxInst_5_n8), .Z0_t (SubCellInst_SboxInst_5_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_U13 ( .A0_t (SubCellInst_SboxInst_5_n8), .B0_t (SubCellInst_SboxInst_5_n7), .Z0_t (Feedback[20]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_U12 ( .A0_t (Output[45]), .B0_t (SubCellInst_SboxInst_5_n6), .Z0_t (SubCellInst_SboxInst_5_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_U11 ( .A0_t (Output[44]), .B0_t (SubCellInst_SboxInst_5_n5), .Z0_t (SubCellInst_SboxInst_5_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_U10 ( .A0_t (Output[47]), .B0_t (Output[46]), .Z0_t (SubCellInst_SboxInst_5_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_U9 ( .A0_t (Output[47]), .B0_t (Output[46]), .Z0_t (SubCellInst_SboxInst_5_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U8 ( .A0_t (SubCellInst_SboxInst_5_n10), .B0_t (SubCellInst_SboxInst_5_n3), .Z0_t (Feedback[22]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U7 ( .A0_t (SubCellInst_SboxInst_5_n2), .B0_t (Output[45]), .Z0_t (SubCellInst_SboxInst_5_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U6 ( .A0_t (SubCellInst_SboxInst_5_n1), .B0_t (Output[46]), .Z0_t (SubCellInst_SboxInst_5_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U4 ( .A0_t (Output[47]), .B0_t (Output[44]), .Z0_t (SubCellInst_SboxInst_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U3 ( .A0_t (Output[44]), .B0_t (Output[47]), .Z0_t (SubCellInst_SboxInst_5_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U19 ( .A0_t (SubCellInst_SboxInst_6_n15), .B0_t (SubCellInst_SboxInst_6_n14), .Z0_t (Feedback[25]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U18 ( .A0_t (Output[42]), .B0_t (SubCellInst_SboxInst_6_n13), .Z0_t (SubCellInst_SboxInst_6_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U17 ( .A0_t (Output[43]), .B0_t (Output[40]), .Z0_t (SubCellInst_SboxInst_6_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U16 ( .A0_t (Output[40]), .B0_t (Output[43]), .Z0_t (SubCellInst_SboxInst_6_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U15 ( .A0_t (SubCellInst_SboxInst_6_n10), .B0_t (SubCellInst_SboxInst_6_n9), .Z0_t (Feedback[27]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U14 ( .A0_t (Output[41]), .B0_t (SubCellInst_SboxInst_6_n8), .Z0_t (SubCellInst_SboxInst_6_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_U13 ( .A0_t (SubCellInst_SboxInst_6_n8), .B0_t (SubCellInst_SboxInst_6_n7), .Z0_t (Feedback[24]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_U12 ( .A0_t (Output[41]), .B0_t (SubCellInst_SboxInst_6_n6), .Z0_t (SubCellInst_SboxInst_6_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_U11 ( .A0_t (Output[40]), .B0_t (SubCellInst_SboxInst_6_n5), .Z0_t (SubCellInst_SboxInst_6_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_U10 ( .A0_t (Output[43]), .B0_t (Output[42]), .Z0_t (SubCellInst_SboxInst_6_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_U9 ( .A0_t (Output[43]), .B0_t (Output[42]), .Z0_t (SubCellInst_SboxInst_6_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U8 ( .A0_t (SubCellInst_SboxInst_6_n10), .B0_t (SubCellInst_SboxInst_6_n3), .Z0_t (Feedback[26]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U7 ( .A0_t (SubCellInst_SboxInst_6_n2), .B0_t (Output[41]), .Z0_t (SubCellInst_SboxInst_6_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U6 ( .A0_t (SubCellInst_SboxInst_6_n1), .B0_t (Output[42]), .Z0_t (SubCellInst_SboxInst_6_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U4 ( .A0_t (Output[43]), .B0_t (Output[40]), .Z0_t (SubCellInst_SboxInst_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U3 ( .A0_t (Output[40]), .B0_t (Output[43]), .Z0_t (SubCellInst_SboxInst_6_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U19 ( .A0_t (SubCellInst_SboxInst_7_n15), .B0_t (SubCellInst_SboxInst_7_n14), .Z0_t (Feedback[29]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U18 ( .A0_t (Output[38]), .B0_t (SubCellInst_SboxInst_7_n13), .Z0_t (SubCellInst_SboxInst_7_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U17 ( .A0_t (Output[39]), .B0_t (Output[36]), .Z0_t (SubCellInst_SboxInst_7_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U16 ( .A0_t (Output[36]), .B0_t (Output[39]), .Z0_t (SubCellInst_SboxInst_7_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U15 ( .A0_t (SubCellInst_SboxInst_7_n10), .B0_t (SubCellInst_SboxInst_7_n9), .Z0_t (Feedback[31]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U14 ( .A0_t (Output[37]), .B0_t (SubCellInst_SboxInst_7_n8), .Z0_t (SubCellInst_SboxInst_7_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_U13 ( .A0_t (SubCellInst_SboxInst_7_n8), .B0_t (SubCellInst_SboxInst_7_n7), .Z0_t (Feedback[28]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_U12 ( .A0_t (Output[37]), .B0_t (SubCellInst_SboxInst_7_n6), .Z0_t (SubCellInst_SboxInst_7_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_U11 ( .A0_t (Output[36]), .B0_t (SubCellInst_SboxInst_7_n5), .Z0_t (SubCellInst_SboxInst_7_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_U10 ( .A0_t (Output[39]), .B0_t (Output[38]), .Z0_t (SubCellInst_SboxInst_7_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_U9 ( .A0_t (Output[39]), .B0_t (Output[38]), .Z0_t (SubCellInst_SboxInst_7_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U8 ( .A0_t (SubCellInst_SboxInst_7_n10), .B0_t (SubCellInst_SboxInst_7_n3), .Z0_t (Feedback[30]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U7 ( .A0_t (SubCellInst_SboxInst_7_n2), .B0_t (Output[37]), .Z0_t (SubCellInst_SboxInst_7_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U6 ( .A0_t (SubCellInst_SboxInst_7_n1), .B0_t (Output[38]), .Z0_t (SubCellInst_SboxInst_7_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U4 ( .A0_t (Output[39]), .B0_t (Output[36]), .Z0_t (SubCellInst_SboxInst_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U3 ( .A0_t (Output[36]), .B0_t (Output[39]), .Z0_t (SubCellInst_SboxInst_7_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U19 ( .A0_t (SubCellInst_SboxInst_8_n15), .B0_t (SubCellInst_SboxInst_8_n14), .Z0_t (Feedback[33]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U18 ( .A0_t (Output[16]), .B0_t (SubCellInst_SboxInst_8_n13), .Z0_t (SubCellInst_SboxInst_8_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U17 ( .A0_t (Output[19]), .B0_t (Output[18]), .Z0_t (SubCellInst_SboxInst_8_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U16 ( .A0_t (Output[18]), .B0_t (Output[19]), .Z0_t (SubCellInst_SboxInst_8_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U15 ( .A0_t (SubCellInst_SboxInst_8_n10), .B0_t (SubCellInst_SboxInst_8_n9), .Z0_t (Feedback[35]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U14 ( .A0_t (SubCellInst_SboxInst_8_n8), .B0_t (Output[17]), .Z0_t (SubCellInst_SboxInst_8_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U13 ( .A0_t (SubCellInst_SboxInst_8_n10), .B0_t (SubCellInst_SboxInst_8_n7), .Z0_t (Feedback[34]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U12 ( .A0_t (SubCellInst_SboxInst_8_n6), .B0_t (Output[17]), .Z0_t (SubCellInst_SboxInst_8_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U11 ( .A0_t (SubCellInst_SboxInst_8_n5), .B0_t (Output[18]), .Z0_t (SubCellInst_SboxInst_8_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U10 ( .A0_t (Output[16]), .B0_t (Output[19]), .Z0_t (SubCellInst_SboxInst_8_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U9 ( .A0_t (Output[19]), .B0_t (Output[16]), .Z0_t (SubCellInst_SboxInst_8_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_U8 ( .A0_t (SubCellInst_SboxInst_8_n8), .B0_t (SubCellInst_SboxInst_8_n3), .Z0_t (Feedback[32]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_U7 ( .A0_t (Output[17]), .B0_t (SubCellInst_SboxInst_8_n2), .Z0_t (SubCellInst_SboxInst_8_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_U6 ( .A0_t (Output[16]), .B0_t (SubCellInst_SboxInst_8_n1), .Z0_t (SubCellInst_SboxInst_8_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_U5 ( .A0_t (Output[18]), .B0_t (Output[19]), .Z0_t (SubCellInst_SboxInst_8_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_U3 ( .A0_t (Output[18]), .B0_t (Output[19]), .Z0_t (SubCellInst_SboxInst_8_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U19 ( .A0_t (SubCellInst_SboxInst_9_n15), .B0_t (SubCellInst_SboxInst_9_n14), .Z0_t (Feedback[37]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U18 ( .A0_t (Output[28]), .B0_t (SubCellInst_SboxInst_9_n13), .Z0_t (SubCellInst_SboxInst_9_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U17 ( .A0_t (Output[31]), .B0_t (Output[30]), .Z0_t (SubCellInst_SboxInst_9_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U16 ( .A0_t (Output[30]), .B0_t (Output[31]), .Z0_t (SubCellInst_SboxInst_9_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U15 ( .A0_t (SubCellInst_SboxInst_9_n10), .B0_t (SubCellInst_SboxInst_9_n9), .Z0_t (Feedback[39]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U14 ( .A0_t (SubCellInst_SboxInst_9_n8), .B0_t (Output[29]), .Z0_t (SubCellInst_SboxInst_9_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U13 ( .A0_t (SubCellInst_SboxInst_9_n10), .B0_t (SubCellInst_SboxInst_9_n7), .Z0_t (Feedback[38]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U12 ( .A0_t (SubCellInst_SboxInst_9_n6), .B0_t (Output[29]), .Z0_t (SubCellInst_SboxInst_9_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U11 ( .A0_t (SubCellInst_SboxInst_9_n5), .B0_t (Output[30]), .Z0_t (SubCellInst_SboxInst_9_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U10 ( .A0_t (Output[28]), .B0_t (Output[31]), .Z0_t (SubCellInst_SboxInst_9_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U9 ( .A0_t (Output[31]), .B0_t (Output[28]), .Z0_t (SubCellInst_SboxInst_9_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_U8 ( .A0_t (SubCellInst_SboxInst_9_n8), .B0_t (SubCellInst_SboxInst_9_n3), .Z0_t (Feedback[36]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_U7 ( .A0_t (Output[29]), .B0_t (SubCellInst_SboxInst_9_n2), .Z0_t (SubCellInst_SboxInst_9_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_U6 ( .A0_t (Output[28]), .B0_t (SubCellInst_SboxInst_9_n1), .Z0_t (SubCellInst_SboxInst_9_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_U5 ( .A0_t (Output[30]), .B0_t (Output[31]), .Z0_t (SubCellInst_SboxInst_9_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_U3 ( .A0_t (Output[30]), .B0_t (Output[31]), .Z0_t (SubCellInst_SboxInst_9_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U19 ( .A0_t (SubCellInst_SboxInst_10_n15), .B0_t (SubCellInst_SboxInst_10_n14), .Z0_t (Feedback[41]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U18 ( .A0_t (Output[24]), .B0_t (SubCellInst_SboxInst_10_n13), .Z0_t (SubCellInst_SboxInst_10_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U17 ( .A0_t (Output[27]), .B0_t (Output[26]), .Z0_t (SubCellInst_SboxInst_10_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U16 ( .A0_t (Output[26]), .B0_t (Output[27]), .Z0_t (SubCellInst_SboxInst_10_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U15 ( .A0_t (SubCellInst_SboxInst_10_n10), .B0_t (SubCellInst_SboxInst_10_n9), .Z0_t (Feedback[43]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U14 ( .A0_t (SubCellInst_SboxInst_10_n8), .B0_t (Output[25]), .Z0_t (SubCellInst_SboxInst_10_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U13 ( .A0_t (SubCellInst_SboxInst_10_n10), .B0_t (SubCellInst_SboxInst_10_n7), .Z0_t (Feedback[42]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U12 ( .A0_t (SubCellInst_SboxInst_10_n6), .B0_t (Output[25]), .Z0_t (SubCellInst_SboxInst_10_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U11 ( .A0_t (SubCellInst_SboxInst_10_n5), .B0_t (Output[26]), .Z0_t (SubCellInst_SboxInst_10_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U10 ( .A0_t (Output[24]), .B0_t (Output[27]), .Z0_t (SubCellInst_SboxInst_10_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U9 ( .A0_t (Output[27]), .B0_t (Output[24]), .Z0_t (SubCellInst_SboxInst_10_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_U8 ( .A0_t (SubCellInst_SboxInst_10_n8), .B0_t (SubCellInst_SboxInst_10_n3), .Z0_t (Feedback[40]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_U7 ( .A0_t (Output[25]), .B0_t (SubCellInst_SboxInst_10_n2), .Z0_t (SubCellInst_SboxInst_10_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_U6 ( .A0_t (Output[24]), .B0_t (SubCellInst_SboxInst_10_n1), .Z0_t (SubCellInst_SboxInst_10_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_U5 ( .A0_t (Output[26]), .B0_t (Output[27]), .Z0_t (SubCellInst_SboxInst_10_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_U3 ( .A0_t (Output[26]), .B0_t (Output[27]), .Z0_t (SubCellInst_SboxInst_10_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U19 ( .A0_t (SubCellInst_SboxInst_11_n15), .B0_t (SubCellInst_SboxInst_11_n14), .Z0_t (Feedback[45]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U18 ( .A0_t (Output[20]), .B0_t (SubCellInst_SboxInst_11_n13), .Z0_t (SubCellInst_SboxInst_11_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U17 ( .A0_t (Output[23]), .B0_t (Output[22]), .Z0_t (SubCellInst_SboxInst_11_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U16 ( .A0_t (Output[22]), .B0_t (Output[23]), .Z0_t (SubCellInst_SboxInst_11_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U15 ( .A0_t (SubCellInst_SboxInst_11_n10), .B0_t (SubCellInst_SboxInst_11_n9), .Z0_t (Feedback[47]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U14 ( .A0_t (SubCellInst_SboxInst_11_n8), .B0_t (Output[21]), .Z0_t (SubCellInst_SboxInst_11_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U13 ( .A0_t (SubCellInst_SboxInst_11_n10), .B0_t (SubCellInst_SboxInst_11_n7), .Z0_t (Feedback[46]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U12 ( .A0_t (SubCellInst_SboxInst_11_n6), .B0_t (Output[21]), .Z0_t (SubCellInst_SboxInst_11_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U11 ( .A0_t (SubCellInst_SboxInst_11_n5), .B0_t (Output[22]), .Z0_t (SubCellInst_SboxInst_11_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U10 ( .A0_t (Output[20]), .B0_t (Output[23]), .Z0_t (SubCellInst_SboxInst_11_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U9 ( .A0_t (Output[23]), .B0_t (Output[20]), .Z0_t (SubCellInst_SboxInst_11_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_U8 ( .A0_t (SubCellInst_SboxInst_11_n8), .B0_t (SubCellInst_SboxInst_11_n3), .Z0_t (Feedback[44]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_U7 ( .A0_t (Output[21]), .B0_t (SubCellInst_SboxInst_11_n2), .Z0_t (SubCellInst_SboxInst_11_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_U6 ( .A0_t (Output[20]), .B0_t (SubCellInst_SboxInst_11_n1), .Z0_t (SubCellInst_SboxInst_11_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_U5 ( .A0_t (Output[22]), .B0_t (Output[23]), .Z0_t (SubCellInst_SboxInst_11_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_U3 ( .A0_t (Output[22]), .B0_t (Output[23]), .Z0_t (SubCellInst_SboxInst_11_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U19 ( .A0_t (SubCellInst_SboxInst_12_n15), .B0_t (SubCellInst_SboxInst_12_n14), .Z0_t (Feedback[49]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U18 ( .A0_t (Output[4]), .B0_t (SubCellInst_SboxInst_12_n13), .Z0_t (SubCellInst_SboxInst_12_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U17 ( .A0_t (Output[7]), .B0_t (Output[6]), .Z0_t (SubCellInst_SboxInst_12_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U16 ( .A0_t (Output[6]), .B0_t (Output[7]), .Z0_t (SubCellInst_SboxInst_12_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U15 ( .A0_t (SubCellInst_SboxInst_12_n10), .B0_t (SubCellInst_SboxInst_12_n9), .Z0_t (Feedback[51]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U14 ( .A0_t (SubCellInst_SboxInst_12_n8), .B0_t (Output[5]), .Z0_t (SubCellInst_SboxInst_12_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U13 ( .A0_t (SubCellInst_SboxInst_12_n10), .B0_t (SubCellInst_SboxInst_12_n7), .Z0_t (Feedback[50]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U12 ( .A0_t (SubCellInst_SboxInst_12_n6), .B0_t (Output[5]), .Z0_t (SubCellInst_SboxInst_12_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U11 ( .A0_t (SubCellInst_SboxInst_12_n5), .B0_t (Output[6]), .Z0_t (SubCellInst_SboxInst_12_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U10 ( .A0_t (Output[4]), .B0_t (Output[7]), .Z0_t (SubCellInst_SboxInst_12_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U9 ( .A0_t (Output[7]), .B0_t (Output[4]), .Z0_t (SubCellInst_SboxInst_12_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_U8 ( .A0_t (SubCellInst_SboxInst_12_n8), .B0_t (SubCellInst_SboxInst_12_n3), .Z0_t (Feedback[48]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_U7 ( .A0_t (Output[5]), .B0_t (SubCellInst_SboxInst_12_n2), .Z0_t (SubCellInst_SboxInst_12_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_U6 ( .A0_t (Output[4]), .B0_t (SubCellInst_SboxInst_12_n1), .Z0_t (SubCellInst_SboxInst_12_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_U5 ( .A0_t (Output[6]), .B0_t (Output[7]), .Z0_t (SubCellInst_SboxInst_12_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_U3 ( .A0_t (Output[6]), .B0_t (Output[7]), .Z0_t (SubCellInst_SboxInst_12_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U19 ( .A0_t (SubCellInst_SboxInst_13_n15), .B0_t (SubCellInst_SboxInst_13_n14), .Z0_t (Feedback[53]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U18 ( .A0_t (Output[8]), .B0_t (SubCellInst_SboxInst_13_n13), .Z0_t (SubCellInst_SboxInst_13_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U17 ( .A0_t (Output[11]), .B0_t (Output[10]), .Z0_t (SubCellInst_SboxInst_13_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U16 ( .A0_t (Output[10]), .B0_t (Output[11]), .Z0_t (SubCellInst_SboxInst_13_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U15 ( .A0_t (SubCellInst_SboxInst_13_n10), .B0_t (SubCellInst_SboxInst_13_n9), .Z0_t (Feedback[55]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U14 ( .A0_t (SubCellInst_SboxInst_13_n8), .B0_t (Output[9]), .Z0_t (SubCellInst_SboxInst_13_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U13 ( .A0_t (SubCellInst_SboxInst_13_n10), .B0_t (SubCellInst_SboxInst_13_n7), .Z0_t (Feedback[54]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U12 ( .A0_t (SubCellInst_SboxInst_13_n6), .B0_t (Output[9]), .Z0_t (SubCellInst_SboxInst_13_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U11 ( .A0_t (SubCellInst_SboxInst_13_n5), .B0_t (Output[10]), .Z0_t (SubCellInst_SboxInst_13_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U10 ( .A0_t (Output[8]), .B0_t (Output[11]), .Z0_t (SubCellInst_SboxInst_13_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U9 ( .A0_t (Output[11]), .B0_t (Output[8]), .Z0_t (SubCellInst_SboxInst_13_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_U8 ( .A0_t (SubCellInst_SboxInst_13_n8), .B0_t (SubCellInst_SboxInst_13_n3), .Z0_t (Feedback[52]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_U7 ( .A0_t (Output[9]), .B0_t (SubCellInst_SboxInst_13_n2), .Z0_t (SubCellInst_SboxInst_13_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_U6 ( .A0_t (Output[8]), .B0_t (SubCellInst_SboxInst_13_n1), .Z0_t (SubCellInst_SboxInst_13_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_U5 ( .A0_t (Output[10]), .B0_t (Output[11]), .Z0_t (SubCellInst_SboxInst_13_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_U3 ( .A0_t (Output[10]), .B0_t (Output[11]), .Z0_t (SubCellInst_SboxInst_13_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U19 ( .A0_t (SubCellInst_SboxInst_14_n15), .B0_t (SubCellInst_SboxInst_14_n14), .Z0_t (Feedback[57]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U18 ( .A0_t (Output[12]), .B0_t (SubCellInst_SboxInst_14_n13), .Z0_t (SubCellInst_SboxInst_14_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U17 ( .A0_t (Output[15]), .B0_t (Output[14]), .Z0_t (SubCellInst_SboxInst_14_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U16 ( .A0_t (Output[14]), .B0_t (Output[15]), .Z0_t (SubCellInst_SboxInst_14_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U15 ( .A0_t (SubCellInst_SboxInst_14_n10), .B0_t (SubCellInst_SboxInst_14_n9), .Z0_t (Feedback[59]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U14 ( .A0_t (SubCellInst_SboxInst_14_n8), .B0_t (Output[13]), .Z0_t (SubCellInst_SboxInst_14_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U13 ( .A0_t (SubCellInst_SboxInst_14_n10), .B0_t (SubCellInst_SboxInst_14_n7), .Z0_t (Feedback[58]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U12 ( .A0_t (SubCellInst_SboxInst_14_n6), .B0_t (Output[13]), .Z0_t (SubCellInst_SboxInst_14_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U11 ( .A0_t (SubCellInst_SboxInst_14_n5), .B0_t (Output[14]), .Z0_t (SubCellInst_SboxInst_14_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U10 ( .A0_t (Output[12]), .B0_t (Output[15]), .Z0_t (SubCellInst_SboxInst_14_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U9 ( .A0_t (Output[15]), .B0_t (Output[12]), .Z0_t (SubCellInst_SboxInst_14_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_U8 ( .A0_t (SubCellInst_SboxInst_14_n8), .B0_t (SubCellInst_SboxInst_14_n3), .Z0_t (Feedback[56]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_U7 ( .A0_t (Output[13]), .B0_t (SubCellInst_SboxInst_14_n2), .Z0_t (SubCellInst_SboxInst_14_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_U6 ( .A0_t (Output[12]), .B0_t (SubCellInst_SboxInst_14_n1), .Z0_t (SubCellInst_SboxInst_14_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_U5 ( .A0_t (Output[14]), .B0_t (Output[15]), .Z0_t (SubCellInst_SboxInst_14_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_U3 ( .A0_t (Output[14]), .B0_t (Output[15]), .Z0_t (SubCellInst_SboxInst_14_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U19 ( .A0_t (SubCellInst_SboxInst_15_n15), .B0_t (SubCellInst_SboxInst_15_n14), .Z0_t (Feedback[61]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U18 ( .A0_t (Output[0]), .B0_t (SubCellInst_SboxInst_15_n13), .Z0_t (SubCellInst_SboxInst_15_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U17 ( .A0_t (Output[3]), .B0_t (Output[2]), .Z0_t (SubCellInst_SboxInst_15_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U16 ( .A0_t (Output[2]), .B0_t (Output[3]), .Z0_t (SubCellInst_SboxInst_15_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U15 ( .A0_t (SubCellInst_SboxInst_15_n10), .B0_t (SubCellInst_SboxInst_15_n9), .Z0_t (Feedback[63]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U14 ( .A0_t (SubCellInst_SboxInst_15_n8), .B0_t (Output[1]), .Z0_t (SubCellInst_SboxInst_15_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U13 ( .A0_t (SubCellInst_SboxInst_15_n10), .B0_t (SubCellInst_SboxInst_15_n7), .Z0_t (Feedback[62]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U12 ( .A0_t (SubCellInst_SboxInst_15_n6), .B0_t (Output[1]), .Z0_t (SubCellInst_SboxInst_15_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U11 ( .A0_t (SubCellInst_SboxInst_15_n5), .B0_t (Output[2]), .Z0_t (SubCellInst_SboxInst_15_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U10 ( .A0_t (Output[0]), .B0_t (Output[3]), .Z0_t (SubCellInst_SboxInst_15_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U9 ( .A0_t (Output[3]), .B0_t (Output[0]), .Z0_t (SubCellInst_SboxInst_15_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_U8 ( .A0_t (SubCellInst_SboxInst_15_n8), .B0_t (SubCellInst_SboxInst_15_n3), .Z0_t (Feedback[60]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_U7 ( .A0_t (Output[1]), .B0_t (SubCellInst_SboxInst_15_n2), .Z0_t (SubCellInst_SboxInst_15_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_U6 ( .A0_t (Output[0]), .B0_t (SubCellInst_SboxInst_15_n1), .Z0_t (SubCellInst_SboxInst_15_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_U5 ( .A0_t (Output[2]), .B0_t (Output[3]), .Z0_t (SubCellInst_SboxInst_15_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_U3 ( .A0_t (Output[2]), .B0_t (Output[3]), .Z0_t (SubCellInst_SboxInst_15_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_0_U1_XOR1_U1 ( .A0_t (Key[64]), .B0_t (Key[0]), .Z0_t (KeyMUX_MUXInst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_0_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_0_U1_X), .Z0_t (KeyMUX_MUXInst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_0_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_0_U1_Y), .B0_t (Key[64]), .Z0_t (SelectedKey[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_1_U1_XOR1_U1 ( .A0_t (Key[65]), .B0_t (Key[1]), .Z0_t (KeyMUX_MUXInst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_1_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_1_U1_X), .Z0_t (KeyMUX_MUXInst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_1_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_1_U1_Y), .B0_t (Key[65]), .Z0_t (SelectedKey[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_2_U1_XOR1_U1 ( .A0_t (Key[66]), .B0_t (Key[2]), .Z0_t (KeyMUX_MUXInst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_2_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_2_U1_X), .Z0_t (KeyMUX_MUXInst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_2_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_2_U1_Y), .B0_t (Key[66]), .Z0_t (SelectedKey[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_3_U1_XOR1_U1 ( .A0_t (Key[67]), .B0_t (Key[3]), .Z0_t (KeyMUX_MUXInst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_3_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_3_U1_X), .Z0_t (KeyMUX_MUXInst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_3_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_3_U1_Y), .B0_t (Key[67]), .Z0_t (SelectedKey[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_4_U1_XOR1_U1 ( .A0_t (Key[68]), .B0_t (Key[4]), .Z0_t (KeyMUX_MUXInst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_4_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_4_U1_X), .Z0_t (KeyMUX_MUXInst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_4_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_4_U1_Y), .B0_t (Key[68]), .Z0_t (SelectedKey[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_5_U1_XOR1_U1 ( .A0_t (Key[69]), .B0_t (Key[5]), .Z0_t (KeyMUX_MUXInst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_5_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_5_U1_X), .Z0_t (KeyMUX_MUXInst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_5_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_5_U1_Y), .B0_t (Key[69]), .Z0_t (SelectedKey[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_6_U1_XOR1_U1 ( .A0_t (Key[70]), .B0_t (Key[6]), .Z0_t (KeyMUX_MUXInst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_6_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_6_U1_X), .Z0_t (KeyMUX_MUXInst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_6_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_6_U1_Y), .B0_t (Key[70]), .Z0_t (SelectedKey[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_7_U1_XOR1_U1 ( .A0_t (Key[71]), .B0_t (Key[7]), .Z0_t (KeyMUX_MUXInst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_7_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_7_U1_X), .Z0_t (KeyMUX_MUXInst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_7_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_7_U1_Y), .B0_t (Key[71]), .Z0_t (SelectedKey[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_8_U1_XOR1_U1 ( .A0_t (Key[72]), .B0_t (Key[8]), .Z0_t (KeyMUX_MUXInst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_8_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_8_U1_X), .Z0_t (KeyMUX_MUXInst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_8_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_8_U1_Y), .B0_t (Key[72]), .Z0_t (SelectedKey[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_9_U1_XOR1_U1 ( .A0_t (Key[73]), .B0_t (Key[9]), .Z0_t (KeyMUX_MUXInst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_9_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_9_U1_X), .Z0_t (KeyMUX_MUXInst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_9_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_9_U1_Y), .B0_t (Key[73]), .Z0_t (SelectedKey[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_10_U1_XOR1_U1 ( .A0_t (Key[74]), .B0_t (Key[10]), .Z0_t (KeyMUX_MUXInst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_10_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_10_U1_X), .Z0_t (KeyMUX_MUXInst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_10_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_10_U1_Y), .B0_t (Key[74]), .Z0_t (SelectedKey[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_11_U1_XOR1_U1 ( .A0_t (Key[75]), .B0_t (Key[11]), .Z0_t (KeyMUX_MUXInst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_11_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_11_U1_X), .Z0_t (KeyMUX_MUXInst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_11_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_11_U1_Y), .B0_t (Key[75]), .Z0_t (SelectedKey[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_12_U1_XOR1_U1 ( .A0_t (Key[76]), .B0_t (Key[12]), .Z0_t (KeyMUX_MUXInst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_12_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_12_U1_X), .Z0_t (KeyMUX_MUXInst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_12_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_12_U1_Y), .B0_t (Key[76]), .Z0_t (SelectedKey[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_13_U1_XOR1_U1 ( .A0_t (Key[77]), .B0_t (Key[13]), .Z0_t (KeyMUX_MUXInst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_13_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_13_U1_X), .Z0_t (KeyMUX_MUXInst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_13_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_13_U1_Y), .B0_t (Key[77]), .Z0_t (SelectedKey[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_14_U1_XOR1_U1 ( .A0_t (Key[78]), .B0_t (Key[14]), .Z0_t (KeyMUX_MUXInst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_14_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_14_U1_X), .Z0_t (KeyMUX_MUXInst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_14_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_14_U1_Y), .B0_t (Key[78]), .Z0_t (SelectedKey[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_15_U1_XOR1_U1 ( .A0_t (Key[79]), .B0_t (Key[15]), .Z0_t (KeyMUX_MUXInst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_15_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_15_U1_X), .Z0_t (KeyMUX_MUXInst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_15_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_15_U1_Y), .B0_t (Key[79]), .Z0_t (SelectedKey[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_16_U1_XOR1_U1 ( .A0_t (Key[80]), .B0_t (Key[16]), .Z0_t (KeyMUX_MUXInst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_16_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_16_U1_X), .Z0_t (KeyMUX_MUXInst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_16_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_16_U1_Y), .B0_t (Key[80]), .Z0_t (SelectedKey[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_17_U1_XOR1_U1 ( .A0_t (Key[81]), .B0_t (Key[17]), .Z0_t (KeyMUX_MUXInst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_17_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_17_U1_X), .Z0_t (KeyMUX_MUXInst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_17_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_17_U1_Y), .B0_t (Key[81]), .Z0_t (SelectedKey[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_18_U1_XOR1_U1 ( .A0_t (Key[82]), .B0_t (Key[18]), .Z0_t (KeyMUX_MUXInst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_18_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_18_U1_X), .Z0_t (KeyMUX_MUXInst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_18_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_18_U1_Y), .B0_t (Key[82]), .Z0_t (SelectedKey[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_19_U1_XOR1_U1 ( .A0_t (Key[83]), .B0_t (Key[19]), .Z0_t (KeyMUX_MUXInst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_19_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_19_U1_X), .Z0_t (KeyMUX_MUXInst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_19_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_19_U1_Y), .B0_t (Key[83]), .Z0_t (SelectedKey[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_20_U1_XOR1_U1 ( .A0_t (Key[84]), .B0_t (Key[20]), .Z0_t (KeyMUX_MUXInst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_20_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_20_U1_X), .Z0_t (KeyMUX_MUXInst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_20_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_20_U1_Y), .B0_t (Key[84]), .Z0_t (SelectedKey[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_21_U1_XOR1_U1 ( .A0_t (Key[85]), .B0_t (Key[21]), .Z0_t (KeyMUX_MUXInst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_21_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_21_U1_X), .Z0_t (KeyMUX_MUXInst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_21_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_21_U1_Y), .B0_t (Key[85]), .Z0_t (SelectedKey[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_22_U1_XOR1_U1 ( .A0_t (Key[86]), .B0_t (Key[22]), .Z0_t (KeyMUX_MUXInst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_22_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_22_U1_X), .Z0_t (KeyMUX_MUXInst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_22_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_22_U1_Y), .B0_t (Key[86]), .Z0_t (SelectedKey[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_23_U1_XOR1_U1 ( .A0_t (Key[87]), .B0_t (Key[23]), .Z0_t (KeyMUX_MUXInst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_23_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_23_U1_X), .Z0_t (KeyMUX_MUXInst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_23_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_23_U1_Y), .B0_t (Key[87]), .Z0_t (SelectedKey[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_24_U1_XOR1_U1 ( .A0_t (Key[88]), .B0_t (Key[24]), .Z0_t (KeyMUX_MUXInst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_24_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_24_U1_X), .Z0_t (KeyMUX_MUXInst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_24_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_24_U1_Y), .B0_t (Key[88]), .Z0_t (SelectedKey[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_25_U1_XOR1_U1 ( .A0_t (Key[89]), .B0_t (Key[25]), .Z0_t (KeyMUX_MUXInst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_25_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_25_U1_X), .Z0_t (KeyMUX_MUXInst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_25_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_25_U1_Y), .B0_t (Key[89]), .Z0_t (SelectedKey[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_26_U1_XOR1_U1 ( .A0_t (Key[90]), .B0_t (Key[26]), .Z0_t (KeyMUX_MUXInst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_26_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_26_U1_X), .Z0_t (KeyMUX_MUXInst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_26_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_26_U1_Y), .B0_t (Key[90]), .Z0_t (SelectedKey[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_27_U1_XOR1_U1 ( .A0_t (Key[91]), .B0_t (Key[27]), .Z0_t (KeyMUX_MUXInst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_27_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_27_U1_X), .Z0_t (KeyMUX_MUXInst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_27_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_27_U1_Y), .B0_t (Key[91]), .Z0_t (SelectedKey[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_28_U1_XOR1_U1 ( .A0_t (Key[92]), .B0_t (Key[28]), .Z0_t (KeyMUX_MUXInst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_28_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_28_U1_X), .Z0_t (KeyMUX_MUXInst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_28_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_28_U1_Y), .B0_t (Key[92]), .Z0_t (SelectedKey[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_29_U1_XOR1_U1 ( .A0_t (Key[93]), .B0_t (Key[29]), .Z0_t (KeyMUX_MUXInst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_29_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_29_U1_X), .Z0_t (KeyMUX_MUXInst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_29_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_29_U1_Y), .B0_t (Key[93]), .Z0_t (SelectedKey[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_30_U1_XOR1_U1 ( .A0_t (Key[94]), .B0_t (Key[30]), .Z0_t (KeyMUX_MUXInst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_30_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_30_U1_X), .Z0_t (KeyMUX_MUXInst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_30_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_30_U1_Y), .B0_t (Key[94]), .Z0_t (SelectedKey[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_31_U1_XOR1_U1 ( .A0_t (Key[95]), .B0_t (Key[31]), .Z0_t (KeyMUX_MUXInst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_31_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_31_U1_X), .Z0_t (KeyMUX_MUXInst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_31_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_31_U1_Y), .B0_t (Key[95]), .Z0_t (SelectedKey[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_32_U1_XOR1_U1 ( .A0_t (Key[96]), .B0_t (Key[32]), .Z0_t (KeyMUX_MUXInst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_32_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_32_U1_X), .Z0_t (KeyMUX_MUXInst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_32_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_32_U1_Y), .B0_t (Key[96]), .Z0_t (SelectedKey[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_33_U1_XOR1_U1 ( .A0_t (Key[97]), .B0_t (Key[33]), .Z0_t (KeyMUX_MUXInst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_33_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_33_U1_X), .Z0_t (KeyMUX_MUXInst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_33_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_33_U1_Y), .B0_t (Key[97]), .Z0_t (SelectedKey[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_34_U1_XOR1_U1 ( .A0_t (Key[98]), .B0_t (Key[34]), .Z0_t (KeyMUX_MUXInst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_34_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_34_U1_X), .Z0_t (KeyMUX_MUXInst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_34_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_34_U1_Y), .B0_t (Key[98]), .Z0_t (SelectedKey[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_35_U1_XOR1_U1 ( .A0_t (Key[99]), .B0_t (Key[35]), .Z0_t (KeyMUX_MUXInst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_35_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_35_U1_X), .Z0_t (KeyMUX_MUXInst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_35_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_35_U1_Y), .B0_t (Key[99]), .Z0_t (SelectedKey[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_36_U1_XOR1_U1 ( .A0_t (Key[100]), .B0_t (Key[36]), .Z0_t (KeyMUX_MUXInst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_36_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_36_U1_X), .Z0_t (KeyMUX_MUXInst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_36_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_36_U1_Y), .B0_t (Key[100]), .Z0_t (SelectedKey[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_37_U1_XOR1_U1 ( .A0_t (Key[101]), .B0_t (Key[37]), .Z0_t (KeyMUX_MUXInst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_37_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_37_U1_X), .Z0_t (KeyMUX_MUXInst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_37_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_37_U1_Y), .B0_t (Key[101]), .Z0_t (SelectedKey[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_38_U1_XOR1_U1 ( .A0_t (Key[102]), .B0_t (Key[38]), .Z0_t (KeyMUX_MUXInst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_38_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_38_U1_X), .Z0_t (KeyMUX_MUXInst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_38_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_38_U1_Y), .B0_t (Key[102]), .Z0_t (SelectedKey[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_39_U1_XOR1_U1 ( .A0_t (Key[103]), .B0_t (Key[39]), .Z0_t (KeyMUX_MUXInst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_39_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_39_U1_X), .Z0_t (KeyMUX_MUXInst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_39_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_39_U1_Y), .B0_t (Key[103]), .Z0_t (SelectedKey[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_40_U1_XOR1_U1 ( .A0_t (Key[104]), .B0_t (Key[40]), .Z0_t (KeyMUX_MUXInst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_40_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_40_U1_X), .Z0_t (KeyMUX_MUXInst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_40_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_40_U1_Y), .B0_t (Key[104]), .Z0_t (SelectedKey[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_41_U1_XOR1_U1 ( .A0_t (Key[105]), .B0_t (Key[41]), .Z0_t (KeyMUX_MUXInst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_41_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_41_U1_X), .Z0_t (KeyMUX_MUXInst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_41_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_41_U1_Y), .B0_t (Key[105]), .Z0_t (SelectedKey[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_42_U1_XOR1_U1 ( .A0_t (Key[106]), .B0_t (Key[42]), .Z0_t (KeyMUX_MUXInst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_42_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_42_U1_X), .Z0_t (KeyMUX_MUXInst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_42_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_42_U1_Y), .B0_t (Key[106]), .Z0_t (SelectedKey[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_43_U1_XOR1_U1 ( .A0_t (Key[107]), .B0_t (Key[43]), .Z0_t (KeyMUX_MUXInst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_43_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_43_U1_X), .Z0_t (KeyMUX_MUXInst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_43_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_43_U1_Y), .B0_t (Key[107]), .Z0_t (SelectedKey[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_44_U1_XOR1_U1 ( .A0_t (Key[108]), .B0_t (Key[44]), .Z0_t (KeyMUX_MUXInst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_44_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_44_U1_X), .Z0_t (KeyMUX_MUXInst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_44_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_44_U1_Y), .B0_t (Key[108]), .Z0_t (SelectedKey[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_45_U1_XOR1_U1 ( .A0_t (Key[109]), .B0_t (Key[45]), .Z0_t (KeyMUX_MUXInst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_45_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_45_U1_X), .Z0_t (KeyMUX_MUXInst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_45_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_45_U1_Y), .B0_t (Key[109]), .Z0_t (SelectedKey[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_46_U1_XOR1_U1 ( .A0_t (Key[110]), .B0_t (Key[46]), .Z0_t (KeyMUX_MUXInst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_46_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_46_U1_X), .Z0_t (KeyMUX_MUXInst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_46_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_46_U1_Y), .B0_t (Key[110]), .Z0_t (SelectedKey[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_47_U1_XOR1_U1 ( .A0_t (Key[111]), .B0_t (Key[47]), .Z0_t (KeyMUX_MUXInst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_47_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_47_U1_X), .Z0_t (KeyMUX_MUXInst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_47_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_47_U1_Y), .B0_t (Key[111]), .Z0_t (SelectedKey[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_48_U1_XOR1_U1 ( .A0_t (Key[112]), .B0_t (Key[48]), .Z0_t (KeyMUX_MUXInst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_48_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_48_U1_X), .Z0_t (KeyMUX_MUXInst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_48_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_48_U1_Y), .B0_t (Key[112]), .Z0_t (SelectedKey[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_49_U1_XOR1_U1 ( .A0_t (Key[113]), .B0_t (Key[49]), .Z0_t (KeyMUX_MUXInst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_49_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_49_U1_X), .Z0_t (KeyMUX_MUXInst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_49_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_49_U1_Y), .B0_t (Key[113]), .Z0_t (SelectedKey[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_50_U1_XOR1_U1 ( .A0_t (Key[114]), .B0_t (Key[50]), .Z0_t (KeyMUX_MUXInst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_50_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_50_U1_X), .Z0_t (KeyMUX_MUXInst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_50_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_50_U1_Y), .B0_t (Key[114]), .Z0_t (SelectedKey[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_51_U1_XOR1_U1 ( .A0_t (Key[115]), .B0_t (Key[51]), .Z0_t (KeyMUX_MUXInst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_51_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_51_U1_X), .Z0_t (KeyMUX_MUXInst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_51_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_51_U1_Y), .B0_t (Key[115]), .Z0_t (SelectedKey[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_52_U1_XOR1_U1 ( .A0_t (Key[116]), .B0_t (Key[52]), .Z0_t (KeyMUX_MUXInst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_52_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_52_U1_X), .Z0_t (KeyMUX_MUXInst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_52_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_52_U1_Y), .B0_t (Key[116]), .Z0_t (SelectedKey[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_53_U1_XOR1_U1 ( .A0_t (Key[117]), .B0_t (Key[53]), .Z0_t (KeyMUX_MUXInst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_53_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_53_U1_X), .Z0_t (KeyMUX_MUXInst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_53_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_53_U1_Y), .B0_t (Key[117]), .Z0_t (SelectedKey[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_54_U1_XOR1_U1 ( .A0_t (Key[118]), .B0_t (Key[54]), .Z0_t (KeyMUX_MUXInst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_54_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_54_U1_X), .Z0_t (KeyMUX_MUXInst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_54_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_54_U1_Y), .B0_t (Key[118]), .Z0_t (SelectedKey[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_55_U1_XOR1_U1 ( .A0_t (Key[119]), .B0_t (Key[55]), .Z0_t (KeyMUX_MUXInst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_55_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_55_U1_X), .Z0_t (KeyMUX_MUXInst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_55_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_55_U1_Y), .B0_t (Key[119]), .Z0_t (SelectedKey[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_56_U1_XOR1_U1 ( .A0_t (Key[120]), .B0_t (Key[56]), .Z0_t (KeyMUX_MUXInst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_56_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_56_U1_X), .Z0_t (KeyMUX_MUXInst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_56_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_56_U1_Y), .B0_t (Key[120]), .Z0_t (SelectedKey[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_57_U1_XOR1_U1 ( .A0_t (Key[121]), .B0_t (Key[57]), .Z0_t (KeyMUX_MUXInst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_57_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_57_U1_X), .Z0_t (KeyMUX_MUXInst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_57_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_57_U1_Y), .B0_t (Key[121]), .Z0_t (SelectedKey[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_58_U1_XOR1_U1 ( .A0_t (Key[122]), .B0_t (Key[58]), .Z0_t (KeyMUX_MUXInst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_58_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_58_U1_X), .Z0_t (KeyMUX_MUXInst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_58_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_58_U1_Y), .B0_t (Key[122]), .Z0_t (SelectedKey[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_59_U1_XOR1_U1 ( .A0_t (Key[123]), .B0_t (Key[59]), .Z0_t (KeyMUX_MUXInst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_59_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_59_U1_X), .Z0_t (KeyMUX_MUXInst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_59_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_59_U1_Y), .B0_t (Key[123]), .Z0_t (SelectedKey[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_60_U1_XOR1_U1 ( .A0_t (Key[124]), .B0_t (Key[60]), .Z0_t (KeyMUX_MUXInst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_60_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_60_U1_X), .Z0_t (KeyMUX_MUXInst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_60_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_60_U1_Y), .B0_t (Key[124]), .Z0_t (SelectedKey[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_61_U1_XOR1_U1 ( .A0_t (Key[125]), .B0_t (Key[61]), .Z0_t (KeyMUX_MUXInst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_61_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_61_U1_X), .Z0_t (KeyMUX_MUXInst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_61_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_61_U1_Y), .B0_t (Key[125]), .Z0_t (SelectedKey[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_62_U1_XOR1_U1 ( .A0_t (Key[126]), .B0_t (Key[62]), .Z0_t (KeyMUX_MUXInst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_62_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_62_U1_X), .Z0_t (KeyMUX_MUXInst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_62_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_62_U1_Y), .B0_t (Key[126]), .Z0_t (SelectedKey[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_63_U1_XOR1_U1 ( .A0_t (Key[127]), .B0_t (Key[63]), .Z0_t (KeyMUX_MUXInst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_63_U1_AND1_U1 ( .A0_t (selects[0]), .B0_t (KeyMUX_MUXInst_63_U1_X), .Z0_t (KeyMUX_MUXInst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_63_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_63_U1_Y), .B0_t (Key[127]), .Z0_t (SelectedKey[63]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_0_U1 ( .A0_t (FSMReg[0]), .B0_t (rst), .Z0_t (RoundConstant_0) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_1_U2 ( .A0_t (rst), .B0_t (FSMReg[1]), .Z0_t (FSMUpdate[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_2_U2 ( .A0_t (rst), .B0_t (FSMReg[2]), .Z0_t (FSMUpdate[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_3_U1 ( .A0_t (FSMReg[3]), .B0_t (rst), .Z0_t (RoundConstant_4_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_4_U2 ( .A0_t (rst), .B0_t (FSMReg[4]), .Z0_t (FSMUpdate[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_5_U2 ( .A0_t (rst), .B0_t (FSMReg[5]), .Z0_t (FSMUpdate[4]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_6_U2 ( .A0_t (rst), .B0_t (FSMReg[6]), .Z0_t (FSMUpdate[5]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) FSMUpdateInst_U2 ( .A0_t (FSMUpdate[0]), .B0_t (RoundConstant_0), .Z0_t (FSMReg[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) FSMUpdateInst_U1 ( .A0_t (FSMUpdate[3]), .B0_t (RoundConstant_4_), .Z0_t (FSMReg[6]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMSignalsInst_U6 ( .A0_t (RoundConstant_0), .B0_t (FSMSignalsInst_n5), .Z0_t (done) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_U5 ( .A0_t (FSMSignalsInst_n4), .B0_t (FSMSignalsInst_n3), .Z0_t (FSMSignalsInst_n5) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_U4 ( .A0_t (FSMSignalsInst_n2), .B0_t (FSMSignalsInst_n1), .Z0_t (FSMSignalsInst_n3) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_U3 ( .A0_t (RoundConstant_4_), .B0_t (FSMUpdate[0]), .Z0_t (FSMSignalsInst_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_U2 ( .A0_t (FSMUpdate[4]), .B0_t (FSMUpdate[3]), .Z0_t (FSMSignalsInst_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_U1 ( .A0_t (FSMUpdate[1]), .B0_t (FSMUpdate[5]), .Z0_t (FSMSignalsInst_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) selectsMUX_MUXInst_0_U2 ( .A0_t (rst), .B0_t (selectsReg[0]), .Z0_t (selects[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) selectsMUX_MUXInst_1_U2 ( .A0_t (rst), .B0_t (selectsReg[1]), .Z0_t (selects[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b0)) selectsUpdateInst_U2 ( .A0_t (selects[1]), .B0_t (selects[0]), .Z0_t (selectsReg[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_984 ( .A0_t (FSMUpdate[5]), .B0_t (1'b0), .Z0_t (FSMReg[5]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_985 ( .A0_t (FSMUpdate[4]), .B0_t (1'b0), .Z0_t (FSMReg[4]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_986 ( .A0_t (FSMUpdate[3]), .B0_t (1'b0), .Z0_t (FSMReg[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_987 ( .A0_t (FSMUpdate[1]), .B0_t (1'b0), .Z0_t (FSMReg[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_988 ( .A0_t (FSMUpdate[0]), .B0_t (1'b0), .Z0_t (FSMReg[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_989 ( .A0_t (selects[0]), .B0_t (1'b0), .Z0_t (selectsReg[0]) ) ;

    /* register cells */
endmodule
