
module XOR_forMUX_0 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_0 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_511 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_0 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_0 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_0 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_511 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_256 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_256 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_256 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_0 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_0 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_256 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_510 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_255 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_509 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_255 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_510 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_255 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_509 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_255 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_255 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_255 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_255 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_255 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_255 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_508 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_254 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_507 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_254 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_508 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_254 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_507 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_254 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_254 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_254 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_254 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_254 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_254 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_506 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_253 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_505 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_253 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_506 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_253 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_505 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_253 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_253 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_253 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_253 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_253 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_253 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_504 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_252 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_503 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_252 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_504 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_252 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_503 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_252 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_252 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_252 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_252 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_252 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_252 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_502 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_251 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_501 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_251 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_502 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_251 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_501 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_251 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_251 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_251 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_251 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_251 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_251 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_500 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_250 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_499 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_250 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_500 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_250 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_499 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_250 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_250 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_250 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_250 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_250 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_250 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_498 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_249 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_497 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_249 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_498 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_249 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_497 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_249 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_249 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_249 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_249 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_249 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_249 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_496 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_248 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_495 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_248 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_496 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_248 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_495 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_248 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_248 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_248 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_248 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_248 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_248 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_494 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_247 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_493 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_247 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_494 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_247 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_493 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_247 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_247 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_247 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_247 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_247 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_247 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_492 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_246 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_491 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_246 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_492 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_246 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_491 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_246 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_246 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_246 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_246 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_246 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_246 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_490 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_245 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_489 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_245 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_490 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_245 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_489 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_245 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_245 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_245 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_245 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_245 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_245 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_488 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_244 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_487 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_244 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_488 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_244 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_487 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_244 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_244 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_244 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_244 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_244 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_244 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_486 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_243 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_485 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_243 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_486 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_243 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_485 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_243 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_243 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_243 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_243 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_243 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_243 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_484 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_242 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_483 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_242 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_484 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_242 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_483 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_242 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_242 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_242 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_242 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_242 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_242 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_482 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_241 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_481 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_241 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_482 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_241 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_481 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_241 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_241 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_241 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_241 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_241 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_241 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_480 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_240 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_479 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_240 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_480 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_240 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_479 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_240 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_240 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_240 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_240 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_240 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_240 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_478 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_239 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_477 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_239 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_478 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_239 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_477 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_239 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_239 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_239 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_239 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_239 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_239 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_476 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_238 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_475 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_238 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_476 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_238 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_475 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_238 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_238 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_238 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_238 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_238 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_238 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_474 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_237 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_473 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_237 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_474 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_237 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_473 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_237 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_237 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_237 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_237 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_237 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_237 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_472 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_236 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_471 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_236 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_472 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_236 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_471 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_236 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_236 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_236 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_236 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_236 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_236 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_470 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_235 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_469 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_235 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_470 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_235 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_469 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_235 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_235 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_235 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_235 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_235 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_235 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_468 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_234 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_467 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_234 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_468 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_234 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_467 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_234 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_234 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_234 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_234 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_234 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_234 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_466 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_233 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_465 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_233 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_466 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_233 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_465 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_233 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_233 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_233 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_233 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_233 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_233 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_464 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_232 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_463 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_232 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_464 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_232 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_463 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_232 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_232 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_232 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_232 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_232 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_232 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_462 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_231 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_461 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_231 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_462 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_231 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_461 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_231 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_231 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_231 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_231 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_231 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_231 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_460 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_230 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_459 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_230 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_460 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_230 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_459 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_230 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_230 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_230 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_230 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_230 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_230 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_458 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_229 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_457 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_229 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_458 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_229 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_457 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_229 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_229 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_229 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_229 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_229 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_229 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_456 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_228 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_455 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_228 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_456 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_228 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_455 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_228 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_228 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_228 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_228 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_228 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_228 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_454 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_227 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_453 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_227 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_454 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_227 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_453 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_227 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_227 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_227 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_227 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_227 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_227 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_452 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_226 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_451 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_226 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_452 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_226 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_451 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_226 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_226 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_226 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_226 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_226 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_226 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_450 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_225 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_449 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_225 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_450 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_225 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_449 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_225 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_225 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_225 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_225 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_225 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_225 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_448 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_224 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_447 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_224 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_448 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_224 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_447 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_224 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_224 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_224 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_224 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_224 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_224 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_446 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_223 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_445 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_223 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_446 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_223 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_445 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_223 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_223 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_223 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_223 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_223 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_223 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_444 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_222 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_443 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_222 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_444 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_222 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_443 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_222 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_222 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_222 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_222 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_222 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_222 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_442 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_221 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_441 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_221 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_442 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_221 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_441 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_221 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_221 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_221 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_221 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_221 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_221 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_440 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_220 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_439 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_220 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_440 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_220 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_439 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_220 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_220 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_220 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_220 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_220 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_220 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_438 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_219 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_437 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_219 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_438 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_219 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_437 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_219 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_219 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_219 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_219 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_219 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_219 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_436 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_218 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_435 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_218 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_436 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_218 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_435 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_218 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_218 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_218 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_218 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_218 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_218 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_434 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_217 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_433 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_217 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_434 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_217 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_433 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_217 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_217 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_217 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_217 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_217 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_217 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_432 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_216 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_431 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_216 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_432 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_216 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_431 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_216 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_216 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_216 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_216 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_216 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_216 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_430 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_215 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_429 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_215 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_430 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_215 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_429 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_215 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_215 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_215 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_215 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_215 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_215 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_428 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_214 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_427 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_214 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_428 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_214 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_427 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_214 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_214 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_214 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_214 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_214 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_214 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_426 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_213 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_425 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_213 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_426 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_213 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_425 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_213 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_213 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_213 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_213 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_213 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_213 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_424 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_212 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_423 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_212 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_424 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_212 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_423 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_212 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_212 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_212 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_212 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_212 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_212 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_422 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_211 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_421 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_211 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_422 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_211 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_421 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_211 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_211 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_211 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_211 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_211 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_211 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_420 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_210 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_419 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_210 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_420 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_210 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_419 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_210 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_210 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_210 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_210 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_210 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_210 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_418 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_209 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_417 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_209 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_418 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_209 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_417 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_209 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_209 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_209 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_209 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_209 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_209 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_416 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_208 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_415 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_208 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_416 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_208 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_415 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_208 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_208 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_208 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_208 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_208 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_208 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_414 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_207 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_413 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_207 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_414 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_207 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_413 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_207 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_207 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_207 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_207 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_207 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_207 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_412 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_206 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_411 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_206 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_412 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_206 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_411 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_206 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_206 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_206 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_206 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_206 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_206 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_410 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_205 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_409 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_205 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_410 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_205 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_409 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_205 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_205 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_205 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_205 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_205 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_205 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_408 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_204 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_407 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_204 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_408 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_204 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_407 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_204 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_204 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_204 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_204 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_204 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_204 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_406 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_203 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_405 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_203 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_406 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_203 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_405 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_203 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_203 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_203 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_203 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_203 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_203 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_404 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_202 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_403 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_202 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_404 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_202 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_403 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_202 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_202 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_202 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_202 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_202 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_202 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_402 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_201 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_401 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_201 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_402 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_201 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_401 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_201 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_201 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_201 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_201 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_201 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_201 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_400 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_200 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_399 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_200 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_400 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_200 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_399 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_200 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_200 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_200 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_200 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_200 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_200 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_398 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_199 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_397 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_199 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_398 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_199 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_397 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_199 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_199 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_199 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_199 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_199 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_199 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_396 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_198 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_395 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_198 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_396 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_198 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_395 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_198 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_198 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_198 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_198 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_198 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_198 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_394 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_197 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_393 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_197 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_394 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_197 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_393 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_197 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_197 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_197 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_197 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_197 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_197 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_392 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_196 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_391 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_196 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_392 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_196 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_391 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_196 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_196 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_196 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_196 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_196 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_196 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_390 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_195 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_389 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_195 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_390 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_195 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_389 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_195 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_195 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_195 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_195 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_195 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_195 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_388 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_194 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_387 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_194 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_388 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_194 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_387 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_194 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_194 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_194 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_194 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_194 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_194 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_386 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_193 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_385 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_193 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_386 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_193 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_385 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_193 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_193 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_193 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_193 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_193 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_193 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_384 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_192 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_383 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_192 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_384 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_192 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_383 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_192 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_192 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_192 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_192 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_192 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_192 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_382 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_191 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_381 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_191 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_382 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_191 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_381 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_191 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_191 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_191 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_191 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_191 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_191 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_380 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_190 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_379 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_190 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_380 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_190 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_379 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_190 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_190 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_190 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_190 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_190 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_190 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_378 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_189 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_377 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_189 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_378 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_189 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_377 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_189 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_189 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_189 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_189 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_189 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_189 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_376 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_188 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_375 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_188 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_376 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_188 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_375 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_188 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_188 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_188 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_188 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_188 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_188 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_374 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_187 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_373 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_187 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_374 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_187 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_373 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_187 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_187 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_187 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_187 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_187 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_187 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_372 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_186 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_371 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_186 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_372 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_186 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_371 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_186 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_186 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_186 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_186 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_186 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_186 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_370 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_185 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_369 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_185 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_370 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_185 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_369 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_185 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_185 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_185 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_185 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_185 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_185 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_368 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_184 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_367 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_184 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_368 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_184 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_367 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_184 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_184 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_184 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_184 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_184 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_184 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_366 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_183 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_365 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_183 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_366 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_183 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_365 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_183 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_183 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_183 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_183 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_183 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_183 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_364 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_182 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_363 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_182 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_364 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_182 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_363 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_182 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_182 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_182 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_182 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_182 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_182 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_362 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_181 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_361 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_181 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_362 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_181 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_361 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_181 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_181 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_181 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_181 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_181 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_181 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_360 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_180 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_359 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_180 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_360 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_180 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_359 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_180 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_180 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_180 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_180 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_180 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_180 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_358 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_179 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_357 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_179 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_358 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_179 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_357 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_179 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_179 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_179 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_179 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_179 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_179 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_356 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_178 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_355 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_178 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_356 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_178 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_355 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_178 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_178 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_178 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_178 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_178 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_178 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_354 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_177 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_353 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_177 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_354 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_177 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_353 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_177 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_177 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_177 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_177 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_177 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_177 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_352 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_176 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_351 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_176 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_352 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_176 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_351 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_176 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_176 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_176 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_176 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_176 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_176 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_350 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_175 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_349 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_175 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_350 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_175 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_349 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_175 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_175 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_175 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_175 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_175 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_175 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_348 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_174 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_347 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_174 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_348 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_174 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_347 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_174 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_174 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_174 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_174 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_174 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_174 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_346 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_173 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_345 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_173 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_346 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_173 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_345 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_173 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_173 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_173 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_173 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_173 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_173 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_344 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_172 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_343 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_172 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_344 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_172 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_343 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_172 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_172 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_172 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_172 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_172 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_172 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_342 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_171 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_341 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_171 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_342 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_171 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_341 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_171 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_171 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_171 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_171 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_171 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_171 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_340 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_170 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_339 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_170 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_340 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_170 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_339 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_170 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_170 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_170 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_170 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_170 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_170 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_338 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_169 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_337 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_169 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_338 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_169 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_337 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_169 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_169 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_169 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_169 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_169 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_169 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_336 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_168 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_335 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_168 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_336 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_168 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_335 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_168 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_168 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_168 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_168 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_168 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_168 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_334 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_167 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_333 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_167 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_334 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_167 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_333 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_167 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_167 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_167 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_167 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_167 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_167 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_332 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_166 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_331 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_166 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_332 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_166 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_331 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_166 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_166 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_166 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_166 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_166 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_166 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_330 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_165 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_329 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_165 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_330 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_165 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_329 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_165 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_165 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_165 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_165 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_165 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_165 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_328 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_164 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_327 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_164 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_328 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_164 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_327 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_164 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_164 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_164 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_164 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_164 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_164 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_326 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_163 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_325 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_163 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_326 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_163 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_325 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_163 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_163 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_163 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_163 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_163 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_163 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_324 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_162 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_323 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_162 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_324 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_162 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_323 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_162 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_162 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_162 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_162 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_162 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_162 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_322 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_161 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_321 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_161 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_322 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_161 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_321 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_161 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_161 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_161 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_161 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_161 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_161 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_320 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_160 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_319 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_160 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_320 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_160 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_319 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_160 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_160 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_160 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_160 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_160 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_160 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_318 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_159 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_317 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_159 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_318 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_159 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_317 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_159 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_159 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_159 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_159 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_159 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_159 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_316 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_158 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_315 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_158 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_316 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_158 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_315 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_158 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_158 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_158 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_158 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_158 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_158 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_314 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_157 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_313 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_157 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_314 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_157 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_313 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_157 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_157 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_157 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_157 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_157 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_157 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_312 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_156 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_311 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_156 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_312 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_156 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_311 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_156 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_156 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_156 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_156 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_156 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_156 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_310 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_155 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_309 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_155 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_310 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_155 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_309 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_155 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_155 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_155 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_155 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_155 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_155 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_308 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_154 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_307 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_154 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_308 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_154 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_307 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_154 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_154 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_154 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_154 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_154 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_154 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_306 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_153 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_305 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_153 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_306 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_153 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_305 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_153 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_153 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_153 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_153 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_153 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_153 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_304 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_152 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_303 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_152 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_304 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_152 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_303 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_152 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_152 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_152 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_152 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_152 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_152 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_302 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_151 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_301 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_151 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_302 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_151 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_301 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_151 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_151 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_151 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_151 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_151 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_151 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_300 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_150 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_299 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_150 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_300 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_150 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_299 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_150 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_150 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_150 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_150 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_150 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_150 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_298 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_149 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_297 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_149 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_298 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_149 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_297 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_149 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_149 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_149 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_149 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_149 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_149 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_296 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_148 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_295 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_148 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_296 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_148 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_295 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_148 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_148 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_148 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_148 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_148 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_148 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_294 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_147 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_293 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_147 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_294 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_147 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_293 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_147 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_147 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_147 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_147 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_147 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_147 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_292 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_146 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_291 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_146 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_292 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_146 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_291 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_146 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_146 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_146 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_146 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_146 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_146 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_290 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_145 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_289 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_145 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_290 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_145 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_289 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_145 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_145 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_145 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_145 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_145 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_145 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_288 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_144 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_287 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_144 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_288 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_144 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_287 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_144 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_144 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_144 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_144 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_144 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_144 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_286 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_143 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_285 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_143 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_286 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_143 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_285 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_143 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_143 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_143 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_143 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_143 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_143 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_284 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_142 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_283 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_142 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_284 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_142 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_283 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_142 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_142 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_142 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_142 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_142 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_142 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_282 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_141 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_281 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_141 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_282 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_141 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_281 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_141 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_141 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_141 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_141 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_141 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_141 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_280 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_140 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_279 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_140 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_280 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_140 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_279 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_140 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_140 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_140 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_140 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_140 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_140 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_278 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_139 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_277 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_139 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_278 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_139 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_277 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_139 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_139 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_139 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_139 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_139 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_139 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_276 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_138 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_275 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_138 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_276 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_138 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_275 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_138 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_138 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_138 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_138 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_138 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_138 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_274 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_137 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_273 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_137 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_274 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_137 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_273 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_137 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_137 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_137 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_137 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_137 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_137 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_272 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_136 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_271 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_136 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_272 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_136 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_271 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_136 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_136 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_136 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_136 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_136 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_136 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_270 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_135 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_269 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_135 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_270 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_135 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_269 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_135 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_135 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_135 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_135 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_135 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_135 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_268 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_134 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_267 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_134 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_268 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_134 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_267 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_134 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_134 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_134 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_134 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_134 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_134 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_266 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_133 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_265 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_133 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_266 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_133 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_265 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_133 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_133 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_133 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_133 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_133 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_133 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_264 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_132 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_263 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_132 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_264 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_132 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_263 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_132 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_132 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_132 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_132 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_132 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_132 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_262 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_131 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_261 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_131 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_262 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_131 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_261 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_131 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_131 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_131 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_131 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_131 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_131 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_260 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_130 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_259 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_130 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_260 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_130 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_259 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_130 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_130 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_130 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_130 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_130 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_130 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_258 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_129 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_257 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_129 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_258 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_129 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_257 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_129 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_129 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_129 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_129 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_129 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_129 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module reg_SDE_size128_0 ( clk, D0, D1, sel, Q );
  input [127:0] D0;
  input [127:0] D1;
  output [127:0] Q;
  input clk, sel;
  wire   n6, n7, n8, n9, n10;

  ff_SDE_0 Inst_ff_SDE_0 ( .clk(clk), .D0(D0[0]), .D1(D1[0]), .sel(n6), .Q(
        Q[0]) );
  ff_SDE_255 Inst_ff_SDE_1 ( .clk(clk), .D0(D0[1]), .D1(D1[1]), .sel(n7), .Q(
        Q[1]) );
  ff_SDE_254 Inst_ff_SDE_2 ( .clk(clk), .D0(D0[2]), .D1(D1[2]), .sel(n8), .Q(
        Q[2]) );
  ff_SDE_253 Inst_ff_SDE_3 ( .clk(clk), .D0(D0[3]), .D1(D1[3]), .sel(n9), .Q(
        Q[3]) );
  ff_SDE_252 Inst_ff_SDE_4 ( .clk(clk), .D0(D0[4]), .D1(D1[4]), .sel(n7), .Q(
        Q[4]) );
  ff_SDE_251 Inst_ff_SDE_5 ( .clk(clk), .D0(D0[5]), .D1(D1[5]), .sel(n6), .Q(
        Q[5]) );
  ff_SDE_250 Inst_ff_SDE_6 ( .clk(clk), .D0(D0[6]), .D1(D1[6]), .sel(n7), .Q(
        Q[6]) );
  ff_SDE_249 Inst_ff_SDE_7 ( .clk(clk), .D0(D0[7]), .D1(D1[7]), .sel(sel), .Q(
        Q[7]) );
  ff_SDE_248 Inst_ff_SDE_8 ( .clk(clk), .D0(D0[8]), .D1(D1[8]), .sel(n6), .Q(
        Q[8]) );
  ff_SDE_247 Inst_ff_SDE_9 ( .clk(clk), .D0(D0[9]), .D1(D1[9]), .sel(sel), .Q(
        Q[9]) );
  ff_SDE_246 Inst_ff_SDE_10 ( .clk(clk), .D0(D0[10]), .D1(D1[10]), .sel(sel), 
        .Q(Q[10]) );
  ff_SDE_245 Inst_ff_SDE_11 ( .clk(clk), .D0(D0[11]), .D1(D1[11]), .sel(sel), 
        .Q(Q[11]) );
  ff_SDE_244 Inst_ff_SDE_12 ( .clk(clk), .D0(D0[12]), .D1(D1[12]), .sel(sel), 
        .Q(Q[12]) );
  ff_SDE_243 Inst_ff_SDE_13 ( .clk(clk), .D0(D0[13]), .D1(D1[13]), .sel(sel), 
        .Q(Q[13]) );
  ff_SDE_242 Inst_ff_SDE_14 ( .clk(clk), .D0(D0[14]), .D1(D1[14]), .sel(sel), 
        .Q(Q[14]) );
  ff_SDE_241 Inst_ff_SDE_15 ( .clk(clk), .D0(D0[15]), .D1(D1[15]), .sel(sel), 
        .Q(Q[15]) );
  ff_SDE_240 Inst_ff_SDE_16 ( .clk(clk), .D0(D0[16]), .D1(D1[16]), .sel(sel), 
        .Q(Q[16]) );
  ff_SDE_239 Inst_ff_SDE_17 ( .clk(clk), .D0(D0[17]), .D1(D1[17]), .sel(sel), 
        .Q(Q[17]) );
  ff_SDE_238 Inst_ff_SDE_18 ( .clk(clk), .D0(D0[18]), .D1(D1[18]), .sel(sel), 
        .Q(Q[18]) );
  ff_SDE_237 Inst_ff_SDE_19 ( .clk(clk), .D0(D0[19]), .D1(D1[19]), .sel(sel), 
        .Q(Q[19]) );
  ff_SDE_236 Inst_ff_SDE_20 ( .clk(clk), .D0(D0[20]), .D1(D1[20]), .sel(n7), 
        .Q(Q[20]) );
  ff_SDE_235 Inst_ff_SDE_21 ( .clk(clk), .D0(D0[21]), .D1(D1[21]), .sel(n8), 
        .Q(Q[21]) );
  ff_SDE_234 Inst_ff_SDE_22 ( .clk(clk), .D0(D0[22]), .D1(D1[22]), .sel(n9), 
        .Q(Q[22]) );
  ff_SDE_233 Inst_ff_SDE_23 ( .clk(clk), .D0(D0[23]), .D1(D1[23]), .sel(n8), 
        .Q(Q[23]) );
  ff_SDE_232 Inst_ff_SDE_24 ( .clk(clk), .D0(D0[24]), .D1(D1[24]), .sel(n6), 
        .Q(Q[24]) );
  ff_SDE_231 Inst_ff_SDE_25 ( .clk(clk), .D0(D0[25]), .D1(D1[25]), .sel(n7), 
        .Q(Q[25]) );
  ff_SDE_230 Inst_ff_SDE_26 ( .clk(clk), .D0(D0[26]), .D1(D1[26]), .sel(n7), 
        .Q(Q[26]) );
  ff_SDE_229 Inst_ff_SDE_27 ( .clk(clk), .D0(D0[27]), .D1(D1[27]), .sel(sel), 
        .Q(Q[27]) );
  ff_SDE_228 Inst_ff_SDE_28 ( .clk(clk), .D0(D0[28]), .D1(D1[28]), .sel(sel), 
        .Q(Q[28]) );
  ff_SDE_227 Inst_ff_SDE_29 ( .clk(clk), .D0(D0[29]), .D1(D1[29]), .sel(sel), 
        .Q(Q[29]) );
  ff_SDE_226 Inst_ff_SDE_30 ( .clk(clk), .D0(D0[30]), .D1(D1[30]), .sel(sel), 
        .Q(Q[30]) );
  ff_SDE_225 Inst_ff_SDE_31 ( .clk(clk), .D0(D0[31]), .D1(D1[31]), .sel(sel), 
        .Q(Q[31]) );
  ff_SDE_224 Inst_ff_SDE_32 ( .clk(clk), .D0(D0[32]), .D1(D1[32]), .sel(n8), 
        .Q(Q[32]) );
  ff_SDE_223 Inst_ff_SDE_33 ( .clk(clk), .D0(D0[33]), .D1(D1[33]), .sel(n9), 
        .Q(Q[33]) );
  ff_SDE_222 Inst_ff_SDE_34 ( .clk(clk), .D0(D0[34]), .D1(D1[34]), .sel(n9), 
        .Q(Q[34]) );
  ff_SDE_221 Inst_ff_SDE_35 ( .clk(clk), .D0(D0[35]), .D1(D1[35]), .sel(n7), 
        .Q(Q[35]) );
  ff_SDE_220 Inst_ff_SDE_36 ( .clk(clk), .D0(D0[36]), .D1(D1[36]), .sel(n8), 
        .Q(Q[36]) );
  ff_SDE_219 Inst_ff_SDE_37 ( .clk(clk), .D0(D0[37]), .D1(D1[37]), .sel(n6), 
        .Q(Q[37]) );
  ff_SDE_218 Inst_ff_SDE_38 ( .clk(clk), .D0(D0[38]), .D1(D1[38]), .sel(sel), 
        .Q(Q[38]) );
  ff_SDE_217 Inst_ff_SDE_39 ( .clk(clk), .D0(D0[39]), .D1(D1[39]), .sel(sel), 
        .Q(Q[39]) );
  ff_SDE_216 Inst_ff_SDE_40 ( .clk(clk), .D0(D0[40]), .D1(D1[40]), .sel(sel), 
        .Q(Q[40]) );
  ff_SDE_215 Inst_ff_SDE_41 ( .clk(clk), .D0(D0[41]), .D1(D1[41]), .sel(sel), 
        .Q(Q[41]) );
  ff_SDE_214 Inst_ff_SDE_42 ( .clk(clk), .D0(D0[42]), .D1(D1[42]), .sel(sel), 
        .Q(Q[42]) );
  ff_SDE_213 Inst_ff_SDE_43 ( .clk(clk), .D0(D0[43]), .D1(D1[43]), .sel(sel), 
        .Q(Q[43]) );
  ff_SDE_212 Inst_ff_SDE_44 ( .clk(clk), .D0(D0[44]), .D1(D1[44]), .sel(n9), 
        .Q(Q[44]) );
  ff_SDE_211 Inst_ff_SDE_45 ( .clk(clk), .D0(D0[45]), .D1(D1[45]), .sel(n6), 
        .Q(Q[45]) );
  ff_SDE_210 Inst_ff_SDE_46 ( .clk(clk), .D0(D0[46]), .D1(D1[46]), .sel(n8), 
        .Q(Q[46]) );
  ff_SDE_209 Inst_ff_SDE_47 ( .clk(clk), .D0(D0[47]), .D1(D1[47]), .sel(n6), 
        .Q(Q[47]) );
  ff_SDE_208 Inst_ff_SDE_48 ( .clk(clk), .D0(D0[48]), .D1(D1[48]), .sel(sel), 
        .Q(Q[48]) );
  ff_SDE_207 Inst_ff_SDE_49 ( .clk(clk), .D0(D0[49]), .D1(D1[49]), .sel(sel), 
        .Q(Q[49]) );
  ff_SDE_206 Inst_ff_SDE_50 ( .clk(clk), .D0(D0[50]), .D1(D1[50]), .sel(sel), 
        .Q(Q[50]) );
  ff_SDE_205 Inst_ff_SDE_51 ( .clk(clk), .D0(D0[51]), .D1(D1[51]), .sel(sel), 
        .Q(Q[51]) );
  ff_SDE_204 Inst_ff_SDE_52 ( .clk(clk), .D0(D0[52]), .D1(D1[52]), .sel(n7), 
        .Q(Q[52]) );
  ff_SDE_203 Inst_ff_SDE_53 ( .clk(clk), .D0(D0[53]), .D1(D1[53]), .sel(n8), 
        .Q(Q[53]) );
  ff_SDE_202 Inst_ff_SDE_54 ( .clk(clk), .D0(D0[54]), .D1(D1[54]), .sel(n9), 
        .Q(Q[54]) );
  ff_SDE_201 Inst_ff_SDE_55 ( .clk(clk), .D0(D0[55]), .D1(D1[55]), .sel(n7), 
        .Q(Q[55]) );
  ff_SDE_200 Inst_ff_SDE_56 ( .clk(clk), .D0(D0[56]), .D1(D1[56]), .sel(n9), 
        .Q(Q[56]) );
  ff_SDE_199 Inst_ff_SDE_57 ( .clk(clk), .D0(D0[57]), .D1(D1[57]), .sel(n8), 
        .Q(Q[57]) );
  ff_SDE_198 Inst_ff_SDE_58 ( .clk(clk), .D0(D0[58]), .D1(D1[58]), .sel(n6), 
        .Q(Q[58]) );
  ff_SDE_197 Inst_ff_SDE_59 ( .clk(clk), .D0(D0[59]), .D1(D1[59]), .sel(n7), 
        .Q(Q[59]) );
  ff_SDE_196 Inst_ff_SDE_60 ( .clk(clk), .D0(D0[60]), .D1(D1[60]), .sel(n8), 
        .Q(Q[60]) );
  ff_SDE_195 Inst_ff_SDE_61 ( .clk(clk), .D0(D0[61]), .D1(D1[61]), .sel(n9), 
        .Q(Q[61]) );
  ff_SDE_194 Inst_ff_SDE_62 ( .clk(clk), .D0(D0[62]), .D1(D1[62]), .sel(n9), 
        .Q(Q[62]) );
  ff_SDE_193 Inst_ff_SDE_63 ( .clk(clk), .D0(D0[63]), .D1(D1[63]), .sel(n6), 
        .Q(Q[63]) );
  ff_SDE_192 Inst_ff_SDE_64 ( .clk(clk), .D0(D0[64]), .D1(D1[64]), .sel(n7), 
        .Q(Q[64]) );
  ff_SDE_191 Inst_ff_SDE_65 ( .clk(clk), .D0(D0[65]), .D1(D1[65]), .sel(n8), 
        .Q(Q[65]) );
  ff_SDE_190 Inst_ff_SDE_66 ( .clk(clk), .D0(D0[66]), .D1(D1[66]), .sel(n9), 
        .Q(Q[66]) );
  ff_SDE_189 Inst_ff_SDE_67 ( .clk(clk), .D0(D0[67]), .D1(D1[67]), .sel(n6), 
        .Q(Q[67]) );
  ff_SDE_188 Inst_ff_SDE_68 ( .clk(clk), .D0(D0[68]), .D1(D1[68]), .sel(n7), 
        .Q(Q[68]) );
  ff_SDE_187 Inst_ff_SDE_69 ( .clk(clk), .D0(D0[69]), .D1(D1[69]), .sel(n8), 
        .Q(Q[69]) );
  ff_SDE_186 Inst_ff_SDE_70 ( .clk(clk), .D0(D0[70]), .D1(D1[70]), .sel(n9), 
        .Q(Q[70]) );
  ff_SDE_185 Inst_ff_SDE_71 ( .clk(clk), .D0(D0[71]), .D1(D1[71]), .sel(n6), 
        .Q(Q[71]) );
  ff_SDE_184 Inst_ff_SDE_72 ( .clk(clk), .D0(D0[72]), .D1(D1[72]), .sel(n7), 
        .Q(Q[72]) );
  ff_SDE_183 Inst_ff_SDE_73 ( .clk(clk), .D0(D0[73]), .D1(D1[73]), .sel(n8), 
        .Q(Q[73]) );
  ff_SDE_182 Inst_ff_SDE_74 ( .clk(clk), .D0(D0[74]), .D1(D1[74]), .sel(n9), 
        .Q(Q[74]) );
  ff_SDE_181 Inst_ff_SDE_75 ( .clk(clk), .D0(D0[75]), .D1(D1[75]), .sel(n6), 
        .Q(Q[75]) );
  ff_SDE_180 Inst_ff_SDE_76 ( .clk(clk), .D0(D0[76]), .D1(D1[76]), .sel(n7), 
        .Q(Q[76]) );
  ff_SDE_179 Inst_ff_SDE_77 ( .clk(clk), .D0(D0[77]), .D1(D1[77]), .sel(n8), 
        .Q(Q[77]) );
  ff_SDE_178 Inst_ff_SDE_78 ( .clk(clk), .D0(D0[78]), .D1(D1[78]), .sel(n9), 
        .Q(Q[78]) );
  ff_SDE_177 Inst_ff_SDE_79 ( .clk(clk), .D0(D0[79]), .D1(D1[79]), .sel(n6), 
        .Q(Q[79]) );
  ff_SDE_176 Inst_ff_SDE_80 ( .clk(clk), .D0(D0[80]), .D1(D1[80]), .sel(n9), 
        .Q(Q[80]) );
  ff_SDE_175 Inst_ff_SDE_81 ( .clk(clk), .D0(D0[81]), .D1(D1[81]), .sel(n9), 
        .Q(Q[81]) );
  ff_SDE_174 Inst_ff_SDE_82 ( .clk(clk), .D0(D0[82]), .D1(D1[82]), .sel(n9), 
        .Q(Q[82]) );
  ff_SDE_173 Inst_ff_SDE_83 ( .clk(clk), .D0(D0[83]), .D1(D1[83]), .sel(n9), 
        .Q(Q[83]) );
  ff_SDE_172 Inst_ff_SDE_84 ( .clk(clk), .D0(D0[84]), .D1(D1[84]), .sel(n9), 
        .Q(Q[84]) );
  ff_SDE_171 Inst_ff_SDE_85 ( .clk(clk), .D0(D0[85]), .D1(D1[85]), .sel(n9), 
        .Q(Q[85]) );
  ff_SDE_170 Inst_ff_SDE_86 ( .clk(clk), .D0(D0[86]), .D1(D1[86]), .sel(n9), 
        .Q(Q[86]) );
  ff_SDE_169 Inst_ff_SDE_87 ( .clk(clk), .D0(D0[87]), .D1(D1[87]), .sel(n9), 
        .Q(Q[87]) );
  ff_SDE_168 Inst_ff_SDE_88 ( .clk(clk), .D0(D0[88]), .D1(D1[88]), .sel(n9), 
        .Q(Q[88]) );
  ff_SDE_167 Inst_ff_SDE_89 ( .clk(clk), .D0(D0[89]), .D1(D1[89]), .sel(n9), 
        .Q(Q[89]) );
  ff_SDE_166 Inst_ff_SDE_90 ( .clk(clk), .D0(D0[90]), .D1(D1[90]), .sel(n9), 
        .Q(Q[90]) );
  ff_SDE_165 Inst_ff_SDE_91 ( .clk(clk), .D0(D0[91]), .D1(D1[91]), .sel(n9), 
        .Q(Q[91]) );
  ff_SDE_164 Inst_ff_SDE_92 ( .clk(clk), .D0(D0[92]), .D1(D1[92]), .sel(n8), 
        .Q(Q[92]) );
  ff_SDE_163 Inst_ff_SDE_93 ( .clk(clk), .D0(D0[93]), .D1(D1[93]), .sel(n8), 
        .Q(Q[93]) );
  ff_SDE_162 Inst_ff_SDE_94 ( .clk(clk), .D0(D0[94]), .D1(D1[94]), .sel(n8), 
        .Q(Q[94]) );
  ff_SDE_161 Inst_ff_SDE_95 ( .clk(clk), .D0(D0[95]), .D1(D1[95]), .sel(n8), 
        .Q(Q[95]) );
  ff_SDE_160 Inst_ff_SDE_96 ( .clk(clk), .D0(D0[96]), .D1(D1[96]), .sel(n8), 
        .Q(Q[96]) );
  ff_SDE_159 Inst_ff_SDE_97 ( .clk(clk), .D0(D0[97]), .D1(D1[97]), .sel(n8), 
        .Q(Q[97]) );
  ff_SDE_158 Inst_ff_SDE_98 ( .clk(clk), .D0(D0[98]), .D1(D1[98]), .sel(n8), 
        .Q(Q[98]) );
  ff_SDE_157 Inst_ff_SDE_99 ( .clk(clk), .D0(D0[99]), .D1(D1[99]), .sel(n8), 
        .Q(Q[99]) );
  ff_SDE_156 Inst_ff_SDE_100 ( .clk(clk), .D0(D0[100]), .D1(D1[100]), .sel(n8), 
        .Q(Q[100]) );
  ff_SDE_155 Inst_ff_SDE_101 ( .clk(clk), .D0(D0[101]), .D1(D1[101]), .sel(n8), 
        .Q(Q[101]) );
  ff_SDE_154 Inst_ff_SDE_102 ( .clk(clk), .D0(D0[102]), .D1(D1[102]), .sel(n8), 
        .Q(Q[102]) );
  ff_SDE_153 Inst_ff_SDE_103 ( .clk(clk), .D0(D0[103]), .D1(D1[103]), .sel(n8), 
        .Q(Q[103]) );
  ff_SDE_152 Inst_ff_SDE_104 ( .clk(clk), .D0(D0[104]), .D1(D1[104]), .sel(n7), 
        .Q(Q[104]) );
  ff_SDE_151 Inst_ff_SDE_105 ( .clk(clk), .D0(D0[105]), .D1(D1[105]), .sel(n7), 
        .Q(Q[105]) );
  ff_SDE_150 Inst_ff_SDE_106 ( .clk(clk), .D0(D0[106]), .D1(D1[106]), .sel(n7), 
        .Q(Q[106]) );
  ff_SDE_149 Inst_ff_SDE_107 ( .clk(clk), .D0(D0[107]), .D1(D1[107]), .sel(n7), 
        .Q(Q[107]) );
  ff_SDE_148 Inst_ff_SDE_108 ( .clk(clk), .D0(D0[108]), .D1(D1[108]), .sel(n7), 
        .Q(Q[108]) );
  ff_SDE_147 Inst_ff_SDE_109 ( .clk(clk), .D0(D0[109]), .D1(D1[109]), .sel(n7), 
        .Q(Q[109]) );
  ff_SDE_146 Inst_ff_SDE_110 ( .clk(clk), .D0(D0[110]), .D1(D1[110]), .sel(n7), 
        .Q(Q[110]) );
  ff_SDE_145 Inst_ff_SDE_111 ( .clk(clk), .D0(D0[111]), .D1(D1[111]), .sel(n7), 
        .Q(Q[111]) );
  ff_SDE_144 Inst_ff_SDE_112 ( .clk(clk), .D0(D0[112]), .D1(D1[112]), .sel(n7), 
        .Q(Q[112]) );
  ff_SDE_143 Inst_ff_SDE_113 ( .clk(clk), .D0(D0[113]), .D1(D1[113]), .sel(n7), 
        .Q(Q[113]) );
  ff_SDE_142 Inst_ff_SDE_114 ( .clk(clk), .D0(D0[114]), .D1(D1[114]), .sel(n7), 
        .Q(Q[114]) );
  ff_SDE_141 Inst_ff_SDE_115 ( .clk(clk), .D0(D0[115]), .D1(D1[115]), .sel(n7), 
        .Q(Q[115]) );
  ff_SDE_140 Inst_ff_SDE_116 ( .clk(clk), .D0(D0[116]), .D1(D1[116]), .sel(n6), 
        .Q(Q[116]) );
  ff_SDE_139 Inst_ff_SDE_117 ( .clk(clk), .D0(D0[117]), .D1(D1[117]), .sel(n6), 
        .Q(Q[117]) );
  ff_SDE_138 Inst_ff_SDE_118 ( .clk(clk), .D0(D0[118]), .D1(D1[118]), .sel(n6), 
        .Q(Q[118]) );
  ff_SDE_137 Inst_ff_SDE_119 ( .clk(clk), .D0(D0[119]), .D1(D1[119]), .sel(n6), 
        .Q(Q[119]) );
  ff_SDE_136 Inst_ff_SDE_120 ( .clk(clk), .D0(D0[120]), .D1(D1[120]), .sel(n6), 
        .Q(Q[120]) );
  ff_SDE_135 Inst_ff_SDE_121 ( .clk(clk), .D0(D0[121]), .D1(D1[121]), .sel(n6), 
        .Q(Q[121]) );
  ff_SDE_134 Inst_ff_SDE_122 ( .clk(clk), .D0(D0[122]), .D1(D1[122]), .sel(n6), 
        .Q(Q[122]) );
  ff_SDE_133 Inst_ff_SDE_123 ( .clk(clk), .D0(D0[123]), .D1(D1[123]), .sel(n6), 
        .Q(Q[123]) );
  ff_SDE_132 Inst_ff_SDE_124 ( .clk(clk), .D0(D0[124]), .D1(D1[124]), .sel(n6), 
        .Q(Q[124]) );
  ff_SDE_131 Inst_ff_SDE_125 ( .clk(clk), .D0(D0[125]), .D1(D1[125]), .sel(n6), 
        .Q(Q[125]) );
  ff_SDE_130 Inst_ff_SDE_126 ( .clk(clk), .D0(D0[126]), .D1(D1[126]), .sel(n6), 
        .Q(Q[126]) );
  ff_SDE_129 Inst_ff_SDE_127 ( .clk(clk), .D0(D0[127]), .D1(D1[127]), .sel(n6), 
        .Q(Q[127]) );
  INV_X1 U1 ( .A(n10), .ZN(n6) );
  INV_X1 U2 ( .A(n10), .ZN(n7) );
  INV_X1 U3 ( .A(n10), .ZN(n8) );
  INV_X1 U4 ( .A(n10), .ZN(n9) );
  INV_X1 U5 ( .A(sel), .ZN(n10) );
endmodule


module MyXOR_0 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1799 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1798 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1797 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1796 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1795 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1794 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1793 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1792 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1791 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1790 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1789 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1788 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1787 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1786 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1785 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1784 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1783 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1782 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1781 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1780 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1779 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1778 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1777 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1776 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1775 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1774 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_0 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_679 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1773 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_678 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1772 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_677 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_676 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1771 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_675 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1770 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_674 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_673 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1769 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_672 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1768 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1767 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1766 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1765 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1764 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1763 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1762 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1761 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1760 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1759 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_671 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1758 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1757 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1756 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_670 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_669 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_668 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_667 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1755 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_666 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_665 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1754 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1753 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1752 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1751 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1750 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1749 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1748 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1747 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1746 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1745 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_664 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_663 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_662 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_661 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_660 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_659 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_658 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_657 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_656 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_655 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_654 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_653 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_652 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_651 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_650 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_649 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_648 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_647 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1744 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1743 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1742 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1741 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1740 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1739 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1738 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1737 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1736 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1735 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1734 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1733 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1732 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1731 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1730 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1729 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1728 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1727 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1726 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1725 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1724 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1723 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1722 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1721 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1720 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1719 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1718 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1717 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1716 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1715 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1714 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_0 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_79 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_1713 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1712 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1711 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_78 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_77 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_0 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_0 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_1799 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_1798 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_1797 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_1796 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_1795 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_1794 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_1793 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_1792 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_1791 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_1790 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_1789 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_1788 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_1787 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_1786 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_1785 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_1784 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_1783 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_1782 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_1781 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_1780 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_1779 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_1778 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_1777 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_1776 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_1775 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_1774 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_0 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_679 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_1773 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_678 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_1772 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_677 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_676 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_1771 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_675 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_1770 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_674 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_673 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_1769 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_672 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_1768 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_1767 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_1766 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_1765 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_1764 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_1763 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_1762 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_1761 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_1760 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_1759 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_671 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_1758 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_1757 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_1756 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_670 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_669 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_668 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_667 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_1755 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_666 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_665 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_1754 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_1753 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_1752 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_1751 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_1750 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_1749 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_1748 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_1747 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_1746 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_1745 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_664 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_663 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_662 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_661 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_660 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_659 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_658 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_657 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_656 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_655 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_654 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_653 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_652 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_651 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_650 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_649 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_648 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_647 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_1744 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_1743 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_1742 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_1741 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_1740 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_1739 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_1738 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_1737 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_1736 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_1735 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_1734 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_1733 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_1732 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_1731 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_1730 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_1729 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_1728 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_1727 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_1726 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_1725 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_1724 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_1723 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_1722 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_1721 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_1720 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_1719 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_1718 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_1717 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_1716 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_1715 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_1714 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_0 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_79 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_1713 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_1712 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_1711 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_78 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_77 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_1710 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1709 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1708 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1707 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1706 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1705 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1704 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1703 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1702 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1701 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1700 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1699 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1698 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1697 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1696 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1695 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1694 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1693 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1692 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1691 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1690 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1689 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1688 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1687 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1686 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1685 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1684 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_646 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_645 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1683 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_644 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1682 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_643 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_642 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1681 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_641 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1680 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_640 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_639 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1679 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_638 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1678 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1677 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1676 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1675 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1674 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1673 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1672 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1671 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1670 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1669 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_637 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1668 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1667 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1666 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_636 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_635 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_634 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_633 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1665 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_632 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_631 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1664 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1663 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1662 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1661 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1660 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1659 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1658 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1657 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1656 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1655 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_630 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_629 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_628 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_627 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_626 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_625 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_624 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_623 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_622 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_621 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_620 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_619 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_618 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_617 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_616 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_615 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_614 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_613 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1654 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1653 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1652 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1651 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1650 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1649 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1648 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1647 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1646 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1645 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1644 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1643 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1642 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1641 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1640 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1639 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1638 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1637 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1636 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1635 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1634 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1633 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1632 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1631 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1630 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1629 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1628 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1627 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1626 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1625 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1624 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_76 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_75 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_1623 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1622 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1621 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_74 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_73 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_19 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_1710 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_1709 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_1708 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_1707 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_1706 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_1705 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_1704 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_1703 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_1702 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_1701 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_1700 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_1699 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_1698 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_1697 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_1696 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_1695 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_1694 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_1693 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_1692 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_1691 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_1690 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_1689 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_1688 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_1687 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_1686 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_1685 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_1684 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_646 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_645 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_1683 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_644 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_1682 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_643 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_642 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_1681 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_641 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_1680 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_640 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_639 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_1679 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_638 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_1678 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_1677 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_1676 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_1675 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_1674 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_1673 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_1672 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_1671 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_1670 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_1669 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_637 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_1668 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_1667 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_1666 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_636 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_635 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_634 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_633 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_1665 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_632 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_631 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_1664 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_1663 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_1662 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_1661 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_1660 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_1659 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_1658 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_1657 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_1656 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_1655 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_630 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_629 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_628 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_627 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_626 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_625 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_624 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_623 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_622 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_621 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_620 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_619 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_618 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_617 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_616 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_615 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_614 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_613 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_1654 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_1653 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_1652 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_1651 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_1650 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_1649 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_1648 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_1647 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_1646 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_1645 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_1644 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_1643 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_1642 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_1641 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_1640 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_1639 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_1638 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_1637 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_1636 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_1635 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_1634 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_1633 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_1632 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_1631 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_1630 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_1629 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_1628 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_1627 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_1626 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_1625 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_1624 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_76 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_75 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_1623 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_1622 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_1621 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_74 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_73 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_1620 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1619 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1618 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1617 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1616 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1615 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1614 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1613 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1612 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1611 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1610 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1609 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1608 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1607 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1606 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1605 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1604 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1603 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1602 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1601 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1600 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1599 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1598 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1597 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1596 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1595 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1594 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_612 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_611 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1593 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_610 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1592 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_609 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_608 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1591 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_607 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1590 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_606 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_605 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1589 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_604 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1588 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1587 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1586 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1585 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1584 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1583 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1582 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1581 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1580 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1579 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_603 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1578 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1577 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1576 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_602 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_601 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_600 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_599 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1575 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_598 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_597 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1574 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1573 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1572 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1571 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1570 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1569 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1568 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1567 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1566 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1565 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_596 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_595 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_594 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_593 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_592 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_591 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_590 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_589 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_588 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_587 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_586 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_585 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_584 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_583 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_582 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_581 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_580 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_579 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1564 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1563 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1562 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1561 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1560 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1559 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1558 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1557 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1556 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1555 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1554 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1553 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1552 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1551 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1550 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1549 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1548 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1547 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1546 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1545 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1544 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1543 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1542 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1541 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1540 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1539 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1538 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1537 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1536 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1535 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1534 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_72 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_71 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_1533 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1532 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1531 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_70 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_69 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_18 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_1620 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_1619 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_1618 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_1617 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_1616 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_1615 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_1614 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_1613 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_1612 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_1611 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_1610 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_1609 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_1608 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_1607 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_1606 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_1605 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_1604 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_1603 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_1602 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_1601 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_1600 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_1599 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_1598 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_1597 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_1596 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_1595 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_1594 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_612 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_611 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_1593 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_610 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_1592 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_609 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_608 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_1591 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_607 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_1590 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_606 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_605 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_1589 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_604 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_1588 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_1587 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_1586 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_1585 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_1584 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_1583 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_1582 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_1581 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_1580 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_1579 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_603 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_1578 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_1577 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_1576 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_602 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_601 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_600 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_599 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_1575 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_598 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_597 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_1574 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_1573 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_1572 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_1571 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_1570 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_1569 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_1568 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_1567 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_1566 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_1565 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_596 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_595 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_594 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_593 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_592 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_591 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_590 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_589 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_588 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_587 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_586 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_585 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_584 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_583 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_582 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_581 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_580 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_579 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_1564 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_1563 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_1562 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_1561 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_1560 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_1559 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_1558 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_1557 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_1556 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_1555 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_1554 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_1553 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_1552 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_1551 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_1550 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_1549 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_1548 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_1547 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_1546 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_1545 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_1544 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_1543 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_1542 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_1541 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_1540 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_1539 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_1538 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_1537 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_1536 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_1535 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_1534 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_72 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_71 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_1533 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_1532 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_1531 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_70 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_69 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_1530 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1529 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1528 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1527 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1526 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1525 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1524 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1523 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1522 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1521 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1520 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1519 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1518 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1517 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1516 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1515 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1514 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1513 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1512 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1511 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1510 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1509 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1508 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1507 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1506 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1505 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1504 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_578 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_577 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1503 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_576 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1502 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_575 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_574 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1501 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_573 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1500 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_572 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_571 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1499 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_570 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1498 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1497 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1496 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1495 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1494 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1493 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1492 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1491 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1490 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1489 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_569 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1488 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1487 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1486 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_568 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_567 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_566 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_565 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1485 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_564 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_563 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1484 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1483 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1482 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1481 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1480 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1479 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1478 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1477 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1476 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1475 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_562 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_561 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_560 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_559 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_558 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_557 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_556 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_555 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_554 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_553 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_552 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_551 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_550 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_549 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_548 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_547 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_546 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_545 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1474 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1473 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1472 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1471 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1470 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1469 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1468 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1467 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1466 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1465 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1464 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1463 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1462 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1461 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1460 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1459 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1458 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1457 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1456 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1455 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1454 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1453 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1452 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1451 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1450 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1449 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1448 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1447 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1446 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1445 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1444 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_68 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_67 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_1443 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1442 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1441 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_66 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_65 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_17 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_1530 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_1529 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_1528 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_1527 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_1526 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_1525 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_1524 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_1523 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_1522 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_1521 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_1520 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_1519 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_1518 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_1517 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_1516 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_1515 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_1514 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_1513 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_1512 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_1511 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_1510 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_1509 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_1508 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_1507 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_1506 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_1505 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_1504 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_578 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_577 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_1503 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_576 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_1502 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_575 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_574 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_1501 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_573 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_1500 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_572 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_571 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_1499 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_570 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_1498 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_1497 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_1496 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_1495 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_1494 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_1493 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_1492 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_1491 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_1490 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_1489 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_569 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_1488 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_1487 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_1486 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_568 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_567 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_566 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_565 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_1485 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_564 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_563 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_1484 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_1483 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_1482 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_1481 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_1480 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_1479 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_1478 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_1477 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_1476 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_1475 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_562 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_561 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_560 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_559 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_558 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_557 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_556 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_555 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_554 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_553 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_552 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_551 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_550 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_549 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_548 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_547 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_546 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_545 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_1474 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_1473 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_1472 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_1471 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_1470 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_1469 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_1468 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_1467 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_1466 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_1465 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_1464 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_1463 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_1462 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_1461 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_1460 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_1459 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_1458 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_1457 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_1456 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_1455 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_1454 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_1453 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_1452 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_1451 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_1450 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_1449 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_1448 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_1447 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_1446 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_1445 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_1444 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_68 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_67 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_1443 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_1442 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_1441 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_66 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_65 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_1440 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1439 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1438 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1437 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1436 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1435 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1434 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1433 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1432 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1431 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1430 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1429 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1428 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1427 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1426 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1425 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1424 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1423 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1422 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1421 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1420 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1419 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1418 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1417 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1416 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1415 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1414 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_544 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_543 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1413 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_542 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1412 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_541 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_540 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1411 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_539 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1410 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_538 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_537 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1409 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_536 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1408 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1407 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1406 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1405 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1404 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1403 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1402 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1401 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1400 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1399 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_535 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1398 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1397 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1396 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_534 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_533 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_532 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_531 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1395 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_530 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_529 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1394 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1393 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1392 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1391 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1390 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1389 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1388 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1387 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1386 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1385 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_528 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_527 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_526 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_525 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_524 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_523 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_522 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_521 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_520 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_519 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_518 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_517 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_516 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_515 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_514 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_513 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_512 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_511 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1384 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1383 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1382 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1381 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1380 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1379 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1378 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1377 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1376 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1375 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1374 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1373 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1372 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1371 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1370 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1369 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1368 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1367 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1366 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1365 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1364 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1363 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1362 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1361 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1360 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1359 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1358 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1357 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1356 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1355 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1354 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_64 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_63 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_1353 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1352 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1351 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_62 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_61 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_16 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_1440 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_1439 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_1438 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_1437 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_1436 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_1435 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_1434 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_1433 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_1432 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_1431 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_1430 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_1429 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_1428 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_1427 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_1426 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_1425 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_1424 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_1423 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_1422 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_1421 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_1420 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_1419 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_1418 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_1417 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_1416 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_1415 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_1414 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_544 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_543 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_1413 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_542 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_1412 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_541 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_540 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_1411 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_539 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_1410 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_538 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_537 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_1409 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_536 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_1408 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_1407 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_1406 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_1405 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_1404 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_1403 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_1402 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_1401 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_1400 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_1399 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_535 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_1398 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_1397 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_1396 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_534 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_533 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_532 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_531 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_1395 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_530 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_529 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_1394 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_1393 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_1392 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_1391 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_1390 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_1389 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_1388 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_1387 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_1386 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_1385 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_528 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_527 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_526 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_525 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_524 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_523 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_522 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_521 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_520 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_519 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_518 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_517 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_516 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_515 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_514 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_513 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_512 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_511 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_1384 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_1383 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_1382 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_1381 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_1380 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_1379 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_1378 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_1377 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_1376 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_1375 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_1374 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_1373 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_1372 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_1371 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_1370 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_1369 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_1368 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_1367 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_1366 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_1365 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_1364 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_1363 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_1362 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_1361 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_1360 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_1359 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_1358 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_1357 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_1356 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_1355 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_1354 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_64 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_63 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_1353 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_1352 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_1351 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_62 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_61 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_1350 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1349 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1348 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1347 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1346 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1345 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1344 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1343 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1342 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1341 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1340 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1339 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1338 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1337 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1336 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1335 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1334 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1333 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1332 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1331 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1330 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1329 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1328 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1327 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1326 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1325 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1324 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_510 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_509 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1323 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_508 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1322 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_507 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_506 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1321 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_505 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1320 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_504 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_503 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1319 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_502 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1318 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1317 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1316 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1315 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1314 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1313 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1312 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1311 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1310 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1309 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_501 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1308 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1307 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1306 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_500 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_499 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_498 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_497 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1305 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_496 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_495 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1304 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1303 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1302 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1301 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1300 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1299 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1298 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1297 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1296 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1295 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_494 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_493 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_492 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_491 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_490 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_489 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_488 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_487 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_486 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_485 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_484 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_483 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_482 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_481 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_480 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_479 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_478 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_477 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1294 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1293 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1292 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1291 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1290 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1289 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1288 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1287 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1286 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1285 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1284 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1283 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1282 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1281 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1280 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1279 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1278 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1277 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1276 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1275 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1274 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1273 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1272 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1271 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1270 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1269 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1268 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1267 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1266 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1265 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1264 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_60 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_59 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_1263 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1262 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1261 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_58 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_57 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_15 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_1350 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_1349 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_1348 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_1347 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_1346 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_1345 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_1344 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_1343 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_1342 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_1341 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_1340 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_1339 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_1338 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_1337 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_1336 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_1335 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_1334 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_1333 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_1332 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_1331 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_1330 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_1329 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_1328 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_1327 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_1326 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_1325 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_1324 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_510 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_509 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_1323 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_508 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_1322 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_507 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_506 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_1321 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_505 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_1320 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_504 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_503 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_1319 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_502 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_1318 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_1317 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_1316 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_1315 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_1314 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_1313 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_1312 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_1311 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_1310 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_1309 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_501 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_1308 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_1307 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_1306 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_500 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_499 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_498 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_497 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_1305 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_496 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_495 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_1304 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_1303 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_1302 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_1301 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_1300 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_1299 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_1298 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_1297 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_1296 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_1295 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_494 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_493 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_492 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_491 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_490 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_489 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_488 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_487 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_486 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_485 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_484 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_483 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_482 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_481 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_480 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_479 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_478 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_477 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_1294 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_1293 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_1292 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_1291 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_1290 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_1289 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_1288 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_1287 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_1286 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_1285 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_1284 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_1283 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_1282 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_1281 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_1280 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_1279 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_1278 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_1277 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_1276 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_1275 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_1274 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_1273 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_1272 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_1271 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_1270 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_1269 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_1268 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_1267 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_1266 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_1265 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_1264 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_60 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_59 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_1263 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_1262 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_1261 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_58 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_57 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_1260 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1259 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1258 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1257 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1256 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1255 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1254 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1253 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1252 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1251 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1250 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1249 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1248 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1247 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1246 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1245 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1244 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1243 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1242 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1241 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1240 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1239 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1238 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1237 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1236 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1235 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1234 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_476 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_475 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1233 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_474 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1232 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_473 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_472 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1231 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_471 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1230 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_470 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_469 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1229 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_468 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1228 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1227 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1226 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1225 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1224 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1223 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1222 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1221 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1220 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1219 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_467 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1218 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1217 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1216 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_466 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_465 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_464 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_463 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1215 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_462 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_461 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1214 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1213 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1212 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1211 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1210 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1209 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1208 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1207 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1206 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1205 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_460 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_459 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_458 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_457 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_456 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_455 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_454 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_453 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_452 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_451 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_450 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_449 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_448 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_447 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_446 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_445 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_444 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_443 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1204 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1203 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1202 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1201 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1200 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1199 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1198 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1197 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1196 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1195 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1194 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1193 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1192 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1191 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1190 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1189 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1188 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1187 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1186 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1185 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1184 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1183 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1182 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1181 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1180 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1179 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1178 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1177 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1176 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1175 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1174 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_56 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_55 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_1173 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1172 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1171 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_54 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_53 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_14 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_1260 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_1259 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_1258 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_1257 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_1256 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_1255 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_1254 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_1253 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_1252 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_1251 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_1250 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_1249 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_1248 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_1247 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_1246 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_1245 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_1244 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_1243 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_1242 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_1241 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_1240 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_1239 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_1238 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_1237 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_1236 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_1235 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_1234 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_476 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_475 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_1233 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_474 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_1232 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_473 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_472 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_1231 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_471 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_1230 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_470 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_469 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_1229 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_468 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_1228 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_1227 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_1226 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_1225 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_1224 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_1223 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_1222 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_1221 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_1220 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_1219 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_467 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_1218 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_1217 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_1216 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_466 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_465 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_464 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_463 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_1215 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_462 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_461 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_1214 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_1213 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_1212 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_1211 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_1210 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_1209 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_1208 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_1207 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_1206 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_1205 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_460 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_459 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_458 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_457 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_456 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_455 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_454 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_453 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_452 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_451 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_450 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_449 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_448 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_447 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_446 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_445 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_444 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_443 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_1204 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_1203 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_1202 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_1201 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_1200 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_1199 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_1198 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_1197 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_1196 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_1195 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_1194 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_1193 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_1192 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_1191 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_1190 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_1189 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_1188 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_1187 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_1186 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_1185 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_1184 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_1183 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_1182 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_1181 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_1180 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_1179 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_1178 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_1177 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_1176 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_1175 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_1174 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_56 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_55 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_1173 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_1172 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_1171 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_54 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_53 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_1170 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1169 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1168 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1167 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1166 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1165 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1164 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1163 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1162 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1161 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1160 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1159 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1158 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1157 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1156 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1155 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1154 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1153 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1152 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1151 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1150 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1149 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1148 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1147 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1146 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1145 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1144 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_442 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_441 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1143 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_440 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1142 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_439 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_438 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1141 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_437 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1140 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_436 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_435 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1139 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_434 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1138 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1137 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1136 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1135 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1134 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1133 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1132 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1131 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1130 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1129 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_433 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1128 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1127 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1126 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_432 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_431 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_430 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_429 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1125 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_428 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_427 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1124 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1123 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1122 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1121 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1120 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1119 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1118 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1117 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1116 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1115 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_426 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_425 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_424 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_423 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_422 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_421 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_420 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_419 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_418 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_417 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_416 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_415 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_414 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_413 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_412 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_411 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_410 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_409 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1114 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1113 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1112 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1111 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1110 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1109 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1108 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1107 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1106 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1105 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1104 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1103 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1102 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1101 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1100 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1099 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1098 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1097 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1096 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1095 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1094 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1093 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1092 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1091 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1090 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1089 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1088 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1087 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1086 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1085 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1084 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_52 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_51 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_1083 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1082 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1081 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_50 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_49 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_13 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_1170 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_1169 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_1168 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_1167 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_1166 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_1165 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_1164 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_1163 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_1162 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_1161 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_1160 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_1159 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_1158 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_1157 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_1156 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_1155 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_1154 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_1153 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_1152 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_1151 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_1150 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_1149 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_1148 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_1147 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_1146 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_1145 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_1144 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_442 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_441 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_1143 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_440 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_1142 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_439 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_438 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_1141 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_437 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_1140 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_436 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_435 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_1139 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_434 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_1138 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_1137 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_1136 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_1135 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_1134 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_1133 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_1132 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_1131 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_1130 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_1129 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_433 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_1128 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_1127 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_1126 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_432 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_431 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_430 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_429 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_1125 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_428 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_427 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_1124 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_1123 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_1122 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_1121 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_1120 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_1119 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_1118 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_1117 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_1116 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_1115 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_426 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_425 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_424 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_423 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_422 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_421 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_420 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_419 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_418 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_417 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_416 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_415 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_414 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_413 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_412 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_411 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_410 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_409 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_1114 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_1113 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_1112 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_1111 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_1110 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_1109 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_1108 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_1107 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_1106 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_1105 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_1104 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_1103 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_1102 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_1101 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_1100 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_1099 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_1098 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_1097 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_1096 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_1095 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_1094 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_1093 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_1092 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_1091 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_1090 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_1089 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_1088 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_1087 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_1086 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_1085 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_1084 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_52 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_51 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_1083 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_1082 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_1081 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_50 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_49 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_1080 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1079 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1078 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1077 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1076 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1075 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1074 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1073 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1072 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1071 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1070 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1069 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1068 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1067 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1066 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1065 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1064 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1063 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1062 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1061 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1060 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1059 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1058 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1057 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1056 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1055 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1054 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_408 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_407 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1053 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_406 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1052 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_405 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_404 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1051 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_403 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1050 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_402 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_401 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1049 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_400 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1048 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1047 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1046 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1045 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1044 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1043 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1042 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1041 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1040 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1039 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_399 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1038 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1037 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1036 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_398 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_397 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_396 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_395 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1035 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_394 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_393 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1034 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1033 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1032 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1031 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1030 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1029 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1028 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1027 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1026 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1025 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_392 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_391 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_390 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_389 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_388 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_387 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_386 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_385 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_384 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_383 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_382 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_381 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_380 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_379 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_378 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_377 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_376 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_375 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_1024 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1023 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1022 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1021 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1020 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1019 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1018 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1017 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1016 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1015 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1014 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1013 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1012 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1011 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1010 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1009 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1008 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1007 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1006 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1005 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1004 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1003 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1002 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1001 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1000 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_999 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_998 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_997 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_996 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_995 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_994 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_48 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_47 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_993 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_992 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_991 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_46 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_45 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_12 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_1080 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_1079 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_1078 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_1077 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_1076 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_1075 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_1074 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_1073 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_1072 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_1071 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_1070 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_1069 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_1068 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_1067 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_1066 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_1065 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_1064 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_1063 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_1062 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_1061 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_1060 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_1059 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_1058 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_1057 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_1056 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_1055 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_1054 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_408 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_407 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_1053 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_406 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_1052 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_405 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_404 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_1051 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_403 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_1050 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_402 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_401 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_1049 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_400 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_1048 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_1047 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_1046 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_1045 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_1044 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_1043 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_1042 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_1041 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_1040 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_1039 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_399 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_1038 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_1037 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_1036 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_398 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_397 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_396 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_395 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_1035 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_394 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_393 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_1034 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_1033 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_1032 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_1031 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_1030 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_1029 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_1028 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_1027 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_1026 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_1025 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_392 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_391 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_390 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_389 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_388 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_387 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_386 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_385 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_384 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_383 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_382 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_381 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_380 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_379 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_378 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_377 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_376 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_375 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_1024 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_1023 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_1022 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_1021 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_1020 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_1019 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_1018 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_1017 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_1016 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_1015 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_1014 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_1013 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_1012 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_1011 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_1010 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_1009 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_1008 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_1007 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_1006 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_1005 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_1004 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_1003 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_1002 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_1001 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_1000 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_999 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_998 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_997 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_996 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_995 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_994 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_48 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_47 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_993 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_992 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_991 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_46 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_45 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_990 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_989 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_988 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_987 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_986 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_985 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_984 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_983 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_982 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_981 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_980 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_979 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_978 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_977 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_976 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_975 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_974 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_973 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_972 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_971 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_970 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_969 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_968 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_967 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_966 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_965 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_964 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_374 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_373 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_963 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_372 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_962 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_371 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_370 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_961 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_369 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_960 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_368 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_367 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_959 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_366 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_958 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_957 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_956 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_955 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_954 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_953 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_952 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_951 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_950 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_949 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_365 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_948 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_947 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_946 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_364 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_363 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_362 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_361 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_945 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_360 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_359 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_944 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_943 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_942 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_941 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_940 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_939 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_938 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_937 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_936 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_935 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_358 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_357 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_356 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_355 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_354 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_353 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_352 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_351 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_350 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_349 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_348 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_347 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_346 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_345 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_344 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_343 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_342 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_341 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_934 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_933 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_932 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_931 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_930 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_929 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_928 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_927 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_926 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_925 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_924 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_923 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_922 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_921 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_920 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_919 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_918 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_917 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_916 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_915 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_914 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_913 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_912 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_911 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_910 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_909 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_908 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_907 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_906 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_905 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_904 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_44 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_43 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_903 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_902 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_901 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_42 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_41 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_11 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_990 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_989 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_988 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_987 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_986 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_985 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_984 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_983 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_982 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_981 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_980 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_979 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_978 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_977 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_976 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_975 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_974 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_973 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_972 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_971 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_970 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_969 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_968 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_967 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_966 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_965 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_964 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_374 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_373 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_963 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_372 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_962 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_371 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_370 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_961 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_369 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_960 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_368 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_367 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_959 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_366 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_958 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_957 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_956 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_955 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_954 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_953 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_952 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_951 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_950 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_949 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_365 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_948 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_947 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_946 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_364 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_363 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_362 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_361 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_945 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_360 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_359 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_944 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_943 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_942 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_941 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_940 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_939 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_938 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_937 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_936 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_935 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_358 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_357 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_356 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_355 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_354 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_353 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_352 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_351 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_350 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_349 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_348 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_347 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_346 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_345 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_344 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_343 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_342 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_341 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_934 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_933 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_932 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_931 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_930 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_929 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_928 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_927 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_926 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_925 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_924 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_923 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_922 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_921 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_920 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_919 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_918 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_917 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_916 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_915 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_914 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_913 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_912 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_911 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_910 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_909 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_908 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_907 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_906 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_905 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_904 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_44 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_43 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_903 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_902 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_901 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_42 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_41 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_900 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_899 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_898 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_897 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_896 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_895 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_894 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_893 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_892 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_891 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_890 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_889 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_888 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_887 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_886 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_885 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_884 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_883 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_882 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_881 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_880 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_879 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_878 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_877 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_876 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_875 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_874 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_340 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_339 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_873 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_338 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_872 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_337 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_336 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_871 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_335 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_870 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_334 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_333 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_869 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_332 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_868 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_867 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_866 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_865 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_864 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_863 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_862 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_861 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_860 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_859 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_331 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_858 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_857 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_856 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_330 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_329 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_328 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_327 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_855 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_326 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_325 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_854 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_853 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_852 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_851 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_850 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_849 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_848 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_847 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_846 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_845 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_324 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_323 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_322 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_321 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_320 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_319 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_318 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_317 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_316 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_315 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_314 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_313 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_312 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_311 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_310 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_309 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_308 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_307 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_844 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_843 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_842 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_841 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_840 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_839 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_838 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_837 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_836 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_835 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_834 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_833 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_832 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_831 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_830 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_829 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_828 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_827 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_826 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_825 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_824 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_823 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_822 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_821 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_820 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_819 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_818 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_817 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_816 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_815 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_814 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_40 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_39 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_813 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_812 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_811 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_38 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_37 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_10 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_900 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_899 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_898 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_897 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_896 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_895 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_894 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_893 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_892 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_891 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_890 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_889 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_888 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_887 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_886 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_885 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_884 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_883 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_882 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_881 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_880 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_879 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_878 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_877 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_876 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_875 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_874 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_340 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_339 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_873 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_338 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_872 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_337 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_336 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_871 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_335 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_870 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_334 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_333 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_869 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_332 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_868 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_867 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_866 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_865 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_864 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_863 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_862 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_861 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_860 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_859 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_331 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_858 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_857 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_856 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_330 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_329 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_328 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_327 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_855 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_326 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_325 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_854 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_853 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_852 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_851 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_850 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_849 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_848 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_847 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_846 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_845 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_324 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_323 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_322 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_321 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_320 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_319 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_318 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_317 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_316 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_315 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_314 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_313 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_312 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_311 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_310 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_309 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_308 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_307 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_844 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_843 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_842 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_841 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_840 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_839 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_838 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_837 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_836 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_835 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_834 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_833 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_832 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_831 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_830 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_829 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_828 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_827 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_826 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_825 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_824 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_823 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_822 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_821 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_820 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_819 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_818 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_817 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_816 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_815 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_814 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_40 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_39 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_813 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_812 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_811 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_38 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_37 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_810 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_809 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_808 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_807 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_806 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_805 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_804 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_803 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_802 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_801 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_800 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_799 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_798 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_797 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_796 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_795 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_794 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_793 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_792 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_791 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_790 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_789 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_788 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_787 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_786 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_785 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_784 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_306 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_305 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_783 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_304 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_782 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_303 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_302 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_781 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_301 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_780 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_300 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_299 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_779 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_298 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_778 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_777 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_776 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_775 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_774 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_773 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_772 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_771 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_770 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_769 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_297 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_768 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_767 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_766 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_296 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_295 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_294 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_293 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_765 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_292 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_291 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_764 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_763 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_762 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_761 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_760 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_759 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_758 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_757 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_756 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_755 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_290 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_289 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_288 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_287 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_286 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_285 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_284 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_283 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_282 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_281 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_280 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_279 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_278 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_277 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_276 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_275 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_274 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_273 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_754 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_753 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_752 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_751 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_750 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_749 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_748 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_747 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_746 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_745 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_744 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_743 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_742 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_741 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_740 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_739 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_738 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_737 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_736 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_735 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_734 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_733 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_732 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_731 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_730 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_729 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_728 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_727 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_726 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_725 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_724 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_36 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_35 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_723 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_722 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_721 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_34 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_33 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_9 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_810 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_809 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_808 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_807 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_806 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_805 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_804 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_803 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_802 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_801 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_800 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_799 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_798 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_797 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_796 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_795 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_794 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_793 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_792 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_791 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_790 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_789 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_788 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_787 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_786 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_785 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_784 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_306 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_305 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_783 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_304 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_782 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_303 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_302 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_781 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_301 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_780 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_300 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_299 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_779 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_298 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_778 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_777 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_776 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_775 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_774 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_773 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_772 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_771 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_770 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_769 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_297 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_768 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_767 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_766 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_296 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_295 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_294 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_293 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_765 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_292 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_291 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_764 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_763 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_762 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_761 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_760 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_759 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_758 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_757 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_756 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_755 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_290 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_289 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_288 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_287 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_286 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_285 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_284 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_283 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_282 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_281 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_280 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_279 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_278 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_277 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_276 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_275 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_274 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_273 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_754 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_753 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_752 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_751 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_750 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_749 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_748 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_747 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_746 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_745 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_744 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_743 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_742 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_741 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_740 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_739 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_738 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_737 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_736 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_735 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_734 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_733 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_732 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_731 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_730 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_729 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_728 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_727 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_726 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_725 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_724 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_36 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_35 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_723 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_722 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_721 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_34 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_33 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_720 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_719 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_718 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_717 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_716 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_715 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_714 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_713 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_712 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_711 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_710 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_709 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_708 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_707 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_706 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_705 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_704 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_703 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_702 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_701 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_700 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_699 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_698 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_697 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_696 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_695 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_694 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_272 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_271 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_693 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_270 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_692 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_269 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_268 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_691 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_267 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_690 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_266 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_265 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_689 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_264 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_688 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_687 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_686 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_685 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_684 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_683 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_682 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_681 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_680 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_679 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_263 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_678 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_677 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_676 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_262 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_261 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_260 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_259 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_675 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_258 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_257 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_674 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_673 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_672 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_671 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_670 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_669 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_668 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_667 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_666 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_665 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_256 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_255 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_254 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_253 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_252 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_251 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_250 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_249 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_248 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_247 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_246 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_245 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_244 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_243 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_242 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_241 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_240 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_239 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_664 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_663 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_662 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_661 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_660 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_659 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_658 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_657 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_656 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_655 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_654 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_653 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_652 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_651 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_650 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_649 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_648 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_647 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_646 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_645 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_644 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_643 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_642 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_641 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_640 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_639 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_638 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_637 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_636 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_635 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_634 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_32 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_31 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_633 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_632 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_631 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_30 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_29 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_8 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_720 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_719 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_718 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_717 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_716 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_715 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_714 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_713 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_712 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_711 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_710 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_709 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_708 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_707 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_706 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_705 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_704 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_703 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_702 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_701 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_700 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_699 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_698 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_697 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_696 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_695 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_694 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_272 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_271 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_693 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_270 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_692 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_269 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_268 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_691 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_267 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_690 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_266 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_265 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_689 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_264 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_688 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_687 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_686 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_685 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_684 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_683 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_682 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_681 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_680 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_679 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_263 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_678 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_677 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_676 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_262 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_261 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_260 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_259 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_675 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_258 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_257 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_674 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_673 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_672 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_671 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_670 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_669 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_668 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_667 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_666 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_665 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_256 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_255 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_254 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_253 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_252 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_251 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_250 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_249 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_248 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_247 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_246 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_245 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_244 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_243 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_242 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_241 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_240 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_239 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_664 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_663 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_662 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_661 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_660 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_659 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_658 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_657 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_656 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_655 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_654 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_653 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_652 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_651 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_650 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_649 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_648 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_647 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_646 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_645 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_644 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_643 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_642 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_641 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_640 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_639 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_638 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_637 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_636 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_635 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_634 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_32 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_31 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_633 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_632 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_631 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_30 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_29 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_630 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_629 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_628 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_627 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_626 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_625 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_624 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_623 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_622 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_621 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_620 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_619 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_618 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_617 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_616 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_615 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_614 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_613 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_612 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_611 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_610 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_609 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_608 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_607 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_606 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_605 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_604 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_238 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_237 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_603 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_236 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_602 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_235 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_234 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_601 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_233 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_600 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_232 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_231 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_599 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_230 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_598 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_597 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_596 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_595 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_594 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_593 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_592 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_591 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_590 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_589 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_229 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_588 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_587 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_586 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_228 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_227 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_226 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_225 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_585 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_224 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_223 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_584 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_583 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_582 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_581 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_580 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_579 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_578 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_577 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_576 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_575 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_222 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_221 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_220 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_219 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_218 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_217 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_216 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_215 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_214 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_213 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_212 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_211 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_210 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_209 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_208 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_207 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_206 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_205 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_574 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_573 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_572 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_571 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_570 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_569 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_568 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_567 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_566 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_565 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_564 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_563 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_562 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_561 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_560 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_559 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_558 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_557 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_556 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_555 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_554 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_553 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_552 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_551 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_550 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_549 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_548 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_547 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_546 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_545 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_544 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_28 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_27 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_543 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_542 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_541 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_26 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_25 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_7 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_630 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_629 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_628 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_627 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_626 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_625 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_624 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_623 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_622 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_621 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_620 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_619 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_618 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_617 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_616 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_615 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_614 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_613 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_612 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_611 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_610 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_609 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_608 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_607 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_606 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_605 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_604 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_238 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_237 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_603 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_236 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_602 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_235 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_234 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_601 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_233 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_600 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_232 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_231 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_599 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_230 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_598 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_597 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_596 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_595 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_594 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_593 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_592 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_591 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_590 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_589 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_229 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_588 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_587 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_586 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_228 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_227 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_226 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_225 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_585 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_224 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_223 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_584 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_583 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_582 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_581 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_580 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_579 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_578 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_577 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_576 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_575 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_222 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_221 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_220 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_219 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_218 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_217 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_216 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_215 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_214 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_213 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_212 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_211 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_210 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_209 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_208 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_207 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_206 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_205 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_574 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_573 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_572 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_571 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_570 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_569 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_568 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_567 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_566 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_565 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_564 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_563 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_562 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_561 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_560 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_559 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_558 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_557 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_556 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_555 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_554 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_553 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_552 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_551 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_550 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_549 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_548 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_547 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_546 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_545 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_544 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_28 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_27 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_543 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_542 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_541 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_26 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_25 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_540 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_539 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_538 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_537 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_536 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_535 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_534 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_533 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_532 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_531 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_530 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_529 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_528 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_527 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_526 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_525 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_524 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_523 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_522 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_521 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_520 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_519 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_518 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_517 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_516 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_515 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_514 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_204 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_203 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_513 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_202 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_512 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_201 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_200 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_511 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_199 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_510 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_198 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_197 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_509 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_196 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_508 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_507 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_506 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_505 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_504 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_503 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_502 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_501 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_500 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_499 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_195 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_498 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_497 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_496 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_194 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_193 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_192 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_191 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_495 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_190 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_189 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_494 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_493 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_492 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_491 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_490 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_489 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_488 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_487 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_486 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_485 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_188 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_187 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_186 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_185 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_184 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_183 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_182 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_181 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_180 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_179 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_178 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_177 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_176 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_175 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_174 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_173 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_172 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_171 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_484 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_483 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_482 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_481 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_480 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_479 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_478 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_477 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_476 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_475 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_474 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_473 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_472 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_471 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_470 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_469 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_468 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_467 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_466 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_465 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_464 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_463 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_462 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_461 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_460 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_459 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_458 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_457 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_456 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_455 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_454 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_24 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_23 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_453 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_452 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_451 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_22 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_21 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_6 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_540 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_539 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_538 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_537 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_536 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_535 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_534 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_533 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_532 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_531 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_530 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_529 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_528 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_527 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_526 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_525 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_524 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_523 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_522 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_521 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_520 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_519 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_518 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_517 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_516 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_515 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_514 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_204 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_203 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_513 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_202 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_512 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_201 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_200 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_511 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_199 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_510 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_198 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_197 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_509 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_196 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_508 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_507 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_506 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_505 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_504 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_503 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_502 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_501 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_500 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_499 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_195 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_498 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_497 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_496 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_194 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_193 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_192 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_191 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_495 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_190 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_189 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_494 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_493 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_492 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_491 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_490 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_489 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_488 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_487 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_486 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_485 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_188 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_187 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_186 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_185 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_184 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_183 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_182 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_181 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_180 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_179 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_178 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_177 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_176 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_175 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_174 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_173 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_172 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_171 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_484 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_483 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_482 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_481 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_480 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_479 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_478 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_477 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_476 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_475 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_474 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_473 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_472 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_471 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_470 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_469 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_468 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_467 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_466 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_465 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_464 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_463 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_462 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_461 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_460 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_459 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_458 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_457 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_456 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_455 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_454 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_24 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_23 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_453 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_452 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_451 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_22 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_21 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_450 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_449 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_448 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_447 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_446 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_445 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_444 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_443 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_442 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_441 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_440 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_439 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_438 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_437 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_436 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_435 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_434 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_433 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_432 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_431 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_430 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_429 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_428 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_427 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_426 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_425 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_424 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_170 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_169 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_423 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_168 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_422 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_167 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_166 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_421 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_165 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_420 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_164 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_163 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_419 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_162 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_418 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_417 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_416 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_415 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_414 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_413 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_412 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_411 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_410 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_409 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_161 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_408 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_407 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_406 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_160 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_159 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_158 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_157 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_405 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_156 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_155 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_404 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_403 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_402 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_401 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_400 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_399 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_398 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_397 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_396 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_395 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_154 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_153 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_152 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_151 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_150 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_149 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_148 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_147 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_146 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_145 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_144 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_143 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_142 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_141 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_140 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_139 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_138 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_137 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_394 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_393 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_392 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_391 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_390 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_389 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_388 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_387 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_386 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_385 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_384 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_383 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_382 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_381 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_380 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_379 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_378 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_377 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_376 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_375 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_374 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_373 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_372 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_371 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_370 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_369 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_368 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_367 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_366 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_365 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_364 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_20 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_19 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_363 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_362 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_361 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_18 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_17 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_5 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_450 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_449 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_448 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_447 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_446 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_445 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_444 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_443 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_442 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_441 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_440 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_439 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_438 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_437 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_436 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_435 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_434 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_433 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_432 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_431 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_430 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_429 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_428 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_427 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_426 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_425 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_424 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_170 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_169 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_423 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_168 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_422 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_167 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_166 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_421 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_165 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_420 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_164 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_163 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_419 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_162 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_418 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_417 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_416 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_415 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_414 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_413 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_412 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_411 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_410 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_409 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_161 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_408 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_407 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_406 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_160 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_159 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_158 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_157 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_405 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_156 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_155 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_404 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_403 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_402 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_401 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_400 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_399 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_398 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_397 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_396 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_395 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_154 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_153 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_152 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_151 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_150 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_149 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_148 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_147 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_146 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_145 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_144 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_143 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_142 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_141 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_140 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_139 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_138 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_137 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_394 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_393 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_392 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_391 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_390 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_389 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_388 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_387 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_386 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_385 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_384 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_383 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_382 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_381 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_380 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_379 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_378 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_377 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_376 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_375 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_374 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_373 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_372 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_371 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_370 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_369 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_368 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_367 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_366 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_365 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_364 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_20 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_19 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_363 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_362 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_361 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_18 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_17 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module SubBytes ( input0, output0 );
  input [127:0] input0;
  output [127:0] output0;


  Sbox_0 Inst_Sbox_0 ( .x(input0[7:0]), .y(output0[7:0]) );
  Sbox_19 Inst_Sbox_1 ( .x(input0[15:8]), .y(output0[15:8]) );
  Sbox_18 Inst_Sbox_2 ( .x(input0[23:16]), .y(output0[23:16]) );
  Sbox_17 Inst_Sbox_3 ( .x(input0[31:24]), .y(output0[31:24]) );
  Sbox_16 Inst_Sbox_4 ( .x(input0[39:32]), .y(output0[39:32]) );
  Sbox_15 Inst_Sbox_5 ( .x(input0[47:40]), .y(output0[47:40]) );
  Sbox_14 Inst_Sbox_6 ( .x(input0[55:48]), .y(output0[55:48]) );
  Sbox_13 Inst_Sbox_7 ( .x(input0[63:56]), .y(output0[63:56]) );
  Sbox_12 Inst_Sbox_8 ( .x(input0[71:64]), .y(output0[71:64]) );
  Sbox_11 Inst_Sbox_9 ( .x(input0[79:72]), .y(output0[79:72]) );
  Sbox_10 Inst_Sbox_10 ( .x(input0[87:80]), .y(output0[87:80]) );
  Sbox_9 Inst_Sbox_11 ( .x(input0[95:88]), .y(output0[95:88]) );
  Sbox_8 Inst_Sbox_12 ( .x(input0[103:96]), .y(output0[103:96]) );
  Sbox_7 Inst_Sbox_13 ( .x(input0[111:104]), .y(output0[111:104]) );
  Sbox_6 Inst_Sbox_14 ( .x(input0[119:112]), .y(output0[119:112]) );
  Sbox_5 Inst_Sbox_15 ( .x(input0[127:120]), .y(output0[127:120]) );
endmodule


module ShiftRows ( input0, output0 );
  input [127:0] input0;
  output [127:0] output0;

  assign output0[127] = input0[127];
  assign output0[126] = input0[126];
  assign output0[125] = input0[125];
  assign output0[124] = input0[124];
  assign output0[123] = input0[123];
  assign output0[122] = input0[122];
  assign output0[121] = input0[121];
  assign output0[120] = input0[120];
  assign output0[119] = input0[87];
  assign output0[118] = input0[86];
  assign output0[117] = input0[85];
  assign output0[116] = input0[84];
  assign output0[115] = input0[83];
  assign output0[114] = input0[82];
  assign output0[113] = input0[81];
  assign output0[112] = input0[80];
  assign output0[111] = input0[47];
  assign output0[110] = input0[46];
  assign output0[109] = input0[45];
  assign output0[108] = input0[44];
  assign output0[107] = input0[43];
  assign output0[106] = input0[42];
  assign output0[105] = input0[41];
  assign output0[104] = input0[40];
  assign output0[103] = input0[7];
  assign output0[102] = input0[6];
  assign output0[101] = input0[5];
  assign output0[100] = input0[4];
  assign output0[99] = input0[3];
  assign output0[98] = input0[2];
  assign output0[97] = input0[1];
  assign output0[96] = input0[0];
  assign output0[95] = input0[95];
  assign output0[94] = input0[94];
  assign output0[93] = input0[93];
  assign output0[92] = input0[92];
  assign output0[91] = input0[91];
  assign output0[90] = input0[90];
  assign output0[89] = input0[89];
  assign output0[88] = input0[88];
  assign output0[87] = input0[55];
  assign output0[86] = input0[54];
  assign output0[85] = input0[53];
  assign output0[84] = input0[52];
  assign output0[83] = input0[51];
  assign output0[82] = input0[50];
  assign output0[81] = input0[49];
  assign output0[80] = input0[48];
  assign output0[79] = input0[15];
  assign output0[78] = input0[14];
  assign output0[77] = input0[13];
  assign output0[76] = input0[12];
  assign output0[75] = input0[11];
  assign output0[74] = input0[10];
  assign output0[73] = input0[9];
  assign output0[72] = input0[8];
  assign output0[71] = input0[103];
  assign output0[70] = input0[102];
  assign output0[69] = input0[101];
  assign output0[68] = input0[100];
  assign output0[67] = input0[99];
  assign output0[66] = input0[98];
  assign output0[65] = input0[97];
  assign output0[64] = input0[96];
  assign output0[63] = input0[63];
  assign output0[62] = input0[62];
  assign output0[61] = input0[61];
  assign output0[60] = input0[60];
  assign output0[59] = input0[59];
  assign output0[58] = input0[58];
  assign output0[57] = input0[57];
  assign output0[56] = input0[56];
  assign output0[55] = input0[23];
  assign output0[54] = input0[22];
  assign output0[53] = input0[21];
  assign output0[52] = input0[20];
  assign output0[51] = input0[19];
  assign output0[50] = input0[18];
  assign output0[49] = input0[17];
  assign output0[48] = input0[16];
  assign output0[47] = input0[111];
  assign output0[46] = input0[110];
  assign output0[45] = input0[109];
  assign output0[44] = input0[108];
  assign output0[43] = input0[107];
  assign output0[42] = input0[106];
  assign output0[41] = input0[105];
  assign output0[40] = input0[104];
  assign output0[39] = input0[71];
  assign output0[38] = input0[70];
  assign output0[37] = input0[69];
  assign output0[36] = input0[68];
  assign output0[35] = input0[67];
  assign output0[34] = input0[66];
  assign output0[33] = input0[65];
  assign output0[32] = input0[64];
  assign output0[31] = input0[31];
  assign output0[30] = input0[30];
  assign output0[29] = input0[29];
  assign output0[28] = input0[28];
  assign output0[27] = input0[27];
  assign output0[26] = input0[26];
  assign output0[25] = input0[25];
  assign output0[24] = input0[24];
  assign output0[23] = input0[119];
  assign output0[22] = input0[118];
  assign output0[21] = input0[117];
  assign output0[20] = input0[116];
  assign output0[19] = input0[115];
  assign output0[18] = input0[114];
  assign output0[17] = input0[113];
  assign output0[16] = input0[112];
  assign output0[15] = input0[79];
  assign output0[14] = input0[78];
  assign output0[13] = input0[77];
  assign output0[12] = input0[76];
  assign output0[11] = input0[75];
  assign output0[10] = input0[74];
  assign output0[9] = input0[73];
  assign output0[8] = input0[72];
  assign output0[7] = input0[39];
  assign output0[6] = input0[38];
  assign output0[5] = input0[37];
  assign output0[4] = input0[36];
  assign output0[3] = input0[35];
  assign output0[2] = input0[34];
  assign output0[1] = input0[33];
  assign output0[0] = input0[32];

endmodule


module Mul2_0 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_15 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_14 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_13 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module MixOneColumn_0 ( input0, output0 );
  input [31:0] input0;
  output [31:0] output0;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  wire   [31:0] DoubleBytes;

  Mul2_0 Mul2Inst_0 ( .input0(input0[31:24]), .output0(DoubleBytes[31:24]) );
  Mul2_15 Mul2Inst_1 ( .input0(input0[23:16]), .output0(DoubleBytes[23:16]) );
  Mul2_14 Mul2Inst_2 ( .input0(input0[15:8]), .output0(DoubleBytes[15:8]) );
  Mul2_13 Mul2Inst_3 ( .input0(input0[7:0]), .output0(DoubleBytes[7:0]) );
  XOR2_X1 U1 ( .A(DoubleBytes[0]), .B(input0[24]), .Z(n59) );
  XOR2_X1 U2 ( .A(input0[16]), .B(DoubleBytes[24]), .Z(n23) );
  XNOR2_X1 U3 ( .A(n59), .B(n23), .ZN(n1) );
  XNOR2_X1 U4 ( .A(n1), .B(input0[8]), .ZN(output0[0]) );
  XOR2_X1 U5 ( .A(DoubleBytes[2]), .B(input0[26]), .Z(n37) );
  XNOR2_X1 U6 ( .A(n37), .B(input0[18]), .ZN(n2) );
  XOR2_X1 U7 ( .A(input0[2]), .B(DoubleBytes[10]), .Z(n10) );
  XNOR2_X1 U8 ( .A(n2), .B(n10), .ZN(output0[10]) );
  XOR2_X1 U9 ( .A(DoubleBytes[3]), .B(input0[27]), .Z(n44) );
  XNOR2_X1 U10 ( .A(n44), .B(input0[19]), .ZN(n3) );
  XOR2_X1 U11 ( .A(input0[3]), .B(DoubleBytes[11]), .Z(n12) );
  XNOR2_X1 U12 ( .A(n3), .B(n12), .ZN(output0[11]) );
  XOR2_X1 U13 ( .A(DoubleBytes[4]), .B(input0[28]), .Z(n47) );
  XNOR2_X1 U14 ( .A(n47), .B(input0[20]), .ZN(n4) );
  XOR2_X1 U15 ( .A(input0[4]), .B(DoubleBytes[12]), .Z(n15) );
  XNOR2_X1 U16 ( .A(n4), .B(n15), .ZN(output0[12]) );
  XOR2_X1 U17 ( .A(DoubleBytes[5]), .B(input0[29]), .Z(n50) );
  XNOR2_X1 U18 ( .A(n50), .B(input0[21]), .ZN(n5) );
  XOR2_X1 U19 ( .A(input0[5]), .B(DoubleBytes[13]), .Z(n17) );
  XNOR2_X1 U20 ( .A(n5), .B(n17), .ZN(output0[13]) );
  XOR2_X1 U21 ( .A(DoubleBytes[6]), .B(input0[30]), .Z(n53) );
  XNOR2_X1 U22 ( .A(n53), .B(input0[22]), .ZN(n6) );
  XOR2_X1 U23 ( .A(input0[6]), .B(DoubleBytes[14]), .Z(n19) );
  XNOR2_X1 U24 ( .A(n6), .B(n19), .ZN(output0[14]) );
  XOR2_X1 U25 ( .A(DoubleBytes[7]), .B(input0[31]), .Z(n56) );
  XNOR2_X1 U26 ( .A(n56), .B(input0[23]), .ZN(n7) );
  XOR2_X1 U27 ( .A(input0[7]), .B(DoubleBytes[15]), .Z(n21) );
  XNOR2_X1 U28 ( .A(n7), .B(n21), .ZN(output0[15]) );
  XOR2_X1 U29 ( .A(DoubleBytes[8]), .B(input0[0]), .Z(n60) );
  XNOR2_X1 U30 ( .A(input0[24]), .B(n60), .ZN(n8) );
  XOR2_X1 U31 ( .A(input0[8]), .B(DoubleBytes[16]), .Z(n24) );
  XNOR2_X1 U32 ( .A(n8), .B(n24), .ZN(output0[16]) );
  XOR2_X1 U33 ( .A(DoubleBytes[9]), .B(input0[1]), .Z(n63) );
  XNOR2_X1 U34 ( .A(n63), .B(input0[25]), .ZN(n9) );
  XOR2_X1 U35 ( .A(DoubleBytes[17]), .B(input0[9]), .Z(n26) );
  XNOR2_X1 U36 ( .A(n9), .B(n26), .ZN(output0[17]) );
  XNOR2_X1 U37 ( .A(input0[26]), .B(n10), .ZN(n11) );
  XOR2_X1 U38 ( .A(input0[10]), .B(DoubleBytes[18]), .Z(n29) );
  XNOR2_X1 U39 ( .A(n11), .B(n29), .ZN(output0[18]) );
  XNOR2_X1 U40 ( .A(input0[27]), .B(n12), .ZN(n13) );
  XOR2_X1 U41 ( .A(input0[11]), .B(DoubleBytes[19]), .Z(n31) );
  XNOR2_X1 U42 ( .A(n13), .B(n31), .ZN(output0[19]) );
  XOR2_X1 U43 ( .A(input0[25]), .B(DoubleBytes[1]), .Z(n62) );
  XNOR2_X1 U44 ( .A(input0[9]), .B(n62), .ZN(n14) );
  XOR2_X1 U45 ( .A(input0[17]), .B(DoubleBytes[25]), .Z(n27) );
  XNOR2_X1 U46 ( .A(n14), .B(n27), .ZN(output0[1]) );
  XNOR2_X1 U47 ( .A(input0[28]), .B(n15), .ZN(n16) );
  XOR2_X1 U48 ( .A(input0[12]), .B(DoubleBytes[20]), .Z(n33) );
  XNOR2_X1 U49 ( .A(n16), .B(n33), .ZN(output0[20]) );
  XNOR2_X1 U50 ( .A(input0[29]), .B(n17), .ZN(n18) );
  XOR2_X1 U51 ( .A(input0[13]), .B(DoubleBytes[21]), .Z(n35) );
  XNOR2_X1 U52 ( .A(n18), .B(n35), .ZN(output0[21]) );
  XNOR2_X1 U53 ( .A(input0[30]), .B(n19), .ZN(n20) );
  XOR2_X1 U54 ( .A(input0[14]), .B(DoubleBytes[22]), .Z(n40) );
  XNOR2_X1 U55 ( .A(n20), .B(n40), .ZN(output0[22]) );
  XNOR2_X1 U56 ( .A(input0[31]), .B(n21), .ZN(n22) );
  XOR2_X1 U57 ( .A(input0[15]), .B(DoubleBytes[23]), .Z(n42) );
  XNOR2_X1 U58 ( .A(n22), .B(n42), .ZN(output0[23]) );
  XNOR2_X1 U59 ( .A(n23), .B(input0[0]), .ZN(n25) );
  XNOR2_X1 U60 ( .A(n25), .B(n24), .ZN(output0[24]) );
  XNOR2_X1 U61 ( .A(input0[1]), .B(n26), .ZN(n28) );
  XNOR2_X1 U62 ( .A(n28), .B(n27), .ZN(output0[25]) );
  XNOR2_X1 U63 ( .A(input0[2]), .B(n29), .ZN(n30) );
  XOR2_X1 U64 ( .A(input0[18]), .B(DoubleBytes[26]), .Z(n38) );
  XNOR2_X1 U65 ( .A(n30), .B(n38), .ZN(output0[26]) );
  XNOR2_X1 U66 ( .A(input0[3]), .B(n31), .ZN(n32) );
  XOR2_X1 U67 ( .A(input0[19]), .B(DoubleBytes[27]), .Z(n45) );
  XNOR2_X1 U68 ( .A(n32), .B(n45), .ZN(output0[27]) );
  XNOR2_X1 U69 ( .A(input0[4]), .B(n33), .ZN(n34) );
  XOR2_X1 U70 ( .A(input0[20]), .B(DoubleBytes[28]), .Z(n48) );
  XNOR2_X1 U71 ( .A(n34), .B(n48), .ZN(output0[28]) );
  XNOR2_X1 U72 ( .A(input0[5]), .B(n35), .ZN(n36) );
  XOR2_X1 U73 ( .A(input0[21]), .B(DoubleBytes[29]), .Z(n51) );
  XNOR2_X1 U74 ( .A(n36), .B(n51), .ZN(output0[29]) );
  XNOR2_X1 U75 ( .A(n37), .B(input0[10]), .ZN(n39) );
  XNOR2_X1 U76 ( .A(n39), .B(n38), .ZN(output0[2]) );
  XNOR2_X1 U77 ( .A(input0[6]), .B(n40), .ZN(n41) );
  XOR2_X1 U78 ( .A(input0[22]), .B(DoubleBytes[30]), .Z(n54) );
  XNOR2_X1 U79 ( .A(n41), .B(n54), .ZN(output0[30]) );
  XNOR2_X1 U80 ( .A(input0[7]), .B(n42), .ZN(n43) );
  XOR2_X1 U81 ( .A(input0[23]), .B(DoubleBytes[31]), .Z(n57) );
  XNOR2_X1 U82 ( .A(n43), .B(n57), .ZN(output0[31]) );
  XNOR2_X1 U83 ( .A(n44), .B(input0[11]), .ZN(n46) );
  XNOR2_X1 U84 ( .A(n46), .B(n45), .ZN(output0[3]) );
  XNOR2_X1 U85 ( .A(n47), .B(input0[12]), .ZN(n49) );
  XNOR2_X1 U86 ( .A(n49), .B(n48), .ZN(output0[4]) );
  XNOR2_X1 U87 ( .A(n50), .B(input0[13]), .ZN(n52) );
  XNOR2_X1 U88 ( .A(n52), .B(n51), .ZN(output0[5]) );
  XNOR2_X1 U89 ( .A(n53), .B(input0[14]), .ZN(n55) );
  XNOR2_X1 U90 ( .A(n55), .B(n54), .ZN(output0[6]) );
  XNOR2_X1 U91 ( .A(n56), .B(input0[15]), .ZN(n58) );
  XNOR2_X1 U92 ( .A(n58), .B(n57), .ZN(output0[7]) );
  XNOR2_X1 U93 ( .A(n59), .B(input0[16]), .ZN(n61) );
  XNOR2_X1 U94 ( .A(n61), .B(n60), .ZN(output0[8]) );
  XNOR2_X1 U95 ( .A(n63), .B(n62), .ZN(n64) );
  XNOR2_X1 U96 ( .A(n64), .B(input0[17]), .ZN(output0[9]) );
endmodule


module Mul2_12 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_11 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_10 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_9 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module MixOneColumn_3 ( input0, output0 );
  input [31:0] input0;
  output [31:0] output0;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  wire   [31:0] DoubleBytes;

  Mul2_12 Mul2Inst_0 ( .input0(input0[31:24]), .output0(DoubleBytes[31:24]) );
  Mul2_11 Mul2Inst_1 ( .input0(input0[23:16]), .output0(DoubleBytes[23:16]) );
  Mul2_10 Mul2Inst_2 ( .input0(input0[15:8]), .output0(DoubleBytes[15:8]) );
  Mul2_9 Mul2Inst_3 ( .input0(input0[7:0]), .output0(DoubleBytes[7:0]) );
  XOR2_X1 U1 ( .A(DoubleBytes[0]), .B(input0[24]), .Z(n59) );
  XOR2_X1 U2 ( .A(input0[16]), .B(DoubleBytes[24]), .Z(n23) );
  XNOR2_X1 U3 ( .A(n59), .B(n23), .ZN(n1) );
  XNOR2_X1 U4 ( .A(n1), .B(input0[8]), .ZN(output0[0]) );
  XOR2_X1 U5 ( .A(DoubleBytes[2]), .B(input0[26]), .Z(n37) );
  XNOR2_X1 U6 ( .A(n37), .B(input0[18]), .ZN(n2) );
  XOR2_X1 U7 ( .A(input0[2]), .B(DoubleBytes[10]), .Z(n10) );
  XNOR2_X1 U8 ( .A(n2), .B(n10), .ZN(output0[10]) );
  XOR2_X1 U9 ( .A(DoubleBytes[3]), .B(input0[27]), .Z(n44) );
  XNOR2_X1 U10 ( .A(n44), .B(input0[19]), .ZN(n3) );
  XOR2_X1 U11 ( .A(input0[3]), .B(DoubleBytes[11]), .Z(n12) );
  XNOR2_X1 U12 ( .A(n3), .B(n12), .ZN(output0[11]) );
  XOR2_X1 U13 ( .A(DoubleBytes[4]), .B(input0[28]), .Z(n47) );
  XNOR2_X1 U14 ( .A(n47), .B(input0[20]), .ZN(n4) );
  XOR2_X1 U15 ( .A(input0[4]), .B(DoubleBytes[12]), .Z(n15) );
  XNOR2_X1 U16 ( .A(n4), .B(n15), .ZN(output0[12]) );
  XOR2_X1 U17 ( .A(DoubleBytes[5]), .B(input0[29]), .Z(n50) );
  XNOR2_X1 U18 ( .A(n50), .B(input0[21]), .ZN(n5) );
  XOR2_X1 U19 ( .A(input0[5]), .B(DoubleBytes[13]), .Z(n17) );
  XNOR2_X1 U20 ( .A(n5), .B(n17), .ZN(output0[13]) );
  XOR2_X1 U21 ( .A(DoubleBytes[6]), .B(input0[30]), .Z(n53) );
  XNOR2_X1 U22 ( .A(n53), .B(input0[22]), .ZN(n6) );
  XOR2_X1 U23 ( .A(input0[6]), .B(DoubleBytes[14]), .Z(n19) );
  XNOR2_X1 U24 ( .A(n6), .B(n19), .ZN(output0[14]) );
  XOR2_X1 U25 ( .A(DoubleBytes[7]), .B(input0[31]), .Z(n56) );
  XNOR2_X1 U26 ( .A(n56), .B(input0[23]), .ZN(n7) );
  XOR2_X1 U27 ( .A(input0[7]), .B(DoubleBytes[15]), .Z(n21) );
  XNOR2_X1 U28 ( .A(n7), .B(n21), .ZN(output0[15]) );
  XOR2_X1 U29 ( .A(DoubleBytes[8]), .B(input0[0]), .Z(n60) );
  XNOR2_X1 U30 ( .A(input0[24]), .B(n60), .ZN(n8) );
  XOR2_X1 U31 ( .A(input0[8]), .B(DoubleBytes[16]), .Z(n24) );
  XNOR2_X1 U32 ( .A(n8), .B(n24), .ZN(output0[16]) );
  XOR2_X1 U33 ( .A(DoubleBytes[9]), .B(input0[1]), .Z(n63) );
  XNOR2_X1 U34 ( .A(n63), .B(input0[25]), .ZN(n9) );
  XOR2_X1 U35 ( .A(DoubleBytes[17]), .B(input0[9]), .Z(n26) );
  XNOR2_X1 U36 ( .A(n9), .B(n26), .ZN(output0[17]) );
  XNOR2_X1 U37 ( .A(input0[26]), .B(n10), .ZN(n11) );
  XOR2_X1 U38 ( .A(input0[10]), .B(DoubleBytes[18]), .Z(n29) );
  XNOR2_X1 U39 ( .A(n11), .B(n29), .ZN(output0[18]) );
  XNOR2_X1 U40 ( .A(input0[27]), .B(n12), .ZN(n13) );
  XOR2_X1 U41 ( .A(input0[11]), .B(DoubleBytes[19]), .Z(n31) );
  XNOR2_X1 U42 ( .A(n13), .B(n31), .ZN(output0[19]) );
  XOR2_X1 U43 ( .A(input0[25]), .B(DoubleBytes[1]), .Z(n62) );
  XNOR2_X1 U44 ( .A(input0[9]), .B(n62), .ZN(n14) );
  XOR2_X1 U45 ( .A(input0[17]), .B(DoubleBytes[25]), .Z(n27) );
  XNOR2_X1 U46 ( .A(n14), .B(n27), .ZN(output0[1]) );
  XNOR2_X1 U47 ( .A(input0[28]), .B(n15), .ZN(n16) );
  XOR2_X1 U48 ( .A(input0[12]), .B(DoubleBytes[20]), .Z(n33) );
  XNOR2_X1 U49 ( .A(n16), .B(n33), .ZN(output0[20]) );
  XNOR2_X1 U50 ( .A(input0[29]), .B(n17), .ZN(n18) );
  XOR2_X1 U51 ( .A(input0[13]), .B(DoubleBytes[21]), .Z(n35) );
  XNOR2_X1 U52 ( .A(n18), .B(n35), .ZN(output0[21]) );
  XNOR2_X1 U53 ( .A(input0[30]), .B(n19), .ZN(n20) );
  XOR2_X1 U54 ( .A(input0[14]), .B(DoubleBytes[22]), .Z(n40) );
  XNOR2_X1 U55 ( .A(n20), .B(n40), .ZN(output0[22]) );
  XNOR2_X1 U56 ( .A(input0[31]), .B(n21), .ZN(n22) );
  XOR2_X1 U57 ( .A(input0[15]), .B(DoubleBytes[23]), .Z(n42) );
  XNOR2_X1 U58 ( .A(n22), .B(n42), .ZN(output0[23]) );
  XNOR2_X1 U59 ( .A(n23), .B(input0[0]), .ZN(n25) );
  XNOR2_X1 U60 ( .A(n25), .B(n24), .ZN(output0[24]) );
  XNOR2_X1 U61 ( .A(input0[1]), .B(n26), .ZN(n28) );
  XNOR2_X1 U62 ( .A(n28), .B(n27), .ZN(output0[25]) );
  XNOR2_X1 U63 ( .A(input0[2]), .B(n29), .ZN(n30) );
  XOR2_X1 U64 ( .A(input0[18]), .B(DoubleBytes[26]), .Z(n38) );
  XNOR2_X1 U65 ( .A(n30), .B(n38), .ZN(output0[26]) );
  XNOR2_X1 U66 ( .A(input0[3]), .B(n31), .ZN(n32) );
  XOR2_X1 U67 ( .A(input0[19]), .B(DoubleBytes[27]), .Z(n45) );
  XNOR2_X1 U68 ( .A(n32), .B(n45), .ZN(output0[27]) );
  XNOR2_X1 U69 ( .A(input0[4]), .B(n33), .ZN(n34) );
  XOR2_X1 U70 ( .A(input0[20]), .B(DoubleBytes[28]), .Z(n48) );
  XNOR2_X1 U71 ( .A(n34), .B(n48), .ZN(output0[28]) );
  XNOR2_X1 U72 ( .A(input0[5]), .B(n35), .ZN(n36) );
  XOR2_X1 U73 ( .A(input0[21]), .B(DoubleBytes[29]), .Z(n51) );
  XNOR2_X1 U74 ( .A(n36), .B(n51), .ZN(output0[29]) );
  XNOR2_X1 U75 ( .A(n37), .B(input0[10]), .ZN(n39) );
  XNOR2_X1 U76 ( .A(n39), .B(n38), .ZN(output0[2]) );
  XNOR2_X1 U77 ( .A(input0[6]), .B(n40), .ZN(n41) );
  XOR2_X1 U78 ( .A(input0[22]), .B(DoubleBytes[30]), .Z(n54) );
  XNOR2_X1 U79 ( .A(n41), .B(n54), .ZN(output0[30]) );
  XNOR2_X1 U80 ( .A(input0[7]), .B(n42), .ZN(n43) );
  XOR2_X1 U81 ( .A(input0[23]), .B(DoubleBytes[31]), .Z(n57) );
  XNOR2_X1 U82 ( .A(n43), .B(n57), .ZN(output0[31]) );
  XNOR2_X1 U83 ( .A(n44), .B(input0[11]), .ZN(n46) );
  XNOR2_X1 U84 ( .A(n46), .B(n45), .ZN(output0[3]) );
  XNOR2_X1 U85 ( .A(n47), .B(input0[12]), .ZN(n49) );
  XNOR2_X1 U86 ( .A(n49), .B(n48), .ZN(output0[4]) );
  XNOR2_X1 U87 ( .A(n50), .B(input0[13]), .ZN(n52) );
  XNOR2_X1 U88 ( .A(n52), .B(n51), .ZN(output0[5]) );
  XNOR2_X1 U89 ( .A(n53), .B(input0[14]), .ZN(n55) );
  XNOR2_X1 U90 ( .A(n55), .B(n54), .ZN(output0[6]) );
  XNOR2_X1 U91 ( .A(n56), .B(input0[15]), .ZN(n58) );
  XNOR2_X1 U92 ( .A(n58), .B(n57), .ZN(output0[7]) );
  XNOR2_X1 U93 ( .A(n59), .B(input0[16]), .ZN(n61) );
  XNOR2_X1 U94 ( .A(n61), .B(n60), .ZN(output0[8]) );
  XNOR2_X1 U95 ( .A(n63), .B(n62), .ZN(n64) );
  XNOR2_X1 U96 ( .A(n64), .B(input0[17]), .ZN(output0[9]) );
endmodule


module Mul2_8 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_7 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_6 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_5 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module MixOneColumn_2 ( input0, output0 );
  input [31:0] input0;
  output [31:0] output0;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  wire   [31:0] DoubleBytes;

  Mul2_8 Mul2Inst_0 ( .input0(input0[31:24]), .output0(DoubleBytes[31:24]) );
  Mul2_7 Mul2Inst_1 ( .input0(input0[23:16]), .output0(DoubleBytes[23:16]) );
  Mul2_6 Mul2Inst_2 ( .input0(input0[15:8]), .output0(DoubleBytes[15:8]) );
  Mul2_5 Mul2Inst_3 ( .input0(input0[7:0]), .output0(DoubleBytes[7:0]) );
  XOR2_X1 U1 ( .A(DoubleBytes[0]), .B(input0[24]), .Z(n59) );
  XOR2_X1 U2 ( .A(input0[16]), .B(DoubleBytes[24]), .Z(n23) );
  XNOR2_X1 U3 ( .A(n59), .B(n23), .ZN(n1) );
  XNOR2_X1 U4 ( .A(n1), .B(input0[8]), .ZN(output0[0]) );
  XOR2_X1 U5 ( .A(DoubleBytes[2]), .B(input0[26]), .Z(n37) );
  XNOR2_X1 U6 ( .A(n37), .B(input0[18]), .ZN(n2) );
  XOR2_X1 U7 ( .A(input0[2]), .B(DoubleBytes[10]), .Z(n10) );
  XNOR2_X1 U8 ( .A(n2), .B(n10), .ZN(output0[10]) );
  XOR2_X1 U9 ( .A(DoubleBytes[3]), .B(input0[27]), .Z(n44) );
  XNOR2_X1 U10 ( .A(n44), .B(input0[19]), .ZN(n3) );
  XOR2_X1 U11 ( .A(input0[3]), .B(DoubleBytes[11]), .Z(n12) );
  XNOR2_X1 U12 ( .A(n3), .B(n12), .ZN(output0[11]) );
  XOR2_X1 U13 ( .A(DoubleBytes[4]), .B(input0[28]), .Z(n47) );
  XNOR2_X1 U14 ( .A(n47), .B(input0[20]), .ZN(n4) );
  XOR2_X1 U15 ( .A(input0[4]), .B(DoubleBytes[12]), .Z(n15) );
  XNOR2_X1 U16 ( .A(n4), .B(n15), .ZN(output0[12]) );
  XOR2_X1 U17 ( .A(DoubleBytes[5]), .B(input0[29]), .Z(n50) );
  XNOR2_X1 U18 ( .A(n50), .B(input0[21]), .ZN(n5) );
  XOR2_X1 U19 ( .A(input0[5]), .B(DoubleBytes[13]), .Z(n17) );
  XNOR2_X1 U20 ( .A(n5), .B(n17), .ZN(output0[13]) );
  XOR2_X1 U21 ( .A(DoubleBytes[6]), .B(input0[30]), .Z(n53) );
  XNOR2_X1 U22 ( .A(n53), .B(input0[22]), .ZN(n6) );
  XOR2_X1 U23 ( .A(input0[6]), .B(DoubleBytes[14]), .Z(n19) );
  XNOR2_X1 U24 ( .A(n6), .B(n19), .ZN(output0[14]) );
  XOR2_X1 U25 ( .A(DoubleBytes[7]), .B(input0[31]), .Z(n56) );
  XNOR2_X1 U26 ( .A(n56), .B(input0[23]), .ZN(n7) );
  XOR2_X1 U27 ( .A(input0[7]), .B(DoubleBytes[15]), .Z(n21) );
  XNOR2_X1 U28 ( .A(n7), .B(n21), .ZN(output0[15]) );
  XOR2_X1 U29 ( .A(DoubleBytes[8]), .B(input0[0]), .Z(n60) );
  XNOR2_X1 U30 ( .A(input0[24]), .B(n60), .ZN(n8) );
  XOR2_X1 U31 ( .A(input0[8]), .B(DoubleBytes[16]), .Z(n24) );
  XNOR2_X1 U32 ( .A(n8), .B(n24), .ZN(output0[16]) );
  XOR2_X1 U33 ( .A(DoubleBytes[9]), .B(input0[1]), .Z(n63) );
  XNOR2_X1 U34 ( .A(n63), .B(input0[25]), .ZN(n9) );
  XOR2_X1 U35 ( .A(DoubleBytes[17]), .B(input0[9]), .Z(n26) );
  XNOR2_X1 U36 ( .A(n9), .B(n26), .ZN(output0[17]) );
  XNOR2_X1 U37 ( .A(input0[26]), .B(n10), .ZN(n11) );
  XOR2_X1 U38 ( .A(input0[10]), .B(DoubleBytes[18]), .Z(n29) );
  XNOR2_X1 U39 ( .A(n11), .B(n29), .ZN(output0[18]) );
  XNOR2_X1 U40 ( .A(input0[27]), .B(n12), .ZN(n13) );
  XOR2_X1 U41 ( .A(input0[11]), .B(DoubleBytes[19]), .Z(n31) );
  XNOR2_X1 U42 ( .A(n13), .B(n31), .ZN(output0[19]) );
  XOR2_X1 U43 ( .A(input0[25]), .B(DoubleBytes[1]), .Z(n62) );
  XNOR2_X1 U44 ( .A(input0[9]), .B(n62), .ZN(n14) );
  XOR2_X1 U45 ( .A(input0[17]), .B(DoubleBytes[25]), .Z(n27) );
  XNOR2_X1 U46 ( .A(n14), .B(n27), .ZN(output0[1]) );
  XNOR2_X1 U47 ( .A(input0[28]), .B(n15), .ZN(n16) );
  XOR2_X1 U48 ( .A(input0[12]), .B(DoubleBytes[20]), .Z(n33) );
  XNOR2_X1 U49 ( .A(n16), .B(n33), .ZN(output0[20]) );
  XNOR2_X1 U50 ( .A(input0[29]), .B(n17), .ZN(n18) );
  XOR2_X1 U51 ( .A(input0[13]), .B(DoubleBytes[21]), .Z(n35) );
  XNOR2_X1 U52 ( .A(n18), .B(n35), .ZN(output0[21]) );
  XNOR2_X1 U53 ( .A(input0[30]), .B(n19), .ZN(n20) );
  XOR2_X1 U54 ( .A(input0[14]), .B(DoubleBytes[22]), .Z(n40) );
  XNOR2_X1 U55 ( .A(n20), .B(n40), .ZN(output0[22]) );
  XNOR2_X1 U56 ( .A(input0[31]), .B(n21), .ZN(n22) );
  XOR2_X1 U57 ( .A(input0[15]), .B(DoubleBytes[23]), .Z(n42) );
  XNOR2_X1 U58 ( .A(n22), .B(n42), .ZN(output0[23]) );
  XNOR2_X1 U59 ( .A(n23), .B(input0[0]), .ZN(n25) );
  XNOR2_X1 U60 ( .A(n25), .B(n24), .ZN(output0[24]) );
  XNOR2_X1 U61 ( .A(input0[1]), .B(n26), .ZN(n28) );
  XNOR2_X1 U62 ( .A(n28), .B(n27), .ZN(output0[25]) );
  XNOR2_X1 U63 ( .A(input0[2]), .B(n29), .ZN(n30) );
  XOR2_X1 U64 ( .A(input0[18]), .B(DoubleBytes[26]), .Z(n38) );
  XNOR2_X1 U65 ( .A(n30), .B(n38), .ZN(output0[26]) );
  XNOR2_X1 U66 ( .A(input0[3]), .B(n31), .ZN(n32) );
  XOR2_X1 U67 ( .A(input0[19]), .B(DoubleBytes[27]), .Z(n45) );
  XNOR2_X1 U68 ( .A(n32), .B(n45), .ZN(output0[27]) );
  XNOR2_X1 U69 ( .A(input0[4]), .B(n33), .ZN(n34) );
  XOR2_X1 U70 ( .A(input0[20]), .B(DoubleBytes[28]), .Z(n48) );
  XNOR2_X1 U71 ( .A(n34), .B(n48), .ZN(output0[28]) );
  XNOR2_X1 U72 ( .A(input0[5]), .B(n35), .ZN(n36) );
  XOR2_X1 U73 ( .A(input0[21]), .B(DoubleBytes[29]), .Z(n51) );
  XNOR2_X1 U74 ( .A(n36), .B(n51), .ZN(output0[29]) );
  XNOR2_X1 U75 ( .A(n37), .B(input0[10]), .ZN(n39) );
  XNOR2_X1 U76 ( .A(n39), .B(n38), .ZN(output0[2]) );
  XNOR2_X1 U77 ( .A(input0[6]), .B(n40), .ZN(n41) );
  XOR2_X1 U78 ( .A(input0[22]), .B(DoubleBytes[30]), .Z(n54) );
  XNOR2_X1 U79 ( .A(n41), .B(n54), .ZN(output0[30]) );
  XNOR2_X1 U80 ( .A(input0[7]), .B(n42), .ZN(n43) );
  XOR2_X1 U81 ( .A(input0[23]), .B(DoubleBytes[31]), .Z(n57) );
  XNOR2_X1 U82 ( .A(n43), .B(n57), .ZN(output0[31]) );
  XNOR2_X1 U83 ( .A(n44), .B(input0[11]), .ZN(n46) );
  XNOR2_X1 U84 ( .A(n46), .B(n45), .ZN(output0[3]) );
  XNOR2_X1 U85 ( .A(n47), .B(input0[12]), .ZN(n49) );
  XNOR2_X1 U86 ( .A(n49), .B(n48), .ZN(output0[4]) );
  XNOR2_X1 U87 ( .A(n50), .B(input0[13]), .ZN(n52) );
  XNOR2_X1 U88 ( .A(n52), .B(n51), .ZN(output0[5]) );
  XNOR2_X1 U89 ( .A(n53), .B(input0[14]), .ZN(n55) );
  XNOR2_X1 U90 ( .A(n55), .B(n54), .ZN(output0[6]) );
  XNOR2_X1 U91 ( .A(n56), .B(input0[15]), .ZN(n58) );
  XNOR2_X1 U92 ( .A(n58), .B(n57), .ZN(output0[7]) );
  XNOR2_X1 U93 ( .A(n59), .B(input0[16]), .ZN(n61) );
  XNOR2_X1 U94 ( .A(n61), .B(n60), .ZN(output0[8]) );
  XNOR2_X1 U95 ( .A(n63), .B(n62), .ZN(n64) );
  XNOR2_X1 U96 ( .A(n64), .B(input0[17]), .ZN(output0[9]) );
endmodule


module Mul2_4 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_3 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_2 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module Mul2_1 ( input0, output0 );
  input [7:0] input0;
  output [7:0] output0;

  assign output0[7] = input0[6];
  assign output0[6] = input0[5];
  assign output0[5] = input0[4];
  assign output0[2] = input0[1];
  assign output0[0] = input0[7];

  XOR2_X1 U1 ( .A(input0[7]), .B(input0[0]), .Z(output0[1]) );
  XOR2_X1 U2 ( .A(input0[7]), .B(input0[2]), .Z(output0[3]) );
  XOR2_X1 U3 ( .A(input0[7]), .B(input0[3]), .Z(output0[4]) );
endmodule


module MixOneColumn_1 ( input0, output0 );
  input [31:0] input0;
  output [31:0] output0;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  wire   [31:0] DoubleBytes;

  Mul2_4 Mul2Inst_0 ( .input0(input0[31:24]), .output0(DoubleBytes[31:24]) );
  Mul2_3 Mul2Inst_1 ( .input0(input0[23:16]), .output0(DoubleBytes[23:16]) );
  Mul2_2 Mul2Inst_2 ( .input0(input0[15:8]), .output0(DoubleBytes[15:8]) );
  Mul2_1 Mul2Inst_3 ( .input0(input0[7:0]), .output0(DoubleBytes[7:0]) );
  XOR2_X1 U1 ( .A(DoubleBytes[0]), .B(input0[24]), .Z(n59) );
  XOR2_X1 U2 ( .A(input0[16]), .B(DoubleBytes[24]), .Z(n23) );
  XNOR2_X1 U3 ( .A(n59), .B(n23), .ZN(n1) );
  XNOR2_X1 U4 ( .A(n1), .B(input0[8]), .ZN(output0[0]) );
  XOR2_X1 U5 ( .A(DoubleBytes[2]), .B(input0[26]), .Z(n37) );
  XNOR2_X1 U6 ( .A(n37), .B(input0[18]), .ZN(n2) );
  XOR2_X1 U7 ( .A(input0[2]), .B(DoubleBytes[10]), .Z(n10) );
  XNOR2_X1 U8 ( .A(n2), .B(n10), .ZN(output0[10]) );
  XOR2_X1 U9 ( .A(DoubleBytes[3]), .B(input0[27]), .Z(n44) );
  XNOR2_X1 U10 ( .A(n44), .B(input0[19]), .ZN(n3) );
  XOR2_X1 U11 ( .A(input0[3]), .B(DoubleBytes[11]), .Z(n12) );
  XNOR2_X1 U12 ( .A(n3), .B(n12), .ZN(output0[11]) );
  XOR2_X1 U13 ( .A(DoubleBytes[4]), .B(input0[28]), .Z(n47) );
  XNOR2_X1 U14 ( .A(n47), .B(input0[20]), .ZN(n4) );
  XOR2_X1 U15 ( .A(input0[4]), .B(DoubleBytes[12]), .Z(n15) );
  XNOR2_X1 U16 ( .A(n4), .B(n15), .ZN(output0[12]) );
  XOR2_X1 U17 ( .A(DoubleBytes[5]), .B(input0[29]), .Z(n50) );
  XNOR2_X1 U18 ( .A(n50), .B(input0[21]), .ZN(n5) );
  XOR2_X1 U19 ( .A(input0[5]), .B(DoubleBytes[13]), .Z(n17) );
  XNOR2_X1 U20 ( .A(n5), .B(n17), .ZN(output0[13]) );
  XOR2_X1 U21 ( .A(DoubleBytes[6]), .B(input0[30]), .Z(n53) );
  XNOR2_X1 U22 ( .A(n53), .B(input0[22]), .ZN(n6) );
  XOR2_X1 U23 ( .A(input0[6]), .B(DoubleBytes[14]), .Z(n19) );
  XNOR2_X1 U24 ( .A(n6), .B(n19), .ZN(output0[14]) );
  XOR2_X1 U25 ( .A(DoubleBytes[7]), .B(input0[31]), .Z(n56) );
  XNOR2_X1 U26 ( .A(n56), .B(input0[23]), .ZN(n7) );
  XOR2_X1 U27 ( .A(input0[7]), .B(DoubleBytes[15]), .Z(n21) );
  XNOR2_X1 U28 ( .A(n7), .B(n21), .ZN(output0[15]) );
  XOR2_X1 U29 ( .A(DoubleBytes[8]), .B(input0[0]), .Z(n60) );
  XNOR2_X1 U30 ( .A(input0[24]), .B(n60), .ZN(n8) );
  XOR2_X1 U31 ( .A(input0[8]), .B(DoubleBytes[16]), .Z(n24) );
  XNOR2_X1 U32 ( .A(n8), .B(n24), .ZN(output0[16]) );
  XOR2_X1 U33 ( .A(DoubleBytes[9]), .B(input0[1]), .Z(n63) );
  XNOR2_X1 U34 ( .A(n63), .B(input0[25]), .ZN(n9) );
  XOR2_X1 U35 ( .A(DoubleBytes[17]), .B(input0[9]), .Z(n26) );
  XNOR2_X1 U36 ( .A(n9), .B(n26), .ZN(output0[17]) );
  XNOR2_X1 U37 ( .A(input0[26]), .B(n10), .ZN(n11) );
  XOR2_X1 U38 ( .A(input0[10]), .B(DoubleBytes[18]), .Z(n29) );
  XNOR2_X1 U39 ( .A(n11), .B(n29), .ZN(output0[18]) );
  XNOR2_X1 U40 ( .A(input0[27]), .B(n12), .ZN(n13) );
  XOR2_X1 U41 ( .A(input0[11]), .B(DoubleBytes[19]), .Z(n31) );
  XNOR2_X1 U42 ( .A(n13), .B(n31), .ZN(output0[19]) );
  XOR2_X1 U43 ( .A(input0[25]), .B(DoubleBytes[1]), .Z(n62) );
  XNOR2_X1 U44 ( .A(input0[9]), .B(n62), .ZN(n14) );
  XOR2_X1 U45 ( .A(input0[17]), .B(DoubleBytes[25]), .Z(n27) );
  XNOR2_X1 U46 ( .A(n14), .B(n27), .ZN(output0[1]) );
  XNOR2_X1 U47 ( .A(input0[28]), .B(n15), .ZN(n16) );
  XOR2_X1 U48 ( .A(input0[12]), .B(DoubleBytes[20]), .Z(n33) );
  XNOR2_X1 U49 ( .A(n16), .B(n33), .ZN(output0[20]) );
  XNOR2_X1 U50 ( .A(input0[29]), .B(n17), .ZN(n18) );
  XOR2_X1 U51 ( .A(input0[13]), .B(DoubleBytes[21]), .Z(n35) );
  XNOR2_X1 U52 ( .A(n18), .B(n35), .ZN(output0[21]) );
  XNOR2_X1 U53 ( .A(input0[30]), .B(n19), .ZN(n20) );
  XOR2_X1 U54 ( .A(input0[14]), .B(DoubleBytes[22]), .Z(n40) );
  XNOR2_X1 U55 ( .A(n20), .B(n40), .ZN(output0[22]) );
  XNOR2_X1 U56 ( .A(input0[31]), .B(n21), .ZN(n22) );
  XOR2_X1 U57 ( .A(input0[15]), .B(DoubleBytes[23]), .Z(n42) );
  XNOR2_X1 U58 ( .A(n22), .B(n42), .ZN(output0[23]) );
  XNOR2_X1 U59 ( .A(n23), .B(input0[0]), .ZN(n25) );
  XNOR2_X1 U60 ( .A(n25), .B(n24), .ZN(output0[24]) );
  XNOR2_X1 U61 ( .A(input0[1]), .B(n26), .ZN(n28) );
  XNOR2_X1 U62 ( .A(n28), .B(n27), .ZN(output0[25]) );
  XNOR2_X1 U63 ( .A(input0[2]), .B(n29), .ZN(n30) );
  XOR2_X1 U64 ( .A(input0[18]), .B(DoubleBytes[26]), .Z(n38) );
  XNOR2_X1 U65 ( .A(n30), .B(n38), .ZN(output0[26]) );
  XNOR2_X1 U66 ( .A(input0[3]), .B(n31), .ZN(n32) );
  XOR2_X1 U67 ( .A(input0[19]), .B(DoubleBytes[27]), .Z(n45) );
  XNOR2_X1 U68 ( .A(n32), .B(n45), .ZN(output0[27]) );
  XNOR2_X1 U69 ( .A(input0[4]), .B(n33), .ZN(n34) );
  XOR2_X1 U70 ( .A(input0[20]), .B(DoubleBytes[28]), .Z(n48) );
  XNOR2_X1 U71 ( .A(n34), .B(n48), .ZN(output0[28]) );
  XNOR2_X1 U72 ( .A(input0[5]), .B(n35), .ZN(n36) );
  XOR2_X1 U73 ( .A(input0[21]), .B(DoubleBytes[29]), .Z(n51) );
  XNOR2_X1 U74 ( .A(n36), .B(n51), .ZN(output0[29]) );
  XNOR2_X1 U75 ( .A(n37), .B(input0[10]), .ZN(n39) );
  XNOR2_X1 U76 ( .A(n39), .B(n38), .ZN(output0[2]) );
  XNOR2_X1 U77 ( .A(input0[6]), .B(n40), .ZN(n41) );
  XOR2_X1 U78 ( .A(input0[22]), .B(DoubleBytes[30]), .Z(n54) );
  XNOR2_X1 U79 ( .A(n41), .B(n54), .ZN(output0[30]) );
  XNOR2_X1 U80 ( .A(input0[7]), .B(n42), .ZN(n43) );
  XOR2_X1 U81 ( .A(input0[23]), .B(DoubleBytes[31]), .Z(n57) );
  XNOR2_X1 U82 ( .A(n43), .B(n57), .ZN(output0[31]) );
  XNOR2_X1 U83 ( .A(n44), .B(input0[11]), .ZN(n46) );
  XNOR2_X1 U84 ( .A(n46), .B(n45), .ZN(output0[3]) );
  XNOR2_X1 U85 ( .A(n47), .B(input0[12]), .ZN(n49) );
  XNOR2_X1 U86 ( .A(n49), .B(n48), .ZN(output0[4]) );
  XNOR2_X1 U87 ( .A(n50), .B(input0[13]), .ZN(n52) );
  XNOR2_X1 U88 ( .A(n52), .B(n51), .ZN(output0[5]) );
  XNOR2_X1 U89 ( .A(n53), .B(input0[14]), .ZN(n55) );
  XNOR2_X1 U90 ( .A(n55), .B(n54), .ZN(output0[6]) );
  XNOR2_X1 U91 ( .A(n56), .B(input0[15]), .ZN(n58) );
  XNOR2_X1 U92 ( .A(n58), .B(n57), .ZN(output0[7]) );
  XNOR2_X1 U93 ( .A(n59), .B(input0[16]), .ZN(n61) );
  XNOR2_X1 U94 ( .A(n61), .B(n60), .ZN(output0[8]) );
  XNOR2_X1 U95 ( .A(n63), .B(n62), .ZN(n64) );
  XNOR2_X1 U96 ( .A(n64), .B(input0[17]), .ZN(output0[9]) );
endmodule


module MixColumns ( input0, output0 );
  input [127:0] input0;
  output [127:0] output0;


  MixOneColumn_0 MixOneColumnInst_0 ( .input0(input0[127:96]), .output0(
        output0[127:96]) );
  MixOneColumn_3 MixOneColumnInst_1 ( .input0(input0[95:64]), .output0(
        output0[95:64]) );
  MixOneColumn_2 MixOneColumnInst_2 ( .input0(input0[63:32]), .output0(
        output0[63:32]) );
  MixOneColumn_1 MixOneColumnInst_3 ( .input0(input0[31:0]), .output0(
        output0[31:0]) );
endmodule


module XOR_forMUX_256 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_128 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_255 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_128 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_256 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_128 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_255 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_128 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_128 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_128 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_128 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_128 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_128 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_254 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_127 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_253 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_127 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_254 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_127 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_253 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_127 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_127 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_127 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_127 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_127 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_127 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_252 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_126 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_251 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_126 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_252 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_126 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_251 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_126 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_126 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_126 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_126 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_126 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_126 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_250 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_125 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_249 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_125 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_250 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_125 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_249 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_125 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_125 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_125 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_125 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_125 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_125 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_248 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_124 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_247 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_124 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_248 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_124 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_247 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_124 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_124 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_124 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_124 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_124 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_124 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_246 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_123 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_245 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_123 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_246 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_123 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_245 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_123 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_123 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_123 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_123 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_123 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_123 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_244 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_122 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_243 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_122 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_244 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_122 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_243 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_122 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_122 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_122 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_122 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_122 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_122 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_242 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_121 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_241 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_121 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_242 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_121 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_241 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_121 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_121 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_121 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_121 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_121 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_121 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_240 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_120 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_239 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_120 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_240 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_120 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_239 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_120 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_120 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_120 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_120 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_120 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_120 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_238 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_119 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_237 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_119 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_238 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_119 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_237 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_119 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_119 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_119 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_119 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_119 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_119 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_236 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_118 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_235 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_118 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_236 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_118 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_235 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_118 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_118 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_118 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_118 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_118 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_118 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_234 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_117 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_233 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_117 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_234 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_117 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_233 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_117 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_117 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_117 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_117 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_117 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_117 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_232 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_116 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_231 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_116 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_232 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_116 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_231 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_116 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_116 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_116 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_116 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_116 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_116 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_230 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_115 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_229 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_115 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_230 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_115 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_229 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_115 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_115 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_115 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_115 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_115 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_115 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_228 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_114 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_227 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_114 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_228 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_114 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_227 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_114 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_114 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_114 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_114 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_114 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_114 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_226 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_113 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_225 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_113 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_226 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_113 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_225 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_113 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_113 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_113 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_113 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_113 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_113 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_224 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_112 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_223 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_112 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_224 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_112 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_223 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_112 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_112 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_112 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_112 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_112 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_112 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_222 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_111 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_221 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_111 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_222 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_111 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_221 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_111 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_111 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_111 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_111 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_111 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_111 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_220 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_110 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_219 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_110 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_220 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_110 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_219 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_110 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_110 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_110 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_110 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_110 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_110 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_218 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_109 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_217 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_109 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_218 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_109 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_217 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_109 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_109 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_109 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_109 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_109 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_109 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_216 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_108 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_215 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_108 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_216 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_108 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_215 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_108 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_108 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_108 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_108 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_108 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_108 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_214 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_107 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_213 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_107 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_214 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_107 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_213 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_107 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_107 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_107 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_107 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_107 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_107 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_212 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_106 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_211 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_106 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_212 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_106 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_211 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_106 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_106 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_106 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_106 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_106 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_106 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_210 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_105 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_209 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_105 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_210 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_105 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_209 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_105 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_105 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_105 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_105 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_105 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_105 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_208 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_104 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_207 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_104 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_208 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_104 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_207 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_104 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_104 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_104 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_104 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_104 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_104 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_206 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_103 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_205 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_103 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_206 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_103 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_205 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_103 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_103 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_103 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_103 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_103 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_103 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_204 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_102 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_203 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_102 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_204 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_102 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_203 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_102 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_102 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_102 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_102 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_102 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_102 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_202 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_101 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_201 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_101 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_202 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_101 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_201 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_101 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_101 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_101 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_101 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_101 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_101 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_200 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_100 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_199 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_100 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_200 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_100 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_199 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_100 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_100 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_100 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_100 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_100 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_100 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_198 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_99 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_197 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_99 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_198 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_99 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_197 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_99 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_99 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_99 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_99 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_99 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_99 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_196 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_98 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_195 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_98 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_196 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_98 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_195 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_98 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_98 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_98 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_98 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_98 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_98 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_194 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_97 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_193 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_97 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_194 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_97 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_193 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_97 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_97 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_97 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_97 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_97 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_97 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_192 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_96 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_191 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_96 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_192 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_96 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_191 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_96 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_96 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_96 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_96 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_96 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_96 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_190 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_95 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_189 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_95 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_190 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_95 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_189 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_95 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_95 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_95 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_95 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_95 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_95 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_188 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_94 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_187 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_94 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_188 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_94 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_187 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_94 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_94 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_94 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_94 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_94 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_94 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_186 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_93 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_185 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_93 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_186 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_93 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_185 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_93 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_93 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_93 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_93 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_93 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_93 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_184 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_92 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_183 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_92 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_184 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_92 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_183 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_92 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_92 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_92 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_92 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_92 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_92 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_182 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_91 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_181 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_91 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_182 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_91 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_181 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_91 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_91 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_91 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_91 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_91 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_91 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_180 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_90 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_179 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_90 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_180 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_90 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_179 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_90 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_90 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_90 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_90 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_90 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_90 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_178 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_89 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_177 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_89 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_178 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_89 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_177 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_89 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_89 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_89 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_89 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_89 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_89 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_176 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_88 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_175 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_88 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_176 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_88 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_175 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_88 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_88 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_88 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_88 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_88 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_88 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_174 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_87 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_173 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_87 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_174 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_87 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_173 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_87 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_87 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_87 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_87 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_87 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_87 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_172 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_86 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_171 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_86 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_172 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_86 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_171 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_86 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_86 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_86 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_86 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_86 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_86 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_170 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_85 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_169 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_85 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_170 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_85 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_169 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_85 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_85 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_85 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_85 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_85 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_85 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_168 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_84 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_167 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_84 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_168 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_84 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_167 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_84 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_84 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_84 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_84 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_84 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_84 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_166 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_83 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_165 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_83 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_166 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_83 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_165 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_83 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_83 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_83 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_83 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_83 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_83 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_164 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_82 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_163 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_82 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_164 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_82 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_163 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_82 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_82 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_82 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_82 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_82 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_82 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_162 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_81 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_161 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_81 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_162 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_81 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_161 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_81 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_81 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_81 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_81 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_81 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_81 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_160 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_80 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_159 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_80 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_160 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_80 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_159 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_80 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_80 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_80 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_80 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_80 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_80 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_158 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_79 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_157 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_79 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_158 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_79 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_157 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_79 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_79 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_79 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_79 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_79 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_79 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_156 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_78 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_155 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_78 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_156 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_78 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_155 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_78 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_78 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_78 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_78 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_78 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_78 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_154 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_77 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_153 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_77 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_154 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_77 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_153 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_77 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_77 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_77 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_77 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_77 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_77 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_152 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_76 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_151 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_76 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_152 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_76 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_151 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_76 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_76 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_76 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_76 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_76 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_76 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_150 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_75 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_149 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_75 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_150 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_75 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_149 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_75 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_75 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_75 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_75 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_75 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_75 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_148 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_74 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_147 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_74 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_148 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_74 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_147 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_74 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_74 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_74 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_74 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_74 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_74 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_146 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_73 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_145 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_73 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_146 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_73 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_145 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_73 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_73 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_73 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_73 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_73 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_73 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_144 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_72 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_143 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_72 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_144 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_72 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_143 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_72 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_72 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_72 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_72 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_72 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_72 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_142 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_71 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_141 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_71 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_142 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_71 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_141 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_71 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_71 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_71 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_71 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_71 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_71 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_140 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_70 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_139 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_70 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_140 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_70 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_139 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_70 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_70 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_70 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_70 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_70 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_70 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_138 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_69 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_137 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_69 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_138 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_69 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_137 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_69 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_69 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_69 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_69 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_69 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_69 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_136 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_68 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_135 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_68 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_136 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_68 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_135 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_68 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_68 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_68 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_68 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_68 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_68 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_134 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_67 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_133 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_67 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_134 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_67 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_133 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_67 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_67 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_67 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_67 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_67 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_67 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_132 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_66 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_131 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_66 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_132 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_66 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_131 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_66 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_66 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_66 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_66 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_66 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_66 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_130 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_65 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_129 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_65 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_130 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_65 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_129 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_65 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_65 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_65 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_65 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_65 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_65 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_128 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_64 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_127 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_64 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_128 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_64 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_127 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_64 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_64 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_64 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_64 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_64 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_64 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_126 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_63 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_125 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_63 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_126 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_63 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_125 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_63 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_63 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_63 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_63 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_63 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_63 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_124 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_62 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_123 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_62 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_124 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_62 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_123 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_62 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_62 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_62 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_62 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_62 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_62 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_122 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_61 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_121 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_61 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_122 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_61 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_121 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_61 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_61 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_61 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_61 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_61 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_61 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_120 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_60 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_119 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_60 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_120 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_60 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_119 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_60 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_60 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_60 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_60 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_60 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_60 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_118 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_59 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_117 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_59 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_118 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_59 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_117 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_59 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_59 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_59 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_59 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_59 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_59 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_116 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_58 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_115 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_58 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_116 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_58 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_115 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_58 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_58 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_58 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_58 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_58 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_58 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_114 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_57 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_113 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_57 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_114 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_57 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_113 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_57 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_57 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_57 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_57 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_57 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_57 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_112 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_56 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_111 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_56 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_112 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_56 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_111 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_56 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_56 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_56 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_56 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_56 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_56 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_110 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_55 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_109 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_55 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_110 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_55 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_109 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_55 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_55 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_55 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_55 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_55 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_55 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_108 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_54 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_107 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_54 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_108 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_54 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_107 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_54 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_54 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_54 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_54 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_54 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_54 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_106 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_53 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_105 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_53 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_106 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_53 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_105 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_53 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_53 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_53 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_53 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_53 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_53 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_104 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_52 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_103 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_52 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_104 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_52 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_103 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_52 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_52 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_52 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_52 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_52 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_52 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_102 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_51 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_101 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_51 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_102 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_51 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_101 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_51 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_51 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_51 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_51 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_51 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_51 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_100 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_50 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_99 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_50 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_100 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_50 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_99 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_50 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_50 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_50 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_50 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_50 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_50 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_98 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_49 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_97 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_49 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_98 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_49 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_97 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_49 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_49 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_49 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_49 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_49 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_49 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_96 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_48 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_95 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_48 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_96 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_48 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_95 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_48 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_48 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_48 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_48 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_48 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_48 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_94 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_47 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_93 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_47 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_94 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_47 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_93 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_47 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_47 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_47 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_47 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_47 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_47 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_92 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_46 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_91 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_46 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_92 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_46 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_91 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_46 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_46 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_46 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_46 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_46 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_46 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_90 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_45 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_89 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_45 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_90 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_45 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_89 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_45 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_45 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_45 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_45 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_45 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_45 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_88 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_44 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_87 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_44 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_88 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_44 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_87 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_44 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_44 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_44 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_44 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_44 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_44 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_86 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_43 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_85 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_43 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_86 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_43 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_85 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_43 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_43 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_43 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_43 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_43 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_43 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_84 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_42 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_83 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_42 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_84 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_42 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_83 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_42 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_42 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_42 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_42 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_42 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_42 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_82 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_41 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_81 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_41 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_82 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_41 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_81 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_41 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_41 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_41 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_41 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_41 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_41 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_80 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_40 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_79 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_40 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_80 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_40 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_79 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_40 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_40 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_40 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_40 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_40 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_40 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_78 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_39 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_77 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_39 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_78 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_39 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_77 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_39 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_39 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_39 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_39 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_39 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_39 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_76 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_38 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_75 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_38 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_76 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_38 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_75 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_38 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_38 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_38 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_38 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_38 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_38 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_74 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_37 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_73 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_37 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_74 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_37 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_73 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_37 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_37 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_37 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_37 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_37 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_37 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_72 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_36 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_71 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_36 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_72 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_36 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_71 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_36 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_36 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_36 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_36 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_36 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_36 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_70 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_35 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_69 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_35 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_70 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_35 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_69 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_35 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_35 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_35 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_35 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_35 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_35 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_68 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_34 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_67 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_34 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_68 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_34 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_67 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_34 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_34 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_34 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_34 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_34 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_34 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_66 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_33 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_65 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_33 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_66 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_33 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_65 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_33 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_33 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_33 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_33 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_33 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_33 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_64 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_32 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_63 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_32 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_64 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_32 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_63 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_32 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_32 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_32 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_32 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_32 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_32 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_62 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_31 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_61 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_31 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_62 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_31 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_61 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_31 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_31 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_31 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_31 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_31 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_31 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_60 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_30 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_59 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_30 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_60 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_30 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_59 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_30 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_30 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_30 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_30 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_30 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_30 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_58 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_29 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_57 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_29 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_58 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_29 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_57 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_29 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_29 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_29 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_29 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_29 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_29 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_56 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_28 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_55 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_28 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_56 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_28 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_55 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_28 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_28 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_28 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_28 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_28 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_28 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_54 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_27 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_53 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_27 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_54 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_27 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_53 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_27 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_27 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_27 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_27 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_27 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_27 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_52 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_26 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_51 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_26 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_52 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_26 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_51 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_26 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_26 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_26 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_26 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_26 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_26 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_50 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_25 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_49 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_25 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_50 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_25 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_49 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_25 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_25 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_25 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_25 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_25 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_25 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_48 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_24 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_47 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_24 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_48 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_24 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_47 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_24 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_24 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_24 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_24 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_24 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_24 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_46 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_23 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_45 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_23 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_46 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_23 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_45 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_23 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_23 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_23 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_23 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_23 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_23 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_44 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_22 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_43 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_22 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_44 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_22 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_43 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_22 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_22 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_22 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_22 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_22 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_22 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_42 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_21 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_41 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_21 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_42 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_21 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_41 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_21 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_21 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_21 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_21 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_21 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_21 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_40 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_20 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_39 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_20 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_40 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_20 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_39 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_20 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_20 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_20 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_20 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_20 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_20 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_38 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_19 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_37 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_19 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_38 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_19 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_37 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_19 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_19 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_19 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_19 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_19 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_19 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_36 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_18 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_35 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_18 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_36 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_18 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_35 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_18 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_18 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_18 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_18 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_18 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_18 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_34 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_17 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_33 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_17 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_34 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_17 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_33 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_17 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_17 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_17 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_17 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_17 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_17 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_32 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_16 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_31 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_16 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_32 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_16 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_31 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_16 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_16 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_16 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_16 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_16 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_16 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_30 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_15 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_29 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_15 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_30 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_15 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_29 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_15 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_15 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_15 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_15 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_15 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_15 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_28 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_14 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_27 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_14 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_28 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_14 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_27 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_14 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_14 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_14 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_14 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_14 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_14 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_26 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_13 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_25 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_13 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_26 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_13 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_25 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_13 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_13 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_13 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_13 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_13 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_13 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_24 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_12 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_23 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_12 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_24 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_12 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_23 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_12 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_12 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_12 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_12 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_12 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_12 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_22 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_11 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_21 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_11 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_22 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_11 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_21 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_11 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_11 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_11 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_11 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_11 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_11 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_20 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_10 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_19 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_10 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_20 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_10 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_19 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_10 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_10 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_10 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_10 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_10 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_10 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_18 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_9 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_17 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_9 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_18 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_9 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_17 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_9 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_9 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_9 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_9 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_9 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_9 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_16 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_8 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_15 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_8 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_16 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_8 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_15 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_8 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_8 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_8 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_8 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_8 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_8 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_14 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_7 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_13 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_7 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_14 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_7 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_13 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_7 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_7 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_7 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_7 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_7 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_7 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_12 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_6 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_11 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_6 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_12 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_6 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_11 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_6 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_6 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_6 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_6 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_6 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_6 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_10 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_5 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_9 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_5 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_10 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_5 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_9 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_5 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_5 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_5 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_5 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_5 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_5 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_8 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_4 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_7 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_4 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_8 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_4 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_7 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_4 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_4 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_4 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_4 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_4 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_4 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_6 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_3 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_5 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_3 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_6 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_3 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_5 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_3 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_3 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_3 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_3 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_3 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_3 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_4 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_2 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_3 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_2 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_4 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_2 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_3 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_2 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_2 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_2 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_2 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_2 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_2 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module XOR_forMUX_2 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module AND_forMUX_1 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module XOR_forMUX_1 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MUX_1bit_1 ( S, D0, D1, Q );
  input S, D0, D1;
  output Q;
  wire   X, Y;

  XOR_forMUX_2 XOR1 ( .A(D0), .B(D1), .C(X) );
  AND_forMUX_1 AND1 ( .A(S), .B(X), .C(Y) );
  XOR_forMUX_1 XOR2 ( .A(Y), .B(D0), .C(Q) );
endmodule


module MyDFFs_1 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_1 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_1 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module ff_SDE_1 ( clk, D0, D1, sel, Q );
  input clk, D0, D1, sel;
  output Q;
  wire   next_state;

  MUX_1bit_1 MUX_inst ( .S(sel), .D0(D0), .D1(D1), .Q(next_state) );
  MyDFF_1 current_state_reg ( .D(next_state), .CK(clk), .Q(Q), .QN() );
endmodule


module reg_SDE_size128_1 ( clk, D0, D1, sel, Q );
  input [127:0] D0;
  input [127:0] D1;
  output [127:0] Q;
  input clk, sel;
  wire   n6, n7, n8, n9, n10;

  ff_SDE_128 Inst_ff_SDE_0 ( .clk(clk), .D0(D0[0]), .D1(D1[0]), .sel(n8), .Q(
        Q[0]) );
  ff_SDE_127 Inst_ff_SDE_1 ( .clk(clk), .D0(D0[1]), .D1(D1[1]), .sel(n9), .Q(
        Q[1]) );
  ff_SDE_126 Inst_ff_SDE_2 ( .clk(clk), .D0(D0[2]), .D1(D1[2]), .sel(n6), .Q(
        Q[2]) );
  ff_SDE_125 Inst_ff_SDE_3 ( .clk(clk), .D0(D0[3]), .D1(D1[3]), .sel(n7), .Q(
        Q[3]) );
  ff_SDE_124 Inst_ff_SDE_4 ( .clk(clk), .D0(D0[4]), .D1(D1[4]), .sel(n6), .Q(
        Q[4]) );
  ff_SDE_123 Inst_ff_SDE_5 ( .clk(clk), .D0(D0[5]), .D1(D1[5]), .sel(n7), .Q(
        Q[5]) );
  ff_SDE_122 Inst_ff_SDE_6 ( .clk(clk), .D0(D0[6]), .D1(D1[6]), .sel(n8), .Q(
        Q[6]) );
  ff_SDE_121 Inst_ff_SDE_7 ( .clk(clk), .D0(D0[7]), .D1(D1[7]), .sel(n6), .Q(
        Q[7]) );
  ff_SDE_120 Inst_ff_SDE_8 ( .clk(clk), .D0(D0[8]), .D1(D1[8]), .sel(n7), .Q(
        Q[8]) );
  ff_SDE_119 Inst_ff_SDE_9 ( .clk(clk), .D0(D0[9]), .D1(D1[9]), .sel(n8), .Q(
        Q[9]) );
  ff_SDE_118 Inst_ff_SDE_10 ( .clk(clk), .D0(D0[10]), .D1(D1[10]), .sel(n9), 
        .Q(Q[10]) );
  ff_SDE_117 Inst_ff_SDE_11 ( .clk(clk), .D0(D0[11]), .D1(D1[11]), .sel(n7), 
        .Q(Q[11]) );
  ff_SDE_116 Inst_ff_SDE_12 ( .clk(clk), .D0(D0[12]), .D1(D1[12]), .sel(n6), 
        .Q(Q[12]) );
  ff_SDE_115 Inst_ff_SDE_13 ( .clk(clk), .D0(D0[13]), .D1(D1[13]), .sel(n6), 
        .Q(Q[13]) );
  ff_SDE_114 Inst_ff_SDE_14 ( .clk(clk), .D0(D0[14]), .D1(D1[14]), .sel(n9), 
        .Q(Q[14]) );
  ff_SDE_113 Inst_ff_SDE_15 ( .clk(clk), .D0(D0[15]), .D1(D1[15]), .sel(n8), 
        .Q(Q[15]) );
  ff_SDE_112 Inst_ff_SDE_16 ( .clk(clk), .D0(D0[16]), .D1(D1[16]), .sel(n7), 
        .Q(Q[16]) );
  ff_SDE_111 Inst_ff_SDE_17 ( .clk(clk), .D0(D0[17]), .D1(D1[17]), .sel(n8), 
        .Q(Q[17]) );
  ff_SDE_110 Inst_ff_SDE_18 ( .clk(clk), .D0(D0[18]), .D1(D1[18]), .sel(n9), 
        .Q(Q[18]) );
  ff_SDE_109 Inst_ff_SDE_19 ( .clk(clk), .D0(D0[19]), .D1(D1[19]), .sel(n8), 
        .Q(Q[19]) );
  ff_SDE_108 Inst_ff_SDE_20 ( .clk(clk), .D0(D0[20]), .D1(D1[20]), .sel(n9), 
        .Q(Q[20]) );
  ff_SDE_107 Inst_ff_SDE_21 ( .clk(clk), .D0(D0[21]), .D1(D1[21]), .sel(n6), 
        .Q(Q[21]) );
  ff_SDE_106 Inst_ff_SDE_22 ( .clk(clk), .D0(D0[22]), .D1(D1[22]), .sel(n7), 
        .Q(Q[22]) );
  ff_SDE_105 Inst_ff_SDE_23 ( .clk(clk), .D0(D0[23]), .D1(D1[23]), .sel(n6), 
        .Q(Q[23]) );
  ff_SDE_104 Inst_ff_SDE_24 ( .clk(clk), .D0(D0[24]), .D1(D1[24]), .sel(n7), 
        .Q(Q[24]) );
  ff_SDE_103 Inst_ff_SDE_25 ( .clk(clk), .D0(D0[25]), .D1(D1[25]), .sel(n8), 
        .Q(Q[25]) );
  ff_SDE_102 Inst_ff_SDE_26 ( .clk(clk), .D0(D0[26]), .D1(D1[26]), .sel(n9), 
        .Q(Q[26]) );
  ff_SDE_101 Inst_ff_SDE_27 ( .clk(clk), .D0(D0[27]), .D1(D1[27]), .sel(n7), 
        .Q(Q[27]) );
  ff_SDE_100 Inst_ff_SDE_28 ( .clk(clk), .D0(D0[28]), .D1(D1[28]), .sel(n6), 
        .Q(Q[28]) );
  ff_SDE_99 Inst_ff_SDE_29 ( .clk(clk), .D0(D0[29]), .D1(D1[29]), .sel(n8), 
        .Q(Q[29]) );
  ff_SDE_98 Inst_ff_SDE_30 ( .clk(clk), .D0(D0[30]), .D1(D1[30]), .sel(n9), 
        .Q(Q[30]) );
  ff_SDE_97 Inst_ff_SDE_31 ( .clk(clk), .D0(D0[31]), .D1(D1[31]), .sel(n7), 
        .Q(Q[31]) );
  ff_SDE_96 Inst_ff_SDE_32 ( .clk(clk), .D0(D0[32]), .D1(D1[32]), .sel(n9), 
        .Q(Q[32]) );
  ff_SDE_95 Inst_ff_SDE_33 ( .clk(clk), .D0(D0[33]), .D1(D1[33]), .sel(n7), 
        .Q(Q[33]) );
  ff_SDE_94 Inst_ff_SDE_34 ( .clk(clk), .D0(D0[34]), .D1(D1[34]), .sel(n8), 
        .Q(Q[34]) );
  ff_SDE_93 Inst_ff_SDE_35 ( .clk(clk), .D0(D0[35]), .D1(D1[35]), .sel(n7), 
        .Q(Q[35]) );
  ff_SDE_92 Inst_ff_SDE_36 ( .clk(clk), .D0(D0[36]), .D1(D1[36]), .sel(n8), 
        .Q(Q[36]) );
  ff_SDE_91 Inst_ff_SDE_37 ( .clk(clk), .D0(D0[37]), .D1(D1[37]), .sel(n9), 
        .Q(Q[37]) );
  ff_SDE_90 Inst_ff_SDE_38 ( .clk(clk), .D0(D0[38]), .D1(D1[38]), .sel(n8), 
        .Q(Q[38]) );
  ff_SDE_89 Inst_ff_SDE_39 ( .clk(clk), .D0(D0[39]), .D1(D1[39]), .sel(n9), 
        .Q(Q[39]) );
  ff_SDE_88 Inst_ff_SDE_40 ( .clk(clk), .D0(D0[40]), .D1(D1[40]), .sel(n7), 
        .Q(Q[40]) );
  ff_SDE_87 Inst_ff_SDE_41 ( .clk(clk), .D0(D0[41]), .D1(D1[41]), .sel(n8), 
        .Q(Q[41]) );
  ff_SDE_86 Inst_ff_SDE_42 ( .clk(clk), .D0(D0[42]), .D1(D1[42]), .sel(n9), 
        .Q(Q[42]) );
  ff_SDE_85 Inst_ff_SDE_43 ( .clk(clk), .D0(D0[43]), .D1(D1[43]), .sel(n9), 
        .Q(Q[43]) );
  ff_SDE_84 Inst_ff_SDE_44 ( .clk(clk), .D0(D0[44]), .D1(D1[44]), .sel(n7), 
        .Q(Q[44]) );
  ff_SDE_83 Inst_ff_SDE_45 ( .clk(clk), .D0(D0[45]), .D1(D1[45]), .sel(n7), 
        .Q(Q[45]) );
  ff_SDE_82 Inst_ff_SDE_46 ( .clk(clk), .D0(D0[46]), .D1(D1[46]), .sel(n8), 
        .Q(Q[46]) );
  ff_SDE_81 Inst_ff_SDE_47 ( .clk(clk), .D0(D0[47]), .D1(D1[47]), .sel(n9), 
        .Q(Q[47]) );
  ff_SDE_80 Inst_ff_SDE_48 ( .clk(clk), .D0(D0[48]), .D1(D1[48]), .sel(n8), 
        .Q(Q[48]) );
  ff_SDE_79 Inst_ff_SDE_49 ( .clk(clk), .D0(D0[49]), .D1(D1[49]), .sel(n7), 
        .Q(Q[49]) );
  ff_SDE_78 Inst_ff_SDE_50 ( .clk(clk), .D0(D0[50]), .D1(D1[50]), .sel(n8), 
        .Q(Q[50]) );
  ff_SDE_77 Inst_ff_SDE_51 ( .clk(clk), .D0(D0[51]), .D1(D1[51]), .sel(n9), 
        .Q(Q[51]) );
  ff_SDE_76 Inst_ff_SDE_52 ( .clk(clk), .D0(D0[52]), .D1(D1[52]), .sel(n9), 
        .Q(Q[52]) );
  ff_SDE_75 Inst_ff_SDE_53 ( .clk(clk), .D0(D0[53]), .D1(D1[53]), .sel(n7), 
        .Q(Q[53]) );
  ff_SDE_74 Inst_ff_SDE_54 ( .clk(clk), .D0(D0[54]), .D1(D1[54]), .sel(n8), 
        .Q(Q[54]) );
  ff_SDE_73 Inst_ff_SDE_55 ( .clk(clk), .D0(D0[55]), .D1(D1[55]), .sel(n9), 
        .Q(Q[55]) );
  ff_SDE_72 Inst_ff_SDE_56 ( .clk(clk), .D0(D0[56]), .D1(D1[56]), .sel(n7), 
        .Q(Q[56]) );
  ff_SDE_71 Inst_ff_SDE_57 ( .clk(clk), .D0(D0[57]), .D1(D1[57]), .sel(n8), 
        .Q(Q[57]) );
  ff_SDE_70 Inst_ff_SDE_58 ( .clk(clk), .D0(D0[58]), .D1(D1[58]), .sel(n9), 
        .Q(Q[58]) );
  ff_SDE_69 Inst_ff_SDE_59 ( .clk(clk), .D0(D0[59]), .D1(D1[59]), .sel(n6), 
        .Q(Q[59]) );
  ff_SDE_68 Inst_ff_SDE_60 ( .clk(clk), .D0(D0[60]), .D1(D1[60]), .sel(sel), 
        .Q(Q[60]) );
  ff_SDE_67 Inst_ff_SDE_61 ( .clk(clk), .D0(D0[61]), .D1(D1[61]), .sel(sel), 
        .Q(Q[61]) );
  ff_SDE_66 Inst_ff_SDE_62 ( .clk(clk), .D0(D0[62]), .D1(D1[62]), .sel(n6), 
        .Q(Q[62]) );
  ff_SDE_65 Inst_ff_SDE_63 ( .clk(clk), .D0(D0[63]), .D1(D1[63]), .sel(n6), 
        .Q(Q[63]) );
  ff_SDE_64 Inst_ff_SDE_64 ( .clk(clk), .D0(D0[64]), .D1(D1[64]), .sel(n6), 
        .Q(Q[64]) );
  ff_SDE_63 Inst_ff_SDE_65 ( .clk(clk), .D0(D0[65]), .D1(D1[65]), .sel(n6), 
        .Q(Q[65]) );
  ff_SDE_62 Inst_ff_SDE_66 ( .clk(clk), .D0(D0[66]), .D1(D1[66]), .sel(n6), 
        .Q(Q[66]) );
  ff_SDE_61 Inst_ff_SDE_67 ( .clk(clk), .D0(D0[67]), .D1(D1[67]), .sel(n6), 
        .Q(Q[67]) );
  ff_SDE_60 Inst_ff_SDE_68 ( .clk(clk), .D0(D0[68]), .D1(D1[68]), .sel(n9), 
        .Q(Q[68]) );
  ff_SDE_59 Inst_ff_SDE_69 ( .clk(clk), .D0(D0[69]), .D1(D1[69]), .sel(n9), 
        .Q(Q[69]) );
  ff_SDE_58 Inst_ff_SDE_70 ( .clk(clk), .D0(D0[70]), .D1(D1[70]), .sel(n9), 
        .Q(Q[70]) );
  ff_SDE_57 Inst_ff_SDE_71 ( .clk(clk), .D0(D0[71]), .D1(D1[71]), .sel(n9), 
        .Q(Q[71]) );
  ff_SDE_56 Inst_ff_SDE_72 ( .clk(clk), .D0(D0[72]), .D1(D1[72]), .sel(n9), 
        .Q(Q[72]) );
  ff_SDE_55 Inst_ff_SDE_73 ( .clk(clk), .D0(D0[73]), .D1(D1[73]), .sel(n9), 
        .Q(Q[73]) );
  ff_SDE_54 Inst_ff_SDE_74 ( .clk(clk), .D0(D0[74]), .D1(D1[74]), .sel(n9), 
        .Q(Q[74]) );
  ff_SDE_53 Inst_ff_SDE_75 ( .clk(clk), .D0(D0[75]), .D1(D1[75]), .sel(n9), 
        .Q(Q[75]) );
  ff_SDE_52 Inst_ff_SDE_76 ( .clk(clk), .D0(D0[76]), .D1(D1[76]), .sel(n9), 
        .Q(Q[76]) );
  ff_SDE_51 Inst_ff_SDE_77 ( .clk(clk), .D0(D0[77]), .D1(D1[77]), .sel(n9), 
        .Q(Q[77]) );
  ff_SDE_50 Inst_ff_SDE_78 ( .clk(clk), .D0(D0[78]), .D1(D1[78]), .sel(n9), 
        .Q(Q[78]) );
  ff_SDE_49 Inst_ff_SDE_79 ( .clk(clk), .D0(D0[79]), .D1(D1[79]), .sel(n9), 
        .Q(Q[79]) );
  ff_SDE_48 Inst_ff_SDE_80 ( .clk(clk), .D0(D0[80]), .D1(D1[80]), .sel(n8), 
        .Q(Q[80]) );
  ff_SDE_47 Inst_ff_SDE_81 ( .clk(clk), .D0(D0[81]), .D1(D1[81]), .sel(n8), 
        .Q(Q[81]) );
  ff_SDE_46 Inst_ff_SDE_82 ( .clk(clk), .D0(D0[82]), .D1(D1[82]), .sel(n8), 
        .Q(Q[82]) );
  ff_SDE_45 Inst_ff_SDE_83 ( .clk(clk), .D0(D0[83]), .D1(D1[83]), .sel(n8), 
        .Q(Q[83]) );
  ff_SDE_44 Inst_ff_SDE_84 ( .clk(clk), .D0(D0[84]), .D1(D1[84]), .sel(n8), 
        .Q(Q[84]) );
  ff_SDE_43 Inst_ff_SDE_85 ( .clk(clk), .D0(D0[85]), .D1(D1[85]), .sel(n8), 
        .Q(Q[85]) );
  ff_SDE_42 Inst_ff_SDE_86 ( .clk(clk), .D0(D0[86]), .D1(D1[86]), .sel(n8), 
        .Q(Q[86]) );
  ff_SDE_41 Inst_ff_SDE_87 ( .clk(clk), .D0(D0[87]), .D1(D1[87]), .sel(n8), 
        .Q(Q[87]) );
  ff_SDE_40 Inst_ff_SDE_88 ( .clk(clk), .D0(D0[88]), .D1(D1[88]), .sel(n8), 
        .Q(Q[88]) );
  ff_SDE_39 Inst_ff_SDE_89 ( .clk(clk), .D0(D0[89]), .D1(D1[89]), .sel(n8), 
        .Q(Q[89]) );
  ff_SDE_38 Inst_ff_SDE_90 ( .clk(clk), .D0(D0[90]), .D1(D1[90]), .sel(n8), 
        .Q(Q[90]) );
  ff_SDE_37 Inst_ff_SDE_91 ( .clk(clk), .D0(D0[91]), .D1(D1[91]), .sel(n8), 
        .Q(Q[91]) );
  ff_SDE_36 Inst_ff_SDE_92 ( .clk(clk), .D0(D0[92]), .D1(D1[92]), .sel(n7), 
        .Q(Q[92]) );
  ff_SDE_35 Inst_ff_SDE_93 ( .clk(clk), .D0(D0[93]), .D1(D1[93]), .sel(n7), 
        .Q(Q[93]) );
  ff_SDE_34 Inst_ff_SDE_94 ( .clk(clk), .D0(D0[94]), .D1(D1[94]), .sel(n7), 
        .Q(Q[94]) );
  ff_SDE_33 Inst_ff_SDE_95 ( .clk(clk), .D0(D0[95]), .D1(D1[95]), .sel(n7), 
        .Q(Q[95]) );
  ff_SDE_32 Inst_ff_SDE_96 ( .clk(clk), .D0(D0[96]), .D1(D1[96]), .sel(n7), 
        .Q(Q[96]) );
  ff_SDE_31 Inst_ff_SDE_97 ( .clk(clk), .D0(D0[97]), .D1(D1[97]), .sel(n7), 
        .Q(Q[97]) );
  ff_SDE_30 Inst_ff_SDE_98 ( .clk(clk), .D0(D0[98]), .D1(D1[98]), .sel(n7), 
        .Q(Q[98]) );
  ff_SDE_29 Inst_ff_SDE_99 ( .clk(clk), .D0(D0[99]), .D1(D1[99]), .sel(n7), 
        .Q(Q[99]) );
  ff_SDE_28 Inst_ff_SDE_100 ( .clk(clk), .D0(D0[100]), .D1(D1[100]), .sel(n7), 
        .Q(Q[100]) );
  ff_SDE_27 Inst_ff_SDE_101 ( .clk(clk), .D0(D0[101]), .D1(D1[101]), .sel(n7), 
        .Q(Q[101]) );
  ff_SDE_26 Inst_ff_SDE_102 ( .clk(clk), .D0(D0[102]), .D1(D1[102]), .sel(n7), 
        .Q(Q[102]) );
  ff_SDE_25 Inst_ff_SDE_103 ( .clk(clk), .D0(D0[103]), .D1(D1[103]), .sel(n7), 
        .Q(Q[103]) );
  ff_SDE_24 Inst_ff_SDE_104 ( .clk(clk), .D0(D0[104]), .D1(D1[104]), .sel(n7), 
        .Q(Q[104]) );
  ff_SDE_23 Inst_ff_SDE_105 ( .clk(clk), .D0(D0[105]), .D1(D1[105]), .sel(n8), 
        .Q(Q[105]) );
  ff_SDE_22 Inst_ff_SDE_106 ( .clk(clk), .D0(D0[106]), .D1(D1[106]), .sel(n9), 
        .Q(Q[106]) );
  ff_SDE_21 Inst_ff_SDE_107 ( .clk(clk), .D0(D0[107]), .D1(D1[107]), .sel(n6), 
        .Q(Q[107]) );
  ff_SDE_20 Inst_ff_SDE_108 ( .clk(clk), .D0(D0[108]), .D1(D1[108]), .sel(n6), 
        .Q(Q[108]) );
  ff_SDE_19 Inst_ff_SDE_109 ( .clk(clk), .D0(D0[109]), .D1(D1[109]), .sel(n7), 
        .Q(Q[109]) );
  ff_SDE_18 Inst_ff_SDE_110 ( .clk(clk), .D0(D0[110]), .D1(D1[110]), .sel(n8), 
        .Q(Q[110]) );
  ff_SDE_17 Inst_ff_SDE_111 ( .clk(clk), .D0(D0[111]), .D1(D1[111]), .sel(n9), 
        .Q(Q[111]) );
  ff_SDE_16 Inst_ff_SDE_112 ( .clk(clk), .D0(D0[112]), .D1(D1[112]), .sel(n7), 
        .Q(Q[112]) );
  ff_SDE_15 Inst_ff_SDE_113 ( .clk(clk), .D0(D0[113]), .D1(D1[113]), .sel(n8), 
        .Q(Q[113]) );
  ff_SDE_14 Inst_ff_SDE_114 ( .clk(clk), .D0(D0[114]), .D1(D1[114]), .sel(n9), 
        .Q(Q[114]) );
  ff_SDE_13 Inst_ff_SDE_115 ( .clk(clk), .D0(D0[115]), .D1(D1[115]), .sel(n6), 
        .Q(Q[115]) );
  ff_SDE_12 Inst_ff_SDE_116 ( .clk(clk), .D0(D0[116]), .D1(D1[116]), .sel(n6), 
        .Q(Q[116]) );
  ff_SDE_11 Inst_ff_SDE_117 ( .clk(clk), .D0(D0[117]), .D1(D1[117]), .sel(n6), 
        .Q(Q[117]) );
  ff_SDE_10 Inst_ff_SDE_118 ( .clk(clk), .D0(D0[118]), .D1(D1[118]), .sel(n6), 
        .Q(Q[118]) );
  ff_SDE_9 Inst_ff_SDE_119 ( .clk(clk), .D0(D0[119]), .D1(D1[119]), .sel(n6), 
        .Q(Q[119]) );
  ff_SDE_8 Inst_ff_SDE_120 ( .clk(clk), .D0(D0[120]), .D1(D1[120]), .sel(n6), 
        .Q(Q[120]) );
  ff_SDE_7 Inst_ff_SDE_121 ( .clk(clk), .D0(D0[121]), .D1(D1[121]), .sel(n6), 
        .Q(Q[121]) );
  ff_SDE_6 Inst_ff_SDE_122 ( .clk(clk), .D0(D0[122]), .D1(D1[122]), .sel(n6), 
        .Q(Q[122]) );
  ff_SDE_5 Inst_ff_SDE_123 ( .clk(clk), .D0(D0[123]), .D1(D1[123]), .sel(n6), 
        .Q(Q[123]) );
  ff_SDE_4 Inst_ff_SDE_124 ( .clk(clk), .D0(D0[124]), .D1(D1[124]), .sel(n6), 
        .Q(Q[124]) );
  ff_SDE_3 Inst_ff_SDE_125 ( .clk(clk), .D0(D0[125]), .D1(D1[125]), .sel(n6), 
        .Q(Q[125]) );
  ff_SDE_2 Inst_ff_SDE_126 ( .clk(clk), .D0(D0[126]), .D1(D1[126]), .sel(n6), 
        .Q(Q[126]) );
  ff_SDE_1 Inst_ff_SDE_127 ( .clk(clk), .D0(D0[127]), .D1(D1[127]), .sel(n6), 
        .Q(Q[127]) );
  INV_X1 U1 ( .A(n10), .ZN(n6) );
  INV_X1 U2 ( .A(n10), .ZN(n7) );
  INV_X1 U3 ( .A(n10), .ZN(n8) );
  INV_X1 U4 ( .A(n10), .ZN(n9) );
  INV_X1 U5 ( .A(sel), .ZN(n10) );
endmodule


module MyXOR_360 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_359 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_358 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_357 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_356 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_355 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_354 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_353 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_352 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_351 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_350 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_349 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_348 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_347 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_346 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_345 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_344 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_343 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_342 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_341 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_340 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_339 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_338 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_337 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_336 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_335 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_334 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_136 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_135 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_333 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_134 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_332 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_133 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_132 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_331 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_131 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_330 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_130 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_129 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_329 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_128 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_328 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_327 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_326 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_325 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_324 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_323 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_322 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_321 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_320 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_319 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_127 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_318 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_317 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_316 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_126 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_125 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_124 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_123 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_315 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_122 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_121 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_314 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_313 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_312 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_311 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_310 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_309 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_308 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_307 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_306 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_305 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_120 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_119 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_118 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_117 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_116 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_115 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_114 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_113 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_112 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_111 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_110 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_109 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_108 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_107 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_106 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_105 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_104 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_103 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_304 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_303 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_302 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_301 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_300 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_299 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_298 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_297 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_296 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_295 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_294 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_293 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_292 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_291 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_290 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_289 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_288 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_287 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_286 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_285 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_284 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_283 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_282 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_281 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_280 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_279 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_278 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_277 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_276 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_275 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_274 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_16 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_15 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_273 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_272 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_271 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_14 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_13 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_4 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_360 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_359 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_358 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_357 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_356 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_355 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_354 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_353 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_352 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_351 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_350 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_349 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_348 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_347 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_346 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_345 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_344 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_343 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_342 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_341 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_340 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_339 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_338 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_337 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_336 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_335 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_334 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_136 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_135 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_333 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_134 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_332 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_133 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_132 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_331 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_131 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_330 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_130 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_129 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_329 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_128 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_328 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_327 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_326 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_325 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_324 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_323 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_322 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_321 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_320 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_319 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_127 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_318 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_317 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_316 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_126 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_125 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_124 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_123 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_315 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_122 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_121 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_314 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_313 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_312 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_311 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_310 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_309 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_308 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_307 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_306 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_305 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_120 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_119 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_118 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_117 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_116 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_115 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_114 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_113 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_112 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_111 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_110 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_109 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_108 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_107 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_106 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_105 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_104 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_103 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_304 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_303 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_302 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_301 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_300 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_299 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_298 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_297 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_296 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_295 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_294 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_293 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_292 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_291 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_290 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_289 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_288 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_287 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_286 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_285 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_284 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_283 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_282 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_281 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_280 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_279 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_278 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_277 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_276 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_275 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_274 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_16 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_15 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_273 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_272 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_271 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_14 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_13 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_270 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_269 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_268 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_267 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_266 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_265 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_264 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_263 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_262 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_261 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_260 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_259 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_258 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_257 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_256 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_255 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_254 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_253 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_252 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_251 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_250 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_249 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_248 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_247 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_246 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_245 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_244 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_102 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_101 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_243 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_100 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_242 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_99 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_98 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_241 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_97 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_240 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_96 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_95 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_239 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_94 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_238 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_237 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_236 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_235 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_234 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_233 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_232 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_231 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_230 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_229 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_93 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_228 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_227 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_226 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_92 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_91 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_90 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_89 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_225 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_88 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_87 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_224 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_223 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_222 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_221 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_220 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_219 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_218 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_217 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_216 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_215 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_86 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_85 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_84 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_83 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_82 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_81 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_80 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_79 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_78 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_77 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_76 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_75 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_74 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_73 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_72 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_71 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_70 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_69 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_214 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_213 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_212 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_211 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_210 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_209 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_208 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_207 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_206 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_205 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_204 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_203 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_202 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_201 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_200 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_199 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_198 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_197 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_196 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_195 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_194 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_193 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_192 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_191 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_190 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_189 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_188 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_187 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_186 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_185 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_184 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_12 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_11 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_183 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_182 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_181 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_10 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_9 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_3 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_270 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_269 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_268 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_267 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_266 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_265 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_264 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_263 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_262 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_261 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_260 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_259 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_258 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_257 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_256 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_255 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_254 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_253 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_252 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_251 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_250 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_249 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_248 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_247 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_246 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_245 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_244 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_102 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_101 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_243 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_100 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_242 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_99 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_98 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_241 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_97 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_240 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_96 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_95 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_239 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_94 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_238 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_237 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_236 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_235 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_234 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_233 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_232 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_231 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_230 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_229 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_93 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_228 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_227 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_226 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_92 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_91 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_90 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_89 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_225 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_88 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_87 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_224 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_223 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_222 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_221 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_220 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_219 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_218 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_217 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_216 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_215 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_86 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_85 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_84 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_83 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_82 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_81 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_80 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_79 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_78 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_77 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_76 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_75 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_74 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_73 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_72 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_71 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_70 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_69 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_214 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_213 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_212 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_211 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_210 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_209 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_208 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_207 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_206 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_205 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_204 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_203 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_202 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_201 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_200 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_199 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_198 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_197 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_196 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_195 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_194 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_193 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_192 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_191 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_190 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_189 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_188 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_187 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_186 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_185 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_184 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_12 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_11 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_183 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_182 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_181 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_10 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_9 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_180 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_179 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_178 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_177 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_176 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_175 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_174 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_173 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_172 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_171 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_170 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_169 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_168 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_167 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_166 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_165 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_164 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_163 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_162 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_161 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_160 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_159 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_158 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_157 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_156 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_155 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_154 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_68 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_67 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_153 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_66 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_152 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_65 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_64 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_151 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_63 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_150 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_62 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_61 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_149 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_60 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_148 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_147 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_146 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_145 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_144 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_143 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_142 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_141 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_140 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_139 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_59 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_138 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_137 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_136 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_58 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_57 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_56 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_55 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_135 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_54 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_53 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_134 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_133 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_132 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_131 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_130 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_129 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_128 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_127 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_126 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_125 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_52 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_51 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_50 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_49 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_48 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_47 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_46 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_45 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_44 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_43 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_42 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_41 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_40 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_39 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_38 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_37 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_36 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_35 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_124 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_123 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_122 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_121 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_120 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_119 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_118 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_117 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_116 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_115 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_114 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_113 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_112 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_111 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_110 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_109 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_108 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_107 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_106 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_105 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_104 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_103 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_102 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_101 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_100 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_99 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_98 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_97 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_96 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_95 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_94 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_8 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_7 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_93 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_92 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_91 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_6 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_5 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_2 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_180 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_179 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_178 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_177 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_176 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_175 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_174 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_173 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_172 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_171 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_170 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_169 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_168 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_167 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_166 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_165 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_164 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_163 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_162 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_161 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_160 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_159 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_158 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_157 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_156 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_155 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_154 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_68 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_67 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_153 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_66 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_152 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_65 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_64 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_151 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_63 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_150 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_62 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_61 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_149 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_60 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_148 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_147 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_146 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_145 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_144 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_143 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_142 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_141 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_140 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_139 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_59 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_138 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_137 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_136 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_58 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_57 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_56 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_55 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_135 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_54 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_53 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_134 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_133 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_132 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_131 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_130 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_129 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_128 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_127 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_126 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_125 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_52 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_51 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_50 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_49 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_48 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_47 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_46 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_45 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_44 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_43 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_42 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_41 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_40 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_39 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_38 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_37 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_36 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_35 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_124 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_123 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_122 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_121 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_120 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_119 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_118 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_117 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_116 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_115 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_114 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_113 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_112 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_111 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_110 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_109 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_108 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_107 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_106 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_105 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_104 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_103 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_102 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_101 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_100 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_99 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_98 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_97 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_96 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_95 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_94 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_8 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_7 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_93 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_92 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_91 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_6 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_5 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module MyXOR_90 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_89 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_88 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_87 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_86 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_85 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_84 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_83 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_82 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_81 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_80 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_79 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_78 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_77 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_76 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_75 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_74 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_73 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_72 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_71 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_70 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_69 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_68 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_67 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_66 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_65 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_64 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_34 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_33 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_63 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_32 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_62 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_31 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_30 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_61 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_29 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_60 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_28 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_27 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_59 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_26 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_58 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_57 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_56 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_55 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_54 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_53 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_52 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_51 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_50 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_49 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_25 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_48 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_47 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_46 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_24 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_23 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_22 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_21 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_45 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_20 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_19 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_44 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_43 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_42 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_41 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_40 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_39 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_38 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_37 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_36 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_35 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyAND_18 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_17 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_16 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_15 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_14 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_13 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_12 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_11 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_10 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_9 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_8 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_7 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_6 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_5 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_4 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_3 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_2 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyAND_1 ( A, B, C );
  input A, B;
  output C;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(C) );
endmodule


module MyXOR_34 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_33 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_32 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_31 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_30 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_29 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_28 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_27 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_26 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_25 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_24 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_23 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_22 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_21 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_20 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_19 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_18 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_17 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_16 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_15 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_14 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_13 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_12 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_11 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_10 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_9 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_8 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_7 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_6 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_5 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_4 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_4 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_3 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXOR_3 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_2 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXOR_1 ( A, B, C );
  input A, B;
  output C;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(C) );
endmodule


module MyXNOR_2 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module MyXNOR_1 ( A, B, C );
  input A, B;
  output C;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(C) );
endmodule


module Sbox_1 ( x, y );
  input [7:0] x;
  output [7:0] y;
  wire   T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16,
         T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, M1, M2, M3, M4,
         M5, M6, M7, M8, M9, M10, M11, M12, M13, M14, M15, M16, M17, M18, M19,
         M20, M21, M22, M23, M24, M25, M26, M27, M28, M29, M30, M31, M32, M33,
         M34, M35, M36, M37, M38, M39, M40, M41, M42, M43, M44, M45, M46, M47,
         M48, M49, M50, M51, M52, M53, M54, M55, M56, M57, M58, M59, M60, M61,
         M62, M63, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13,
         L14, L15, L16, L17, L18, L19, L20, L21, L22, L23, L24, L25, L26, L27,
         L28, L29;

  MyXOR_90 XOR_T1 ( .A(x[7]), .B(x[4]), .C(T1) );
  MyXOR_89 XOR_T2 ( .A(x[7]), .B(x[2]), .C(T2) );
  MyXOR_88 XOR_T3 ( .A(x[7]), .B(x[1]), .C(T3) );
  MyXOR_87 XOR_T4 ( .A(x[4]), .B(x[2]), .C(T4) );
  MyXOR_86 XOR_T5 ( .A(x[3]), .B(x[1]), .C(T5) );
  MyXOR_85 XOR_T6 ( .A(T1), .B(T5), .C(T6) );
  MyXOR_84 XOR_T7 ( .A(x[6]), .B(x[5]), .C(T7) );
  MyXOR_83 XOR_T8 ( .A(x[0]), .B(T6), .C(T8) );
  MyXOR_82 XOR_T9 ( .A(x[0]), .B(T7), .C(T9) );
  MyXOR_81 XOR_T10 ( .A(T6), .B(T7), .C(T10) );
  MyXOR_80 XOR_T11 ( .A(x[6]), .B(x[2]), .C(T11) );
  MyXOR_79 XOR_T12 ( .A(x[5]), .B(x[2]), .C(T12) );
  MyXOR_78 XOR_T13 ( .A(T3), .B(T4), .C(T13) );
  MyXOR_77 XOR_T14 ( .A(T6), .B(T11), .C(T14) );
  MyXOR_76 XOR_T15 ( .A(T5), .B(T11), .C(T15) );
  MyXOR_75 XOR_T16 ( .A(T5), .B(T12), .C(T16) );
  MyXOR_74 XOR_T17 ( .A(T9), .B(T16), .C(T17) );
  MyXOR_73 XOR_T18 ( .A(x[4]), .B(x[0]), .C(T18) );
  MyXOR_72 XOR_T19 ( .A(T7), .B(T18), .C(T19) );
  MyXOR_71 XOR_T20 ( .A(T1), .B(T19), .C(T20) );
  MyXOR_70 XOR_T21 ( .A(x[1]), .B(x[0]), .C(T21) );
  MyXOR_69 XOR_T22 ( .A(T7), .B(T21), .C(T22) );
  MyXOR_68 XOR_T23 ( .A(T2), .B(T22), .C(T23) );
  MyXOR_67 XOR_T24 ( .A(T2), .B(T10), .C(T24) );
  MyXOR_66 XOR_T25 ( .A(T20), .B(T17), .C(T25) );
  MyXOR_65 XOR_T26 ( .A(T3), .B(T16), .C(T26) );
  MyXOR_64 XOR_T27 ( .A(T1), .B(T12), .C(T27) );
  MyAND_34 AND_M1 ( .A(T13), .B(T6), .C(M1) );
  MyAND_33 AND_M2 ( .A(T23), .B(T8), .C(M2) );
  MyXOR_63 XOR_M3 ( .A(T14), .B(M1), .C(M3) );
  MyAND_32 AND_M4 ( .A(T19), .B(x[0]), .C(M4) );
  MyXOR_62 XOR_M5 ( .A(M4), .B(M1), .C(M5) );
  MyAND_31 AND_M6 ( .A(T3), .B(T16), .C(M6) );
  MyAND_30 AND_M7 ( .A(T22), .B(T9), .C(M7) );
  MyXOR_61 XOR_M8 ( .A(T26), .B(M6), .C(M8) );
  MyAND_29 AND_M9 ( .A(T20), .B(T17), .C(M9) );
  MyXOR_60 XOR_M10 ( .A(M9), .B(M6), .C(M10) );
  MyAND_28 AND_M11 ( .A(T1), .B(T15), .C(M11) );
  MyAND_27 AND_M12 ( .A(T4), .B(T27), .C(M12) );
  MyXOR_59 XOR_M13 ( .A(M12), .B(M11), .C(M13) );
  MyAND_26 AND_M14 ( .A(T2), .B(T10), .C(M14) );
  MyXOR_58 XOR_M15 ( .A(M14), .B(M11), .C(M15) );
  MyXOR_57 XOR_M16 ( .A(M3), .B(M2), .C(M16) );
  MyXOR_56 XOR_M17 ( .A(M5), .B(T24), .C(M17) );
  MyXOR_55 XOR_M18 ( .A(M8), .B(M7), .C(M18) );
  MyXOR_54 XOR_M19 ( .A(M10), .B(M15), .C(M19) );
  MyXOR_53 XOR_M20 ( .A(M16), .B(M13), .C(M20) );
  MyXOR_52 XOR_M21 ( .A(M17), .B(M15), .C(M21) );
  MyXOR_51 XOR_M22 ( .A(M18), .B(M13), .C(M22) );
  MyXOR_50 XOR_M23 ( .A(M19), .B(T25), .C(M23) );
  MyXOR_49 XOR_M24 ( .A(M22), .B(M23), .C(M24) );
  MyAND_25 AND_M25 ( .A(M22), .B(M20), .C(M25) );
  MyXOR_48 XOR_M26 ( .A(M21), .B(M25), .C(M26) );
  MyXOR_47 XOR_M27 ( .A(M20), .B(M21), .C(M27) );
  MyXOR_46 XOR_M28 ( .A(M23), .B(M25), .C(M28) );
  MyAND_24 AND_M29 ( .A(M28), .B(M27), .C(M29) );
  MyAND_23 AND_M30 ( .A(M26), .B(M24), .C(M30) );
  MyAND_22 AND_M31 ( .A(M20), .B(M23), .C(M31) );
  MyAND_21 AND_M32 ( .A(M27), .B(M31), .C(M32) );
  MyXOR_45 XOR_M33 ( .A(M27), .B(M25), .C(M33) );
  MyAND_20 AND_M34 ( .A(M21), .B(M22), .C(M34) );
  MyAND_19 AND_M35 ( .A(M24), .B(M34), .C(M35) );
  MyXOR_44 XOR_M36 ( .A(M24), .B(M25), .C(M36) );
  MyXOR_43 XOR_M37 ( .A(M21), .B(M29), .C(M37) );
  MyXOR_42 XOR_M38 ( .A(M32), .B(M33), .C(M38) );
  MyXOR_41 XOR_M39 ( .A(M23), .B(M30), .C(M39) );
  MyXOR_40 XOR_M40 ( .A(M35), .B(M36), .C(M40) );
  MyXOR_39 XOR_M41 ( .A(M38), .B(M40), .C(M41) );
  MyXOR_38 XOR_M42 ( .A(M37), .B(M39), .C(M42) );
  MyXOR_37 XOR_M43 ( .A(M37), .B(M38), .C(M43) );
  MyXOR_36 XOR_M44 ( .A(M39), .B(M40), .C(M44) );
  MyXOR_35 XOR_M45 ( .A(M42), .B(M41), .C(M45) );
  MyAND_18 AND_M46 ( .A(M44), .B(T6), .C(M46) );
  MyAND_17 AND_M47 ( .A(M40), .B(T8), .C(M47) );
  MyAND_16 AND_M48 ( .A(M39), .B(x[0]), .C(M48) );
  MyAND_15 AND_M49 ( .A(M43), .B(T16), .C(M49) );
  MyAND_14 AND_M50 ( .A(M38), .B(T9), .C(M50) );
  MyAND_13 AND_M51 ( .A(M37), .B(T17), .C(M51) );
  MyAND_12 AND_M52 ( .A(M42), .B(T15), .C(M52) );
  MyAND_11 AND_M53 ( .A(M45), .B(T27), .C(M53) );
  MyAND_10 AND_M54 ( .A(M41), .B(T10), .C(M54) );
  MyAND_9 AND_M55 ( .A(M44), .B(T13), .C(M55) );
  MyAND_8 AND_M56 ( .A(M40), .B(T23), .C(M56) );
  MyAND_7 AND_M57 ( .A(M39), .B(T19), .C(M57) );
  MyAND_6 AND_M58 ( .A(M43), .B(T3), .C(M58) );
  MyAND_5 AND_M59 ( .A(M38), .B(T22), .C(M59) );
  MyAND_4 AND_M60 ( .A(M37), .B(T20), .C(M60) );
  MyAND_3 AND_M61 ( .A(M42), .B(T1), .C(M61) );
  MyAND_2 AND_M62 ( .A(M45), .B(T4), .C(M62) );
  MyAND_1 AND_M63 ( .A(M41), .B(T2), .C(M63) );
  MyXOR_34 XOR_L0 ( .A(M61), .B(M62), .C(L0) );
  MyXOR_33 XOR_L1 ( .A(M50), .B(M56), .C(L1) );
  MyXOR_32 XOR_L2 ( .A(M46), .B(M48), .C(L2) );
  MyXOR_31 XOR_L3 ( .A(M47), .B(M55), .C(L3) );
  MyXOR_30 XOR_L4 ( .A(M54), .B(M58), .C(L4) );
  MyXOR_29 XOR_L5 ( .A(M49), .B(M61), .C(L5) );
  MyXOR_28 XOR_L6 ( .A(M62), .B(L5), .C(L6) );
  MyXOR_27 XOR_L7 ( .A(M46), .B(L3), .C(L7) );
  MyXOR_26 XOR_L8 ( .A(M51), .B(M59), .C(L8) );
  MyXOR_25 XOR_L9 ( .A(M52), .B(M53), .C(L9) );
  MyXOR_24 XOR_L10 ( .A(M53), .B(L4), .C(L10) );
  MyXOR_23 XOR_L11 ( .A(M60), .B(L2), .C(L11) );
  MyXOR_22 XOR_L12 ( .A(M48), .B(M51), .C(L12) );
  MyXOR_21 XOR_L13 ( .A(M50), .B(L0), .C(L13) );
  MyXOR_20 XOR_L14 ( .A(M52), .B(M61), .C(L14) );
  MyXOR_19 XOR_L15 ( .A(M55), .B(L1), .C(L15) );
  MyXOR_18 XOR_L16 ( .A(M56), .B(L0), .C(L16) );
  MyXOR_17 XOR_L17 ( .A(M57), .B(L1), .C(L17) );
  MyXOR_16 XOR_L18 ( .A(M58), .B(L8), .C(L18) );
  MyXOR_15 XOR_L19 ( .A(M63), .B(L4), .C(L19) );
  MyXOR_14 XOR_L20 ( .A(L0), .B(L1), .C(L20) );
  MyXOR_13 XOR_L21 ( .A(L1), .B(L7), .C(L21) );
  MyXOR_12 XOR_L22 ( .A(L3), .B(L12), .C(L22) );
  MyXOR_11 XOR_L23 ( .A(L18), .B(L2), .C(L23) );
  MyXOR_10 XOR_L24 ( .A(L15), .B(L9), .C(L24) );
  MyXOR_9 XOR_L25 ( .A(L6), .B(L10), .C(L25) );
  MyXOR_8 XOR_L26 ( .A(L7), .B(L9), .C(L26) );
  MyXOR_7 XOR_L27 ( .A(L8), .B(L10), .C(L27) );
  MyXOR_6 XOR_L28 ( .A(L11), .B(L14), .C(L28) );
  MyXOR_5 XOR_L29 ( .A(L11), .B(L17), .C(L29) );
  MyXOR_4 XOR_S0 ( .A(L6), .B(L24), .C(y[7]) );
  MyXNOR_4 XOR_S1 ( .A(L16), .B(L26), .C(y[6]) );
  MyXNOR_3 XOR_S2 ( .A(L19), .B(L28), .C(y[5]) );
  MyXOR_3 XOR_S3 ( .A(L6), .B(L21), .C(y[4]) );
  MyXOR_2 XOR_S4 ( .A(L20), .B(L22), .C(y[3]) );
  MyXOR_1 XOR_S5 ( .A(L25), .B(L29), .C(y[2]) );
  MyXNOR_2 XOR_S6 ( .A(L13), .B(L27), .C(y[1]) );
  MyXNOR_1 XOR_S7 ( .A(L6), .B(L23), .C(y[0]) );
endmodule


module KeySchedCore ( input0, Rcon, output0 );
  input [31:0] input0;
  input [7:0] Rcon;
  output [31:0] output0;
  wire   OutBytes_0__7_, OutBytes_0__6_, OutBytes_0__5_, OutBytes_0__4_,
         OutBytes_0__3_, OutBytes_0__2_, OutBytes_0__1_, OutBytes_0__0_;

  Sbox_4 Inst_Sbox_0 ( .x(input0[23:16]), .y({OutBytes_0__7_, OutBytes_0__6_, 
        OutBytes_0__5_, OutBytes_0__4_, OutBytes_0__3_, OutBytes_0__2_, 
        OutBytes_0__1_, OutBytes_0__0_}) );
  Sbox_3 Inst_Sbox_1 ( .x(input0[15:8]), .y(output0[23:16]) );
  Sbox_2 Inst_Sbox_2 ( .x(input0[7:0]), .y(output0[15:8]) );
  Sbox_1 Inst_Sbox_3 ( .x(input0[31:24]), .y(output0[7:0]) );
  XOR2_X1 U1 ( .A(OutBytes_0__0_), .B(Rcon[0]), .Z(output0[24]) );
  XOR2_X1 U2 ( .A(OutBytes_0__1_), .B(Rcon[1]), .Z(output0[25]) );
  XOR2_X1 U3 ( .A(OutBytes_0__2_), .B(Rcon[2]), .Z(output0[26]) );
  XOR2_X1 U4 ( .A(OutBytes_0__3_), .B(Rcon[3]), .Z(output0[27]) );
  XOR2_X1 U5 ( .A(OutBytes_0__4_), .B(Rcon[4]), .Z(output0[28]) );
  XOR2_X1 U6 ( .A(OutBytes_0__5_), .B(Rcon[5]), .Z(output0[29]) );
  XOR2_X1 U7 ( .A(OutBytes_0__6_), .B(Rcon[6]), .Z(output0[30]) );
  XOR2_X1 U8 ( .A(OutBytes_0__7_), .B(Rcon[7]), .Z(output0[31]) );
endmodule


module KeyExpansion ( input0, Rcon, output0 );
  input [127:0] input0;
  input [7:0] Rcon;
  output [127:0] output0;

  wire   [31:0] tmp;

  KeySchedCore KeySchedCoreInst ( .input0(input0[31:0]), .Rcon(Rcon), 
        .output0(tmp) );
  XOR2_X1 U1 ( .A(input0[96]), .B(tmp[0]), .Z(output0[96]) );
  XOR2_X1 U2 ( .A(input0[64]), .B(output0[96]), .Z(output0[64]) );
  XOR2_X1 U3 ( .A(input0[32]), .B(output0[64]), .Z(output0[32]) );
  XOR2_X1 U4 ( .A(input0[0]), .B(output0[32]), .Z(output0[0]) );
  XOR2_X1 U5 ( .A(input0[100]), .B(tmp[4]), .Z(output0[100]) );
  XOR2_X1 U6 ( .A(input0[101]), .B(tmp[5]), .Z(output0[101]) );
  XOR2_X1 U7 ( .A(input0[102]), .B(tmp[6]), .Z(output0[102]) );
  XOR2_X1 U8 ( .A(input0[103]), .B(tmp[7]), .Z(output0[103]) );
  XOR2_X1 U9 ( .A(input0[104]), .B(tmp[8]), .Z(output0[104]) );
  XOR2_X1 U10 ( .A(input0[105]), .B(tmp[9]), .Z(output0[105]) );
  XOR2_X1 U11 ( .A(input0[106]), .B(tmp[10]), .Z(output0[106]) );
  XOR2_X1 U12 ( .A(input0[107]), .B(tmp[11]), .Z(output0[107]) );
  XOR2_X1 U13 ( .A(input0[108]), .B(tmp[12]), .Z(output0[108]) );
  XOR2_X1 U14 ( .A(input0[109]), .B(tmp[13]), .Z(output0[109]) );
  XOR2_X1 U15 ( .A(input0[74]), .B(output0[106]), .Z(output0[74]) );
  XOR2_X1 U16 ( .A(input0[42]), .B(output0[74]), .Z(output0[42]) );
  XOR2_X1 U17 ( .A(input0[10]), .B(output0[42]), .Z(output0[10]) );
  XOR2_X1 U18 ( .A(input0[110]), .B(tmp[14]), .Z(output0[110]) );
  XOR2_X1 U19 ( .A(input0[111]), .B(tmp[15]), .Z(output0[111]) );
  XOR2_X1 U20 ( .A(input0[112]), .B(tmp[16]), .Z(output0[112]) );
  XOR2_X1 U21 ( .A(input0[113]), .B(tmp[17]), .Z(output0[113]) );
  XOR2_X1 U22 ( .A(input0[114]), .B(tmp[18]), .Z(output0[114]) );
  XOR2_X1 U23 ( .A(input0[115]), .B(tmp[19]), .Z(output0[115]) );
  XOR2_X1 U24 ( .A(input0[116]), .B(tmp[20]), .Z(output0[116]) );
  XOR2_X1 U25 ( .A(input0[117]), .B(tmp[21]), .Z(output0[117]) );
  XOR2_X1 U26 ( .A(input0[118]), .B(tmp[22]), .Z(output0[118]) );
  XOR2_X1 U27 ( .A(input0[119]), .B(tmp[23]), .Z(output0[119]) );
  XOR2_X1 U28 ( .A(input0[75]), .B(output0[107]), .Z(output0[75]) );
  XOR2_X1 U29 ( .A(input0[43]), .B(output0[75]), .Z(output0[43]) );
  XOR2_X1 U30 ( .A(input0[11]), .B(output0[43]), .Z(output0[11]) );
  XOR2_X1 U31 ( .A(input0[120]), .B(tmp[24]), .Z(output0[120]) );
  XOR2_X1 U32 ( .A(input0[121]), .B(tmp[25]), .Z(output0[121]) );
  XOR2_X1 U33 ( .A(input0[122]), .B(tmp[26]), .Z(output0[122]) );
  XOR2_X1 U34 ( .A(input0[123]), .B(tmp[27]), .Z(output0[123]) );
  XOR2_X1 U35 ( .A(input0[124]), .B(tmp[28]), .Z(output0[124]) );
  XOR2_X1 U36 ( .A(input0[125]), .B(tmp[29]), .Z(output0[125]) );
  XOR2_X1 U37 ( .A(input0[126]), .B(tmp[30]), .Z(output0[126]) );
  XOR2_X1 U38 ( .A(input0[127]), .B(tmp[31]), .Z(output0[127]) );
  XOR2_X1 U39 ( .A(input0[76]), .B(output0[108]), .Z(output0[76]) );
  XOR2_X1 U40 ( .A(input0[44]), .B(output0[76]), .Z(output0[44]) );
  XOR2_X1 U41 ( .A(input0[12]), .B(output0[44]), .Z(output0[12]) );
  XOR2_X1 U42 ( .A(input0[77]), .B(output0[109]), .Z(output0[77]) );
  XOR2_X1 U43 ( .A(input0[45]), .B(output0[77]), .Z(output0[45]) );
  XOR2_X1 U44 ( .A(input0[13]), .B(output0[45]), .Z(output0[13]) );
  XOR2_X1 U45 ( .A(input0[78]), .B(output0[110]), .Z(output0[78]) );
  XOR2_X1 U46 ( .A(input0[46]), .B(output0[78]), .Z(output0[46]) );
  XOR2_X1 U47 ( .A(input0[14]), .B(output0[46]), .Z(output0[14]) );
  XOR2_X1 U48 ( .A(input0[79]), .B(output0[111]), .Z(output0[79]) );
  XOR2_X1 U49 ( .A(input0[47]), .B(output0[79]), .Z(output0[47]) );
  XOR2_X1 U50 ( .A(input0[15]), .B(output0[47]), .Z(output0[15]) );
  XOR2_X1 U51 ( .A(input0[80]), .B(output0[112]), .Z(output0[80]) );
  XOR2_X1 U52 ( .A(input0[48]), .B(output0[80]), .Z(output0[48]) );
  XOR2_X1 U53 ( .A(input0[16]), .B(output0[48]), .Z(output0[16]) );
  XOR2_X1 U54 ( .A(input0[81]), .B(output0[113]), .Z(output0[81]) );
  XOR2_X1 U55 ( .A(input0[49]), .B(output0[81]), .Z(output0[49]) );
  XOR2_X1 U56 ( .A(input0[17]), .B(output0[49]), .Z(output0[17]) );
  XOR2_X1 U57 ( .A(input0[82]), .B(output0[114]), .Z(output0[82]) );
  XOR2_X1 U58 ( .A(input0[50]), .B(output0[82]), .Z(output0[50]) );
  XOR2_X1 U59 ( .A(input0[18]), .B(output0[50]), .Z(output0[18]) );
  XOR2_X1 U60 ( .A(input0[83]), .B(output0[115]), .Z(output0[83]) );
  XOR2_X1 U61 ( .A(input0[51]), .B(output0[83]), .Z(output0[51]) );
  XOR2_X1 U62 ( .A(input0[19]), .B(output0[51]), .Z(output0[19]) );
  XOR2_X1 U63 ( .A(input0[97]), .B(tmp[1]), .Z(output0[97]) );
  XOR2_X1 U64 ( .A(input0[65]), .B(output0[97]), .Z(output0[65]) );
  XOR2_X1 U65 ( .A(input0[33]), .B(output0[65]), .Z(output0[33]) );
  XOR2_X1 U66 ( .A(input0[1]), .B(output0[33]), .Z(output0[1]) );
  XOR2_X1 U67 ( .A(input0[84]), .B(output0[116]), .Z(output0[84]) );
  XOR2_X1 U68 ( .A(input0[52]), .B(output0[84]), .Z(output0[52]) );
  XOR2_X1 U69 ( .A(input0[20]), .B(output0[52]), .Z(output0[20]) );
  XOR2_X1 U70 ( .A(input0[85]), .B(output0[117]), .Z(output0[85]) );
  XOR2_X1 U71 ( .A(input0[53]), .B(output0[85]), .Z(output0[53]) );
  XOR2_X1 U72 ( .A(input0[21]), .B(output0[53]), .Z(output0[21]) );
  XOR2_X1 U73 ( .A(input0[86]), .B(output0[118]), .Z(output0[86]) );
  XOR2_X1 U74 ( .A(input0[54]), .B(output0[86]), .Z(output0[54]) );
  XOR2_X1 U75 ( .A(input0[22]), .B(output0[54]), .Z(output0[22]) );
  XOR2_X1 U76 ( .A(input0[87]), .B(output0[119]), .Z(output0[87]) );
  XOR2_X1 U77 ( .A(input0[55]), .B(output0[87]), .Z(output0[55]) );
  XOR2_X1 U78 ( .A(input0[23]), .B(output0[55]), .Z(output0[23]) );
  XOR2_X1 U79 ( .A(input0[88]), .B(output0[120]), .Z(output0[88]) );
  XOR2_X1 U80 ( .A(input0[56]), .B(output0[88]), .Z(output0[56]) );
  XOR2_X1 U81 ( .A(input0[24]), .B(output0[56]), .Z(output0[24]) );
  XOR2_X1 U82 ( .A(input0[89]), .B(output0[121]), .Z(output0[89]) );
  XOR2_X1 U83 ( .A(input0[57]), .B(output0[89]), .Z(output0[57]) );
  XOR2_X1 U84 ( .A(input0[25]), .B(output0[57]), .Z(output0[25]) );
  XOR2_X1 U85 ( .A(input0[90]), .B(output0[122]), .Z(output0[90]) );
  XOR2_X1 U86 ( .A(input0[58]), .B(output0[90]), .Z(output0[58]) );
  XOR2_X1 U87 ( .A(input0[26]), .B(output0[58]), .Z(output0[26]) );
  XOR2_X1 U88 ( .A(input0[91]), .B(output0[123]), .Z(output0[91]) );
  XOR2_X1 U89 ( .A(input0[59]), .B(output0[91]), .Z(output0[59]) );
  XOR2_X1 U90 ( .A(input0[27]), .B(output0[59]), .Z(output0[27]) );
  XOR2_X1 U91 ( .A(input0[92]), .B(output0[124]), .Z(output0[92]) );
  XOR2_X1 U92 ( .A(input0[60]), .B(output0[92]), .Z(output0[60]) );
  XOR2_X1 U93 ( .A(input0[28]), .B(output0[60]), .Z(output0[28]) );
  XOR2_X1 U94 ( .A(input0[93]), .B(output0[125]), .Z(output0[93]) );
  XOR2_X1 U95 ( .A(input0[61]), .B(output0[93]), .Z(output0[61]) );
  XOR2_X1 U96 ( .A(input0[29]), .B(output0[61]), .Z(output0[29]) );
  XOR2_X1 U97 ( .A(input0[98]), .B(tmp[2]), .Z(output0[98]) );
  XOR2_X1 U98 ( .A(input0[66]), .B(output0[98]), .Z(output0[66]) );
  XOR2_X1 U99 ( .A(input0[34]), .B(output0[66]), .Z(output0[34]) );
  XOR2_X1 U100 ( .A(input0[2]), .B(output0[34]), .Z(output0[2]) );
  XOR2_X1 U101 ( .A(input0[94]), .B(output0[126]), .Z(output0[94]) );
  XOR2_X1 U102 ( .A(input0[62]), .B(output0[94]), .Z(output0[62]) );
  XOR2_X1 U103 ( .A(input0[30]), .B(output0[62]), .Z(output0[30]) );
  XOR2_X1 U104 ( .A(input0[95]), .B(output0[127]), .Z(output0[95]) );
  XOR2_X1 U105 ( .A(input0[63]), .B(output0[95]), .Z(output0[63]) );
  XOR2_X1 U106 ( .A(input0[31]), .B(output0[63]), .Z(output0[31]) );
  XOR2_X1 U107 ( .A(input0[99]), .B(tmp[3]), .Z(output0[99]) );
  XOR2_X1 U108 ( .A(input0[67]), .B(output0[99]), .Z(output0[67]) );
  XOR2_X1 U109 ( .A(input0[35]), .B(output0[67]), .Z(output0[35]) );
  XOR2_X1 U110 ( .A(input0[68]), .B(output0[100]), .Z(output0[68]) );
  XOR2_X1 U111 ( .A(input0[36]), .B(output0[68]), .Z(output0[36]) );
  XOR2_X1 U112 ( .A(input0[69]), .B(output0[101]), .Z(output0[69]) );
  XOR2_X1 U113 ( .A(input0[37]), .B(output0[69]), .Z(output0[37]) );
  XOR2_X1 U114 ( .A(input0[70]), .B(output0[102]), .Z(output0[70]) );
  XOR2_X1 U115 ( .A(input0[38]), .B(output0[70]), .Z(output0[38]) );
  XOR2_X1 U116 ( .A(input0[71]), .B(output0[103]), .Z(output0[71]) );
  XOR2_X1 U117 ( .A(input0[39]), .B(output0[71]), .Z(output0[39]) );
  XOR2_X1 U118 ( .A(input0[3]), .B(output0[35]), .Z(output0[3]) );
  XOR2_X1 U119 ( .A(input0[72]), .B(output0[104]), .Z(output0[72]) );
  XOR2_X1 U120 ( .A(input0[40]), .B(output0[72]), .Z(output0[40]) );
  XOR2_X1 U121 ( .A(input0[73]), .B(output0[105]), .Z(output0[73]) );
  XOR2_X1 U122 ( .A(input0[41]), .B(output0[73]), .Z(output0[41]) );
  XOR2_X1 U123 ( .A(input0[4]), .B(output0[36]), .Z(output0[4]) );
  XOR2_X1 U124 ( .A(input0[5]), .B(output0[37]), .Z(output0[5]) );
  XOR2_X1 U125 ( .A(input0[6]), .B(output0[38]), .Z(output0[6]) );
  XOR2_X1 U126 ( .A(input0[7]), .B(output0[39]), .Z(output0[7]) );
  XOR2_X1 U127 ( .A(input0[8]), .B(output0[40]), .Z(output0[8]) );
  XOR2_X1 U128 ( .A(input0[9]), .B(output0[41]), .Z(output0[9]) );
endmodule


module MyDFFs_0 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_0 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_0 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module MyDFFs_259 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_259 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_259 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module MyDFFs_258 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_258 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_258 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module MyDFFs_257 ( D, CK, Q );
  input D, CK;
  output Q;


  DFF_X1 FF ( .D(D), .CK(CK), .Q(Q), .QN() );
endmodule


module MyDFF_257 ( D, CK, Q, QN );
  input D, CK;
  output Q, QN;


  MyDFFs_257 FF ( .D(D), .CK(CK), .Q(Q) );
  INV_X1 U1 ( .A(Q), .ZN(QN) );
endmodule


module counter_size4 ( clk, en, reset, q );
  output [3:0] q;
  input clk, en, reset;
  wire   n27, n26, n1, n25, n24, n2, n3, n4, n5, n6, n7, n8;

  MyDFF_0 count_reg_0_ ( .D(n27), .CK(clk), .Q(q[0]), .QN() );
  MyDFF_259 count_reg_1_ ( .D(n26), .CK(clk), .Q(q[1]), .QN(n1) );
  MyDFF_258 count_reg_2_ ( .D(n25), .CK(clk), .Q(q[2]), .QN() );
  MyDFF_257 count_reg_3_ ( .D(n24), .CK(clk), .Q(q[3]), .QN() );
  NAND2_X1 U1 ( .A1(en), .A2(q[0]), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n6), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n4), .A2(q[2]), .ZN(n2) );
  XOR2_X1 U4 ( .A(q[3]), .B(n2), .Z(n3) );
  NOR2_X1 U5 ( .A1(reset), .A2(n3), .ZN(n24) );
  XNOR2_X1 U6 ( .A(q[2]), .B(n4), .ZN(n5) );
  NOR2_X1 U7 ( .A1(reset), .A2(n5), .ZN(n25) );
  XOR2_X1 U8 ( .A(q[1]), .B(n6), .Z(n7) );
  NOR2_X1 U9 ( .A1(reset), .A2(n7), .ZN(n26) );
  XNOR2_X1 U10 ( .A(q[0]), .B(en), .ZN(n8) );
  NOR2_X1 U11 ( .A1(reset), .A2(n8), .ZN(n27) );
endmodule


module AES ( clk, start, port_in, port_out, done );
  input [7:0] port_in;
  output [7:0] port_out;
  input clk, start;
  output done;
  wire   start_done, n286, n287, notdone, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854;
  wire   [127:0] RoundOutput;
  wire   [127:8] state_shifted;
  wire   [127:120] RoundInput;
  wire   [127:0] ShiftRowsInput;
  wire   [119:0] SubBytesInput;
  wire   [127:0] MixColumnsInput;
  wire   [127:0] MixColumnsOutput;
  wire   [127:0] KeyExpansionOutput;
  wire   [127:8] key_shifted;
  wire   [127:120] RoundKey;
  wire   [5:0] Rcon;
  wire   [3:0] RoundCounter;

  reg_SDE_size128_0 RoundReg ( .clk(clk), .D0(RoundOutput), .D1({state_shifted, 
        port_in}), .sel(start_done), .Q({RoundInput, state_shifted}) );
  SubBytes SubBytesIns ( .input0({port_out, SubBytesInput}), .output0(
        ShiftRowsInput) );
  ShiftRows ShiftRowsIns ( .input0(ShiftRowsInput), .output0(MixColumnsInput)
         );
  MixColumns MixColumnsIns ( .input0(MixColumnsInput), .output0(
        MixColumnsOutput) );
  reg_SDE_size128_1 KeyReg ( .clk(clk), .D0(KeyExpansionOutput), .D1({
        key_shifted, RoundInput}), .sel(start_done), .Q({RoundKey, key_shifted}) );
  KeyExpansion KeyExpansionIns ( .input0({RoundKey, key_shifted}), .Rcon({n286, 
        n287, Rcon}), .output0(KeyExpansionOutput) );
  counter_size4 RoundCounterIns ( .clk(clk), .en(notdone), .reset(start), .q(
        RoundCounter) );
  INV_X8 U1092 ( .A(n845), .ZN(n579) );
  OR2_X1 U1093 ( .A1(start), .A2(done), .ZN(start_done) );
  INV_X1 U1094 ( .A(n579), .ZN(n574) );
  INV_X1 U1095 ( .A(n579), .ZN(n576) );
  INV_X1 U1096 ( .A(n579), .ZN(n575) );
  INV_X1 U1097 ( .A(n579), .ZN(n577) );
  INV_X1 U1098 ( .A(n579), .ZN(n578) );
  NAND2_X1 U1099 ( .A1(RoundCounter[0]), .A2(n587), .ZN(n845) );
  NOR2_X1 U1100 ( .A1(n852), .A2(n580), .ZN(n587) );
  INV_X1 U1101 ( .A(notdone), .ZN(done) );
  NAND2_X1 U1102 ( .A1(n854), .A2(n853), .ZN(notdone) );
  INV_X1 U1103 ( .A(RoundCounter[3]), .ZN(n852) );
  NOR2_X1 U1104 ( .A1(RoundCounter[2]), .A2(n584), .ZN(n854) );
  INV_X1 U1105 ( .A(RoundCounter[1]), .ZN(n584) );
  INV_X1 U1106 ( .A(RoundCounter[2]), .ZN(n851) );
  NOR2_X1 U1107 ( .A1(RoundCounter[0]), .A2(n852), .ZN(n853) );
  NAND2_X1 U1108 ( .A1(n851), .A2(n584), .ZN(n580) );
  NOR2_X1 U1109 ( .A1(RoundCounter[0]), .A2(n580), .ZN(Rcon[0]) );
  NOR2_X1 U1110 ( .A1(RoundCounter[0]), .A2(RoundCounter[3]), .ZN(n849) );
  NOR2_X1 U1111 ( .A1(n849), .A2(n580), .ZN(Rcon[1]) );
  NAND2_X1 U1112 ( .A1(n854), .A2(n849), .ZN(n581) );
  NAND2_X1 U1113 ( .A1(n578), .A2(n581), .ZN(Rcon[2]) );
  NAND2_X1 U1114 ( .A1(RoundCounter[0]), .A2(n852), .ZN(n589) );
  NOR2_X1 U1115 ( .A1(n584), .A2(n589), .ZN(n848) );
  NAND2_X1 U1116 ( .A1(n848), .A2(n851), .ZN(n583) );
  NAND2_X1 U1117 ( .A1(RoundCounter[3]), .A2(Rcon[0]), .ZN(n582) );
  NAND2_X1 U1118 ( .A1(n583), .A2(n582), .ZN(Rcon[3]) );
  INV_X1 U1119 ( .A(n849), .ZN(n585) );
  NAND2_X1 U1120 ( .A1(RoundCounter[2]), .A2(n584), .ZN(n588) );
  NOR2_X1 U1121 ( .A1(n585), .A2(n588), .ZN(n586) );
  OR2_X1 U1122 ( .A1(n587), .A2(n586), .ZN(Rcon[4]) );
  OR2_X1 U1123 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U1124 ( .A1(n578), .A2(n590), .ZN(Rcon[5]) );
  NAND2_X1 U1125 ( .A1(MixColumnsOutput[0]), .A2(n578), .ZN(n592) );
  NAND2_X1 U1126 ( .A1(n579), .A2(MixColumnsInput[0]), .ZN(n591) );
  NAND2_X1 U1127 ( .A1(n592), .A2(n591), .ZN(RoundOutput[0]) );
  NAND2_X1 U1128 ( .A1(MixColumnsOutput[100]), .A2(n578), .ZN(n594) );
  NAND2_X1 U1129 ( .A1(n579), .A2(MixColumnsInput[100]), .ZN(n593) );
  NAND2_X1 U1130 ( .A1(n594), .A2(n593), .ZN(RoundOutput[100]) );
  NAND2_X1 U1131 ( .A1(MixColumnsOutput[101]), .A2(n578), .ZN(n596) );
  NAND2_X1 U1132 ( .A1(n579), .A2(MixColumnsInput[101]), .ZN(n595) );
  NAND2_X1 U1133 ( .A1(n596), .A2(n595), .ZN(RoundOutput[101]) );
  NAND2_X1 U1134 ( .A1(MixColumnsOutput[102]), .A2(n578), .ZN(n598) );
  NAND2_X1 U1135 ( .A1(n579), .A2(MixColumnsInput[102]), .ZN(n597) );
  NAND2_X1 U1136 ( .A1(n598), .A2(n597), .ZN(RoundOutput[102]) );
  NAND2_X1 U1137 ( .A1(MixColumnsOutput[103]), .A2(n578), .ZN(n600) );
  NAND2_X1 U1138 ( .A1(n579), .A2(MixColumnsInput[103]), .ZN(n599) );
  NAND2_X1 U1139 ( .A1(n600), .A2(n599), .ZN(RoundOutput[103]) );
  NAND2_X1 U1140 ( .A1(MixColumnsOutput[104]), .A2(n578), .ZN(n602) );
  NAND2_X1 U1141 ( .A1(n579), .A2(MixColumnsInput[104]), .ZN(n601) );
  NAND2_X1 U1142 ( .A1(n602), .A2(n601), .ZN(RoundOutput[104]) );
  NAND2_X1 U1143 ( .A1(MixColumnsOutput[105]), .A2(n578), .ZN(n604) );
  NAND2_X1 U1144 ( .A1(n579), .A2(MixColumnsInput[105]), .ZN(n603) );
  NAND2_X1 U1145 ( .A1(n604), .A2(n603), .ZN(RoundOutput[105]) );
  NAND2_X1 U1146 ( .A1(MixColumnsOutput[106]), .A2(n578), .ZN(n606) );
  NAND2_X1 U1147 ( .A1(n579), .A2(MixColumnsInput[106]), .ZN(n605) );
  NAND2_X1 U1148 ( .A1(n606), .A2(n605), .ZN(RoundOutput[106]) );
  NAND2_X1 U1149 ( .A1(MixColumnsOutput[107]), .A2(n577), .ZN(n608) );
  NAND2_X1 U1150 ( .A1(n579), .A2(MixColumnsInput[107]), .ZN(n607) );
  NAND2_X1 U1151 ( .A1(n608), .A2(n607), .ZN(RoundOutput[107]) );
  NAND2_X1 U1152 ( .A1(MixColumnsOutput[108]), .A2(n577), .ZN(n610) );
  NAND2_X1 U1153 ( .A1(n579), .A2(MixColumnsInput[108]), .ZN(n609) );
  NAND2_X1 U1154 ( .A1(n610), .A2(n609), .ZN(RoundOutput[108]) );
  NAND2_X1 U1155 ( .A1(MixColumnsOutput[109]), .A2(n577), .ZN(n612) );
  NAND2_X1 U1156 ( .A1(n579), .A2(MixColumnsInput[109]), .ZN(n611) );
  NAND2_X1 U1157 ( .A1(n612), .A2(n611), .ZN(RoundOutput[109]) );
  NAND2_X1 U1158 ( .A1(MixColumnsOutput[10]), .A2(n577), .ZN(n614) );
  NAND2_X1 U1159 ( .A1(n579), .A2(MixColumnsInput[10]), .ZN(n613) );
  NAND2_X1 U1160 ( .A1(n614), .A2(n613), .ZN(RoundOutput[10]) );
  NAND2_X1 U1161 ( .A1(MixColumnsOutput[110]), .A2(n577), .ZN(n616) );
  NAND2_X1 U1162 ( .A1(n579), .A2(MixColumnsInput[110]), .ZN(n615) );
  NAND2_X1 U1163 ( .A1(n616), .A2(n615), .ZN(RoundOutput[110]) );
  NAND2_X1 U1164 ( .A1(MixColumnsOutput[111]), .A2(n577), .ZN(n618) );
  NAND2_X1 U1165 ( .A1(n579), .A2(MixColumnsInput[111]), .ZN(n617) );
  NAND2_X1 U1166 ( .A1(n618), .A2(n617), .ZN(RoundOutput[111]) );
  NAND2_X1 U1167 ( .A1(MixColumnsOutput[112]), .A2(n577), .ZN(n620) );
  NAND2_X1 U1168 ( .A1(n579), .A2(MixColumnsInput[112]), .ZN(n619) );
  NAND2_X1 U1169 ( .A1(n620), .A2(n619), .ZN(RoundOutput[112]) );
  NAND2_X1 U1170 ( .A1(MixColumnsOutput[113]), .A2(n577), .ZN(n622) );
  NAND2_X1 U1171 ( .A1(n579), .A2(MixColumnsInput[113]), .ZN(n621) );
  NAND2_X1 U1172 ( .A1(n622), .A2(n621), .ZN(RoundOutput[113]) );
  NAND2_X1 U1173 ( .A1(MixColumnsOutput[114]), .A2(n577), .ZN(n624) );
  NAND2_X1 U1174 ( .A1(n579), .A2(MixColumnsInput[114]), .ZN(n623) );
  NAND2_X1 U1175 ( .A1(n624), .A2(n623), .ZN(RoundOutput[114]) );
  NAND2_X1 U1176 ( .A1(MixColumnsOutput[115]), .A2(n577), .ZN(n626) );
  NAND2_X1 U1177 ( .A1(n579), .A2(MixColumnsInput[115]), .ZN(n625) );
  NAND2_X1 U1178 ( .A1(n626), .A2(n625), .ZN(RoundOutput[115]) );
  NAND2_X1 U1179 ( .A1(MixColumnsOutput[116]), .A2(n577), .ZN(n628) );
  NAND2_X1 U1180 ( .A1(n579), .A2(MixColumnsInput[116]), .ZN(n627) );
  NAND2_X1 U1181 ( .A1(n628), .A2(n627), .ZN(RoundOutput[116]) );
  NAND2_X1 U1182 ( .A1(MixColumnsOutput[117]), .A2(n577), .ZN(n630) );
  NAND2_X1 U1183 ( .A1(n579), .A2(MixColumnsInput[117]), .ZN(n629) );
  NAND2_X1 U1184 ( .A1(n630), .A2(n629), .ZN(RoundOutput[117]) );
  NAND2_X1 U1185 ( .A1(MixColumnsOutput[118]), .A2(n576), .ZN(n632) );
  NAND2_X1 U1186 ( .A1(n579), .A2(MixColumnsInput[118]), .ZN(n631) );
  NAND2_X1 U1187 ( .A1(n632), .A2(n631), .ZN(RoundOutput[118]) );
  NAND2_X1 U1188 ( .A1(MixColumnsOutput[119]), .A2(n576), .ZN(n634) );
  NAND2_X1 U1189 ( .A1(n579), .A2(MixColumnsInput[119]), .ZN(n633) );
  NAND2_X1 U1190 ( .A1(n634), .A2(n633), .ZN(RoundOutput[119]) );
  NAND2_X1 U1191 ( .A1(MixColumnsOutput[11]), .A2(n576), .ZN(n636) );
  NAND2_X1 U1192 ( .A1(n579), .A2(MixColumnsInput[11]), .ZN(n635) );
  NAND2_X1 U1193 ( .A1(n636), .A2(n635), .ZN(RoundOutput[11]) );
  NAND2_X1 U1194 ( .A1(MixColumnsOutput[120]), .A2(n576), .ZN(n638) );
  NAND2_X1 U1195 ( .A1(n579), .A2(MixColumnsInput[120]), .ZN(n637) );
  NAND2_X1 U1196 ( .A1(n638), .A2(n637), .ZN(RoundOutput[120]) );
  NAND2_X1 U1197 ( .A1(MixColumnsOutput[121]), .A2(n576), .ZN(n640) );
  NAND2_X1 U1198 ( .A1(n579), .A2(MixColumnsInput[121]), .ZN(n639) );
  NAND2_X1 U1199 ( .A1(n640), .A2(n639), .ZN(RoundOutput[121]) );
  NAND2_X1 U1200 ( .A1(MixColumnsOutput[122]), .A2(n576), .ZN(n642) );
  NAND2_X1 U1201 ( .A1(n579), .A2(MixColumnsInput[122]), .ZN(n641) );
  NAND2_X1 U1202 ( .A1(n642), .A2(n641), .ZN(RoundOutput[122]) );
  NAND2_X1 U1203 ( .A1(MixColumnsOutput[123]), .A2(n576), .ZN(n644) );
  NAND2_X1 U1204 ( .A1(n579), .A2(MixColumnsInput[123]), .ZN(n643) );
  NAND2_X1 U1205 ( .A1(n644), .A2(n643), .ZN(RoundOutput[123]) );
  NAND2_X1 U1206 ( .A1(MixColumnsOutput[124]), .A2(n576), .ZN(n646) );
  NAND2_X1 U1207 ( .A1(n579), .A2(MixColumnsInput[124]), .ZN(n645) );
  NAND2_X1 U1208 ( .A1(n646), .A2(n645), .ZN(RoundOutput[124]) );
  NAND2_X1 U1209 ( .A1(MixColumnsOutput[125]), .A2(n576), .ZN(n648) );
  NAND2_X1 U1210 ( .A1(n579), .A2(MixColumnsInput[125]), .ZN(n647) );
  NAND2_X1 U1211 ( .A1(n648), .A2(n647), .ZN(RoundOutput[125]) );
  NAND2_X1 U1212 ( .A1(MixColumnsOutput[126]), .A2(n576), .ZN(n650) );
  NAND2_X1 U1213 ( .A1(n579), .A2(MixColumnsInput[126]), .ZN(n649) );
  NAND2_X1 U1214 ( .A1(n650), .A2(n649), .ZN(RoundOutput[126]) );
  NAND2_X1 U1215 ( .A1(MixColumnsOutput[127]), .A2(n576), .ZN(n652) );
  NAND2_X1 U1216 ( .A1(n579), .A2(MixColumnsInput[127]), .ZN(n651) );
  NAND2_X1 U1217 ( .A1(n652), .A2(n651), .ZN(RoundOutput[127]) );
  NAND2_X1 U1218 ( .A1(MixColumnsOutput[12]), .A2(n576), .ZN(n654) );
  NAND2_X1 U1219 ( .A1(n579), .A2(MixColumnsInput[12]), .ZN(n653) );
  NAND2_X1 U1220 ( .A1(n654), .A2(n653), .ZN(RoundOutput[12]) );
  NAND2_X1 U1221 ( .A1(MixColumnsOutput[13]), .A2(n575), .ZN(n656) );
  NAND2_X1 U1222 ( .A1(n579), .A2(MixColumnsInput[13]), .ZN(n655) );
  NAND2_X1 U1223 ( .A1(n656), .A2(n655), .ZN(RoundOutput[13]) );
  NAND2_X1 U1224 ( .A1(MixColumnsOutput[14]), .A2(n575), .ZN(n658) );
  NAND2_X1 U1225 ( .A1(n579), .A2(MixColumnsInput[14]), .ZN(n657) );
  NAND2_X1 U1226 ( .A1(n658), .A2(n657), .ZN(RoundOutput[14]) );
  NAND2_X1 U1227 ( .A1(MixColumnsOutput[15]), .A2(n575), .ZN(n660) );
  NAND2_X1 U1228 ( .A1(n579), .A2(MixColumnsInput[15]), .ZN(n659) );
  NAND2_X1 U1229 ( .A1(n660), .A2(n659), .ZN(RoundOutput[15]) );
  NAND2_X1 U1230 ( .A1(MixColumnsOutput[16]), .A2(n575), .ZN(n662) );
  NAND2_X1 U1231 ( .A1(n579), .A2(MixColumnsInput[16]), .ZN(n661) );
  NAND2_X1 U1232 ( .A1(n662), .A2(n661), .ZN(RoundOutput[16]) );
  NAND2_X1 U1233 ( .A1(MixColumnsOutput[17]), .A2(n575), .ZN(n664) );
  NAND2_X1 U1234 ( .A1(n579), .A2(MixColumnsInput[17]), .ZN(n663) );
  NAND2_X1 U1235 ( .A1(n664), .A2(n663), .ZN(RoundOutput[17]) );
  NAND2_X1 U1236 ( .A1(MixColumnsOutput[18]), .A2(n575), .ZN(n666) );
  NAND2_X1 U1237 ( .A1(n579), .A2(MixColumnsInput[18]), .ZN(n665) );
  NAND2_X1 U1238 ( .A1(n666), .A2(n665), .ZN(RoundOutput[18]) );
  NAND2_X1 U1239 ( .A1(MixColumnsOutput[19]), .A2(n575), .ZN(n668) );
  NAND2_X1 U1240 ( .A1(n579), .A2(MixColumnsInput[19]), .ZN(n667) );
  NAND2_X1 U1241 ( .A1(n668), .A2(n667), .ZN(RoundOutput[19]) );
  NAND2_X1 U1242 ( .A1(MixColumnsOutput[1]), .A2(n575), .ZN(n670) );
  NAND2_X1 U1243 ( .A1(n579), .A2(MixColumnsInput[1]), .ZN(n669) );
  NAND2_X1 U1244 ( .A1(n670), .A2(n669), .ZN(RoundOutput[1]) );
  NAND2_X1 U1245 ( .A1(MixColumnsOutput[20]), .A2(n575), .ZN(n672) );
  NAND2_X1 U1246 ( .A1(n579), .A2(MixColumnsInput[20]), .ZN(n671) );
  NAND2_X1 U1247 ( .A1(n672), .A2(n671), .ZN(RoundOutput[20]) );
  NAND2_X1 U1248 ( .A1(MixColumnsOutput[21]), .A2(n575), .ZN(n674) );
  NAND2_X1 U1249 ( .A1(n579), .A2(MixColumnsInput[21]), .ZN(n673) );
  NAND2_X1 U1250 ( .A1(n674), .A2(n673), .ZN(RoundOutput[21]) );
  NAND2_X1 U1251 ( .A1(MixColumnsOutput[22]), .A2(n575), .ZN(n676) );
  NAND2_X1 U1252 ( .A1(n579), .A2(MixColumnsInput[22]), .ZN(n675) );
  NAND2_X1 U1253 ( .A1(n676), .A2(n675), .ZN(RoundOutput[22]) );
  NAND2_X1 U1254 ( .A1(MixColumnsOutput[23]), .A2(n575), .ZN(n678) );
  NAND2_X1 U1255 ( .A1(n579), .A2(MixColumnsInput[23]), .ZN(n677) );
  NAND2_X1 U1256 ( .A1(n678), .A2(n677), .ZN(RoundOutput[23]) );
  NAND2_X1 U1257 ( .A1(MixColumnsOutput[24]), .A2(n574), .ZN(n680) );
  NAND2_X1 U1258 ( .A1(n579), .A2(MixColumnsInput[24]), .ZN(n679) );
  NAND2_X1 U1259 ( .A1(n680), .A2(n679), .ZN(RoundOutput[24]) );
  NAND2_X1 U1260 ( .A1(MixColumnsOutput[25]), .A2(n574), .ZN(n682) );
  NAND2_X1 U1261 ( .A1(n579), .A2(MixColumnsInput[25]), .ZN(n681) );
  NAND2_X1 U1262 ( .A1(n682), .A2(n681), .ZN(RoundOutput[25]) );
  NAND2_X1 U1263 ( .A1(MixColumnsOutput[26]), .A2(n574), .ZN(n684) );
  NAND2_X1 U1264 ( .A1(n579), .A2(MixColumnsInput[26]), .ZN(n683) );
  NAND2_X1 U1265 ( .A1(n684), .A2(n683), .ZN(RoundOutput[26]) );
  NAND2_X1 U1266 ( .A1(MixColumnsOutput[27]), .A2(n574), .ZN(n686) );
  NAND2_X1 U1267 ( .A1(n579), .A2(MixColumnsInput[27]), .ZN(n685) );
  NAND2_X1 U1268 ( .A1(n686), .A2(n685), .ZN(RoundOutput[27]) );
  NAND2_X1 U1269 ( .A1(MixColumnsOutput[28]), .A2(n574), .ZN(n688) );
  NAND2_X1 U1270 ( .A1(n579), .A2(MixColumnsInput[28]), .ZN(n687) );
  NAND2_X1 U1271 ( .A1(n688), .A2(n687), .ZN(RoundOutput[28]) );
  NAND2_X1 U1272 ( .A1(MixColumnsOutput[29]), .A2(n574), .ZN(n690) );
  NAND2_X1 U1273 ( .A1(n579), .A2(MixColumnsInput[29]), .ZN(n689) );
  NAND2_X1 U1274 ( .A1(n690), .A2(n689), .ZN(RoundOutput[29]) );
  NAND2_X1 U1275 ( .A1(MixColumnsOutput[2]), .A2(n574), .ZN(n692) );
  NAND2_X1 U1276 ( .A1(n579), .A2(MixColumnsInput[2]), .ZN(n691) );
  NAND2_X1 U1277 ( .A1(n692), .A2(n691), .ZN(RoundOutput[2]) );
  NAND2_X1 U1278 ( .A1(MixColumnsOutput[30]), .A2(n574), .ZN(n694) );
  NAND2_X1 U1279 ( .A1(n579), .A2(MixColumnsInput[30]), .ZN(n693) );
  NAND2_X1 U1280 ( .A1(n694), .A2(n693), .ZN(RoundOutput[30]) );
  NAND2_X1 U1281 ( .A1(MixColumnsOutput[31]), .A2(n574), .ZN(n696) );
  NAND2_X1 U1282 ( .A1(n579), .A2(MixColumnsInput[31]), .ZN(n695) );
  NAND2_X1 U1283 ( .A1(n696), .A2(n695), .ZN(RoundOutput[31]) );
  NAND2_X1 U1284 ( .A1(MixColumnsOutput[32]), .A2(n574), .ZN(n698) );
  NAND2_X1 U1285 ( .A1(n579), .A2(MixColumnsInput[32]), .ZN(n697) );
  NAND2_X1 U1286 ( .A1(n698), .A2(n697), .ZN(RoundOutput[32]) );
  NAND2_X1 U1287 ( .A1(MixColumnsOutput[33]), .A2(n574), .ZN(n700) );
  NAND2_X1 U1288 ( .A1(n579), .A2(MixColumnsInput[33]), .ZN(n699) );
  NAND2_X1 U1289 ( .A1(n700), .A2(n699), .ZN(RoundOutput[33]) );
  NAND2_X1 U1290 ( .A1(MixColumnsOutput[34]), .A2(n574), .ZN(n702) );
  NAND2_X1 U1291 ( .A1(n579), .A2(MixColumnsInput[34]), .ZN(n701) );
  NAND2_X1 U1292 ( .A1(n702), .A2(n701), .ZN(RoundOutput[34]) );
  NAND2_X1 U1293 ( .A1(MixColumnsOutput[35]), .A2(n845), .ZN(n704) );
  NAND2_X1 U1294 ( .A1(n579), .A2(MixColumnsInput[35]), .ZN(n703) );
  NAND2_X1 U1295 ( .A1(n704), .A2(n703), .ZN(RoundOutput[35]) );
  NAND2_X1 U1296 ( .A1(MixColumnsOutput[36]), .A2(n578), .ZN(n706) );
  NAND2_X1 U1297 ( .A1(n579), .A2(MixColumnsInput[36]), .ZN(n705) );
  NAND2_X1 U1298 ( .A1(n706), .A2(n705), .ZN(RoundOutput[36]) );
  NAND2_X1 U1299 ( .A1(MixColumnsOutput[37]), .A2(n578), .ZN(n708) );
  NAND2_X1 U1300 ( .A1(n579), .A2(MixColumnsInput[37]), .ZN(n707) );
  NAND2_X1 U1301 ( .A1(n708), .A2(n707), .ZN(RoundOutput[37]) );
  NAND2_X1 U1302 ( .A1(MixColumnsOutput[38]), .A2(n845), .ZN(n710) );
  NAND2_X1 U1303 ( .A1(n579), .A2(MixColumnsInput[38]), .ZN(n709) );
  NAND2_X1 U1304 ( .A1(n710), .A2(n709), .ZN(RoundOutput[38]) );
  NAND2_X1 U1305 ( .A1(MixColumnsOutput[39]), .A2(n845), .ZN(n712) );
  NAND2_X1 U1306 ( .A1(n579), .A2(MixColumnsInput[39]), .ZN(n711) );
  NAND2_X1 U1307 ( .A1(n712), .A2(n711), .ZN(RoundOutput[39]) );
  NAND2_X1 U1308 ( .A1(MixColumnsOutput[3]), .A2(n578), .ZN(n714) );
  NAND2_X1 U1309 ( .A1(n579), .A2(MixColumnsInput[3]), .ZN(n713) );
  NAND2_X1 U1310 ( .A1(n714), .A2(n713), .ZN(RoundOutput[3]) );
  NAND2_X1 U1311 ( .A1(MixColumnsOutput[40]), .A2(n845), .ZN(n716) );
  NAND2_X1 U1312 ( .A1(n579), .A2(MixColumnsInput[40]), .ZN(n715) );
  NAND2_X1 U1313 ( .A1(n716), .A2(n715), .ZN(RoundOutput[40]) );
  NAND2_X1 U1314 ( .A1(MixColumnsOutput[41]), .A2(n845), .ZN(n718) );
  NAND2_X1 U1315 ( .A1(n579), .A2(MixColumnsInput[41]), .ZN(n717) );
  NAND2_X1 U1316 ( .A1(n718), .A2(n717), .ZN(RoundOutput[41]) );
  NAND2_X1 U1317 ( .A1(MixColumnsOutput[42]), .A2(n845), .ZN(n720) );
  NAND2_X1 U1318 ( .A1(n579), .A2(MixColumnsInput[42]), .ZN(n719) );
  NAND2_X1 U1319 ( .A1(n720), .A2(n719), .ZN(RoundOutput[42]) );
  NAND2_X1 U1320 ( .A1(MixColumnsOutput[43]), .A2(n845), .ZN(n722) );
  NAND2_X1 U1321 ( .A1(n579), .A2(MixColumnsInput[43]), .ZN(n721) );
  NAND2_X1 U1322 ( .A1(n722), .A2(n721), .ZN(RoundOutput[43]) );
  NAND2_X1 U1323 ( .A1(MixColumnsOutput[44]), .A2(n578), .ZN(n724) );
  NAND2_X1 U1324 ( .A1(n579), .A2(MixColumnsInput[44]), .ZN(n723) );
  NAND2_X1 U1325 ( .A1(n724), .A2(n723), .ZN(RoundOutput[44]) );
  NAND2_X1 U1326 ( .A1(MixColumnsOutput[45]), .A2(n578), .ZN(n726) );
  NAND2_X1 U1327 ( .A1(n579), .A2(MixColumnsInput[45]), .ZN(n725) );
  NAND2_X1 U1328 ( .A1(n726), .A2(n725), .ZN(RoundOutput[45]) );
  NAND2_X1 U1329 ( .A1(MixColumnsOutput[46]), .A2(n578), .ZN(n728) );
  NAND2_X1 U1330 ( .A1(n579), .A2(MixColumnsInput[46]), .ZN(n727) );
  NAND2_X1 U1331 ( .A1(n728), .A2(n727), .ZN(RoundOutput[46]) );
  NAND2_X1 U1332 ( .A1(MixColumnsOutput[47]), .A2(n578), .ZN(n730) );
  NAND2_X1 U1333 ( .A1(n579), .A2(MixColumnsInput[47]), .ZN(n729) );
  NAND2_X1 U1334 ( .A1(n730), .A2(n729), .ZN(RoundOutput[47]) );
  NAND2_X1 U1335 ( .A1(MixColumnsOutput[48]), .A2(n578), .ZN(n732) );
  NAND2_X1 U1336 ( .A1(n579), .A2(MixColumnsInput[48]), .ZN(n731) );
  NAND2_X1 U1337 ( .A1(n732), .A2(n731), .ZN(RoundOutput[48]) );
  NAND2_X1 U1338 ( .A1(MixColumnsOutput[49]), .A2(n574), .ZN(n734) );
  NAND2_X1 U1339 ( .A1(n579), .A2(MixColumnsInput[49]), .ZN(n733) );
  NAND2_X1 U1340 ( .A1(n734), .A2(n733), .ZN(RoundOutput[49]) );
  NAND2_X1 U1341 ( .A1(MixColumnsOutput[4]), .A2(n574), .ZN(n736) );
  NAND2_X1 U1342 ( .A1(n579), .A2(MixColumnsInput[4]), .ZN(n735) );
  NAND2_X1 U1343 ( .A1(n736), .A2(n735), .ZN(RoundOutput[4]) );
  NAND2_X1 U1344 ( .A1(MixColumnsOutput[50]), .A2(n576), .ZN(n738) );
  NAND2_X1 U1345 ( .A1(n579), .A2(MixColumnsInput[50]), .ZN(n737) );
  NAND2_X1 U1346 ( .A1(n738), .A2(n737), .ZN(RoundOutput[50]) );
  NAND2_X1 U1347 ( .A1(MixColumnsOutput[51]), .A2(n575), .ZN(n740) );
  NAND2_X1 U1348 ( .A1(n579), .A2(MixColumnsInput[51]), .ZN(n739) );
  NAND2_X1 U1349 ( .A1(n740), .A2(n739), .ZN(RoundOutput[51]) );
  NAND2_X1 U1350 ( .A1(MixColumnsOutput[52]), .A2(n576), .ZN(n742) );
  NAND2_X1 U1351 ( .A1(n579), .A2(MixColumnsInput[52]), .ZN(n741) );
  NAND2_X1 U1352 ( .A1(n742), .A2(n741), .ZN(RoundOutput[52]) );
  NAND2_X1 U1353 ( .A1(MixColumnsOutput[53]), .A2(n578), .ZN(n744) );
  NAND2_X1 U1354 ( .A1(n579), .A2(MixColumnsInput[53]), .ZN(n743) );
  NAND2_X1 U1355 ( .A1(n744), .A2(n743), .ZN(RoundOutput[53]) );
  NAND2_X1 U1356 ( .A1(MixColumnsOutput[54]), .A2(n845), .ZN(n746) );
  NAND2_X1 U1357 ( .A1(n579), .A2(MixColumnsInput[54]), .ZN(n745) );
  NAND2_X1 U1358 ( .A1(n746), .A2(n745), .ZN(RoundOutput[54]) );
  NAND2_X1 U1359 ( .A1(MixColumnsOutput[55]), .A2(n575), .ZN(n748) );
  NAND2_X1 U1360 ( .A1(n579), .A2(MixColumnsInput[55]), .ZN(n747) );
  NAND2_X1 U1361 ( .A1(n748), .A2(n747), .ZN(RoundOutput[55]) );
  NAND2_X1 U1362 ( .A1(MixColumnsOutput[56]), .A2(n845), .ZN(n750) );
  NAND2_X1 U1363 ( .A1(n579), .A2(MixColumnsInput[56]), .ZN(n749) );
  NAND2_X1 U1364 ( .A1(n750), .A2(n749), .ZN(RoundOutput[56]) );
  NAND2_X1 U1365 ( .A1(MixColumnsOutput[57]), .A2(n574), .ZN(n752) );
  NAND2_X1 U1366 ( .A1(n579), .A2(MixColumnsInput[57]), .ZN(n751) );
  NAND2_X1 U1367 ( .A1(n752), .A2(n751), .ZN(RoundOutput[57]) );
  NAND2_X1 U1368 ( .A1(MixColumnsOutput[58]), .A2(n576), .ZN(n754) );
  NAND2_X1 U1369 ( .A1(n579), .A2(MixColumnsInput[58]), .ZN(n753) );
  NAND2_X1 U1370 ( .A1(n754), .A2(n753), .ZN(RoundOutput[58]) );
  NAND2_X1 U1371 ( .A1(MixColumnsOutput[59]), .A2(n577), .ZN(n756) );
  NAND2_X1 U1372 ( .A1(n579), .A2(MixColumnsInput[59]), .ZN(n755) );
  NAND2_X1 U1373 ( .A1(n756), .A2(n755), .ZN(RoundOutput[59]) );
  NAND2_X1 U1374 ( .A1(MixColumnsOutput[5]), .A2(n575), .ZN(n758) );
  NAND2_X1 U1375 ( .A1(n579), .A2(MixColumnsInput[5]), .ZN(n757) );
  NAND2_X1 U1376 ( .A1(n758), .A2(n757), .ZN(RoundOutput[5]) );
  NAND2_X1 U1377 ( .A1(MixColumnsOutput[60]), .A2(n577), .ZN(n760) );
  NAND2_X1 U1378 ( .A1(n579), .A2(MixColumnsInput[60]), .ZN(n759) );
  NAND2_X1 U1379 ( .A1(n760), .A2(n759), .ZN(RoundOutput[60]) );
  NAND2_X1 U1380 ( .A1(MixColumnsOutput[61]), .A2(n845), .ZN(n762) );
  NAND2_X1 U1381 ( .A1(n579), .A2(MixColumnsInput[61]), .ZN(n761) );
  NAND2_X1 U1382 ( .A1(n762), .A2(n761), .ZN(RoundOutput[61]) );
  NAND2_X1 U1383 ( .A1(MixColumnsOutput[62]), .A2(n845), .ZN(n764) );
  NAND2_X1 U1384 ( .A1(n579), .A2(MixColumnsInput[62]), .ZN(n763) );
  NAND2_X1 U1385 ( .A1(n764), .A2(n763), .ZN(RoundOutput[62]) );
  NAND2_X1 U1386 ( .A1(MixColumnsOutput[63]), .A2(n574), .ZN(n766) );
  NAND2_X1 U1387 ( .A1(n579), .A2(MixColumnsInput[63]), .ZN(n765) );
  NAND2_X1 U1388 ( .A1(n766), .A2(n765), .ZN(RoundOutput[63]) );
  NAND2_X1 U1389 ( .A1(MixColumnsOutput[64]), .A2(n574), .ZN(n768) );
  NAND2_X1 U1390 ( .A1(n579), .A2(MixColumnsInput[64]), .ZN(n767) );
  NAND2_X1 U1391 ( .A1(n768), .A2(n767), .ZN(RoundOutput[64]) );
  NAND2_X1 U1392 ( .A1(MixColumnsOutput[65]), .A2(n576), .ZN(n770) );
  NAND2_X1 U1393 ( .A1(n579), .A2(MixColumnsInput[65]), .ZN(n769) );
  NAND2_X1 U1394 ( .A1(n770), .A2(n769), .ZN(RoundOutput[65]) );
  NAND2_X1 U1395 ( .A1(MixColumnsOutput[66]), .A2(n575), .ZN(n772) );
  NAND2_X1 U1396 ( .A1(n579), .A2(MixColumnsInput[66]), .ZN(n771) );
  NAND2_X1 U1397 ( .A1(n772), .A2(n771), .ZN(RoundOutput[66]) );
  NAND2_X1 U1398 ( .A1(MixColumnsOutput[67]), .A2(n577), .ZN(n774) );
  NAND2_X1 U1399 ( .A1(n579), .A2(MixColumnsInput[67]), .ZN(n773) );
  NAND2_X1 U1400 ( .A1(n774), .A2(n773), .ZN(RoundOutput[67]) );
  NAND2_X1 U1401 ( .A1(MixColumnsOutput[68]), .A2(n845), .ZN(n776) );
  NAND2_X1 U1402 ( .A1(n579), .A2(MixColumnsInput[68]), .ZN(n775) );
  NAND2_X1 U1403 ( .A1(n776), .A2(n775), .ZN(RoundOutput[68]) );
  NAND2_X1 U1404 ( .A1(MixColumnsOutput[69]), .A2(n845), .ZN(n778) );
  NAND2_X1 U1405 ( .A1(n579), .A2(MixColumnsInput[69]), .ZN(n777) );
  NAND2_X1 U1406 ( .A1(n778), .A2(n777), .ZN(RoundOutput[69]) );
  NAND2_X1 U1407 ( .A1(MixColumnsOutput[6]), .A2(n845), .ZN(n780) );
  NAND2_X1 U1408 ( .A1(n579), .A2(MixColumnsInput[6]), .ZN(n779) );
  NAND2_X1 U1409 ( .A1(n780), .A2(n779), .ZN(RoundOutput[6]) );
  NAND2_X1 U1410 ( .A1(MixColumnsOutput[70]), .A2(n574), .ZN(n782) );
  NAND2_X1 U1411 ( .A1(n579), .A2(MixColumnsInput[70]), .ZN(n781) );
  NAND2_X1 U1412 ( .A1(n782), .A2(n781), .ZN(RoundOutput[70]) );
  NAND2_X1 U1413 ( .A1(MixColumnsOutput[71]), .A2(n574), .ZN(n784) );
  NAND2_X1 U1414 ( .A1(n579), .A2(MixColumnsInput[71]), .ZN(n783) );
  NAND2_X1 U1415 ( .A1(n784), .A2(n783), .ZN(RoundOutput[71]) );
  NAND2_X1 U1416 ( .A1(MixColumnsOutput[72]), .A2(n574), .ZN(n786) );
  NAND2_X1 U1417 ( .A1(n579), .A2(MixColumnsInput[72]), .ZN(n785) );
  NAND2_X1 U1418 ( .A1(n786), .A2(n785), .ZN(RoundOutput[72]) );
  NAND2_X1 U1419 ( .A1(MixColumnsOutput[73]), .A2(n576), .ZN(n788) );
  NAND2_X1 U1420 ( .A1(n579), .A2(MixColumnsInput[73]), .ZN(n787) );
  NAND2_X1 U1421 ( .A1(n788), .A2(n787), .ZN(RoundOutput[73]) );
  NAND2_X1 U1422 ( .A1(MixColumnsOutput[74]), .A2(n575), .ZN(n790) );
  NAND2_X1 U1423 ( .A1(n579), .A2(MixColumnsInput[74]), .ZN(n789) );
  NAND2_X1 U1424 ( .A1(n790), .A2(n789), .ZN(RoundOutput[74]) );
  NAND2_X1 U1425 ( .A1(MixColumnsOutput[75]), .A2(n577), .ZN(n792) );
  NAND2_X1 U1426 ( .A1(n579), .A2(MixColumnsInput[75]), .ZN(n791) );
  NAND2_X1 U1427 ( .A1(n792), .A2(n791), .ZN(RoundOutput[75]) );
  NAND2_X1 U1428 ( .A1(MixColumnsOutput[76]), .A2(n576), .ZN(n794) );
  NAND2_X1 U1429 ( .A1(n579), .A2(MixColumnsInput[76]), .ZN(n793) );
  NAND2_X1 U1430 ( .A1(n794), .A2(n793), .ZN(RoundOutput[76]) );
  NAND2_X1 U1431 ( .A1(MixColumnsOutput[77]), .A2(n575), .ZN(n796) );
  NAND2_X1 U1432 ( .A1(n579), .A2(MixColumnsInput[77]), .ZN(n795) );
  NAND2_X1 U1433 ( .A1(n796), .A2(n795), .ZN(RoundOutput[77]) );
  NAND2_X1 U1434 ( .A1(MixColumnsOutput[78]), .A2(n845), .ZN(n798) );
  NAND2_X1 U1435 ( .A1(n579), .A2(MixColumnsInput[78]), .ZN(n797) );
  NAND2_X1 U1436 ( .A1(n798), .A2(n797), .ZN(RoundOutput[78]) );
  NAND2_X1 U1437 ( .A1(MixColumnsOutput[79]), .A2(n577), .ZN(n800) );
  NAND2_X1 U1438 ( .A1(n579), .A2(MixColumnsInput[79]), .ZN(n799) );
  NAND2_X1 U1439 ( .A1(n800), .A2(n799), .ZN(RoundOutput[79]) );
  NAND2_X1 U1440 ( .A1(MixColumnsOutput[7]), .A2(n576), .ZN(n802) );
  NAND2_X1 U1441 ( .A1(n579), .A2(MixColumnsInput[7]), .ZN(n801) );
  NAND2_X1 U1442 ( .A1(n802), .A2(n801), .ZN(RoundOutput[7]) );
  NAND2_X1 U1443 ( .A1(MixColumnsOutput[80]), .A2(n575), .ZN(n804) );
  NAND2_X1 U1444 ( .A1(n579), .A2(MixColumnsInput[80]), .ZN(n803) );
  NAND2_X1 U1445 ( .A1(n804), .A2(n803), .ZN(RoundOutput[80]) );
  NAND2_X1 U1446 ( .A1(MixColumnsOutput[81]), .A2(n577), .ZN(n806) );
  NAND2_X1 U1447 ( .A1(n579), .A2(MixColumnsInput[81]), .ZN(n805) );
  NAND2_X1 U1448 ( .A1(n806), .A2(n805), .ZN(RoundOutput[81]) );
  NAND2_X1 U1449 ( .A1(MixColumnsOutput[82]), .A2(n845), .ZN(n808) );
  NAND2_X1 U1450 ( .A1(n579), .A2(MixColumnsInput[82]), .ZN(n807) );
  NAND2_X1 U1451 ( .A1(n808), .A2(n807), .ZN(RoundOutput[82]) );
  NAND2_X1 U1452 ( .A1(MixColumnsOutput[83]), .A2(n576), .ZN(n810) );
  NAND2_X1 U1453 ( .A1(n579), .A2(MixColumnsInput[83]), .ZN(n809) );
  NAND2_X1 U1454 ( .A1(n810), .A2(n809), .ZN(RoundOutput[83]) );
  NAND2_X1 U1455 ( .A1(MixColumnsOutput[84]), .A2(n574), .ZN(n812) );
  NAND2_X1 U1456 ( .A1(n579), .A2(MixColumnsInput[84]), .ZN(n811) );
  NAND2_X1 U1457 ( .A1(n812), .A2(n811), .ZN(RoundOutput[84]) );
  NAND2_X1 U1458 ( .A1(MixColumnsOutput[85]), .A2(n576), .ZN(n814) );
  NAND2_X1 U1459 ( .A1(n579), .A2(MixColumnsInput[85]), .ZN(n813) );
  NAND2_X1 U1460 ( .A1(n814), .A2(n813), .ZN(RoundOutput[85]) );
  NAND2_X1 U1461 ( .A1(MixColumnsOutput[86]), .A2(n575), .ZN(n816) );
  NAND2_X1 U1462 ( .A1(n579), .A2(MixColumnsInput[86]), .ZN(n815) );
  NAND2_X1 U1463 ( .A1(n816), .A2(n815), .ZN(RoundOutput[86]) );
  NAND2_X1 U1464 ( .A1(MixColumnsOutput[87]), .A2(n577), .ZN(n818) );
  NAND2_X1 U1465 ( .A1(n579), .A2(MixColumnsInput[87]), .ZN(n817) );
  NAND2_X1 U1466 ( .A1(n818), .A2(n817), .ZN(RoundOutput[87]) );
  NAND2_X1 U1467 ( .A1(MixColumnsOutput[88]), .A2(n577), .ZN(n820) );
  NAND2_X1 U1468 ( .A1(n579), .A2(MixColumnsInput[88]), .ZN(n819) );
  NAND2_X1 U1469 ( .A1(n820), .A2(n819), .ZN(RoundOutput[88]) );
  NAND2_X1 U1470 ( .A1(MixColumnsOutput[89]), .A2(n845), .ZN(n822) );
  NAND2_X1 U1471 ( .A1(n579), .A2(MixColumnsInput[89]), .ZN(n821) );
  NAND2_X1 U1472 ( .A1(n822), .A2(n821), .ZN(RoundOutput[89]) );
  NAND2_X1 U1473 ( .A1(MixColumnsOutput[8]), .A2(n575), .ZN(n824) );
  NAND2_X1 U1474 ( .A1(n579), .A2(MixColumnsInput[8]), .ZN(n823) );
  NAND2_X1 U1475 ( .A1(n824), .A2(n823), .ZN(RoundOutput[8]) );
  NAND2_X1 U1476 ( .A1(MixColumnsOutput[90]), .A2(n574), .ZN(n826) );
  NAND2_X1 U1477 ( .A1(n579), .A2(MixColumnsInput[90]), .ZN(n825) );
  NAND2_X1 U1478 ( .A1(n826), .A2(n825), .ZN(RoundOutput[90]) );
  NAND2_X1 U1479 ( .A1(MixColumnsOutput[91]), .A2(n576), .ZN(n828) );
  NAND2_X1 U1480 ( .A1(n579), .A2(MixColumnsInput[91]), .ZN(n827) );
  NAND2_X1 U1481 ( .A1(n828), .A2(n827), .ZN(RoundOutput[91]) );
  NAND2_X1 U1482 ( .A1(MixColumnsOutput[92]), .A2(n575), .ZN(n830) );
  NAND2_X1 U1483 ( .A1(n579), .A2(MixColumnsInput[92]), .ZN(n829) );
  NAND2_X1 U1484 ( .A1(n830), .A2(n829), .ZN(RoundOutput[92]) );
  NAND2_X1 U1485 ( .A1(MixColumnsOutput[93]), .A2(n577), .ZN(n832) );
  NAND2_X1 U1486 ( .A1(n579), .A2(MixColumnsInput[93]), .ZN(n831) );
  NAND2_X1 U1487 ( .A1(n832), .A2(n831), .ZN(RoundOutput[93]) );
  NAND2_X1 U1488 ( .A1(MixColumnsOutput[94]), .A2(n575), .ZN(n834) );
  NAND2_X1 U1489 ( .A1(n579), .A2(MixColumnsInput[94]), .ZN(n833) );
  NAND2_X1 U1490 ( .A1(n834), .A2(n833), .ZN(RoundOutput[94]) );
  NAND2_X1 U1491 ( .A1(MixColumnsOutput[95]), .A2(n576), .ZN(n836) );
  NAND2_X1 U1492 ( .A1(n579), .A2(MixColumnsInput[95]), .ZN(n835) );
  NAND2_X1 U1493 ( .A1(n836), .A2(n835), .ZN(RoundOutput[95]) );
  NAND2_X1 U1494 ( .A1(MixColumnsOutput[96]), .A2(n577), .ZN(n838) );
  NAND2_X1 U1495 ( .A1(n579), .A2(MixColumnsInput[96]), .ZN(n837) );
  NAND2_X1 U1496 ( .A1(n838), .A2(n837), .ZN(RoundOutput[96]) );
  NAND2_X1 U1497 ( .A1(MixColumnsOutput[97]), .A2(n578), .ZN(n840) );
  NAND2_X1 U1498 ( .A1(n579), .A2(MixColumnsInput[97]), .ZN(n839) );
  NAND2_X1 U1499 ( .A1(n840), .A2(n839), .ZN(RoundOutput[97]) );
  NAND2_X1 U1500 ( .A1(MixColumnsOutput[98]), .A2(n577), .ZN(n842) );
  NAND2_X1 U1501 ( .A1(n579), .A2(MixColumnsInput[98]), .ZN(n841) );
  NAND2_X1 U1502 ( .A1(n842), .A2(n841), .ZN(RoundOutput[98]) );
  NAND2_X1 U1503 ( .A1(MixColumnsOutput[99]), .A2(n574), .ZN(n844) );
  NAND2_X1 U1504 ( .A1(n579), .A2(MixColumnsInput[99]), .ZN(n843) );
  NAND2_X1 U1505 ( .A1(n844), .A2(n843), .ZN(RoundOutput[99]) );
  NAND2_X1 U1506 ( .A1(MixColumnsOutput[9]), .A2(n578), .ZN(n847) );
  NAND2_X1 U1507 ( .A1(n579), .A2(MixColumnsInput[9]), .ZN(n846) );
  NAND2_X1 U1508 ( .A1(n847), .A2(n846), .ZN(RoundOutput[9]) );
  XOR2_X1 U1509 ( .A(key_shifted[8]), .B(state_shifted[8]), .Z(
        SubBytesInput[0]) );
  XOR2_X1 U1510 ( .A(key_shifted[108]), .B(state_shifted[108]), .Z(
        SubBytesInput[100]) );
  XOR2_X1 U1511 ( .A(key_shifted[109]), .B(state_shifted[109]), .Z(
        SubBytesInput[101]) );
  XOR2_X1 U1512 ( .A(key_shifted[110]), .B(state_shifted[110]), .Z(
        SubBytesInput[102]) );
  XOR2_X1 U1513 ( .A(key_shifted[111]), .B(state_shifted[111]), .Z(
        SubBytesInput[103]) );
  XOR2_X1 U1514 ( .A(key_shifted[112]), .B(state_shifted[112]), .Z(
        SubBytesInput[104]) );
  XOR2_X1 U1515 ( .A(key_shifted[113]), .B(state_shifted[113]), .Z(
        SubBytesInput[105]) );
  XOR2_X1 U1516 ( .A(key_shifted[114]), .B(state_shifted[114]), .Z(
        SubBytesInput[106]) );
  XOR2_X1 U1517 ( .A(key_shifted[115]), .B(state_shifted[115]), .Z(
        SubBytesInput[107]) );
  XOR2_X1 U1518 ( .A(key_shifted[116]), .B(state_shifted[116]), .Z(
        SubBytesInput[108]) );
  XOR2_X1 U1519 ( .A(key_shifted[117]), .B(state_shifted[117]), .Z(
        SubBytesInput[109]) );
  XOR2_X1 U1520 ( .A(key_shifted[18]), .B(state_shifted[18]), .Z(
        SubBytesInput[10]) );
  XOR2_X1 U1521 ( .A(key_shifted[118]), .B(state_shifted[118]), .Z(
        SubBytesInput[110]) );
  XOR2_X1 U1522 ( .A(key_shifted[119]), .B(state_shifted[119]), .Z(
        SubBytesInput[111]) );
  XOR2_X1 U1523 ( .A(key_shifted[120]), .B(state_shifted[120]), .Z(
        SubBytesInput[112]) );
  XOR2_X1 U1524 ( .A(key_shifted[121]), .B(state_shifted[121]), .Z(
        SubBytesInput[113]) );
  XOR2_X1 U1525 ( .A(key_shifted[122]), .B(state_shifted[122]), .Z(
        SubBytesInput[114]) );
  XOR2_X1 U1526 ( .A(key_shifted[123]), .B(state_shifted[123]), .Z(
        SubBytesInput[115]) );
  XOR2_X1 U1527 ( .A(key_shifted[124]), .B(state_shifted[124]), .Z(
        SubBytesInput[116]) );
  XOR2_X1 U1528 ( .A(key_shifted[125]), .B(state_shifted[125]), .Z(
        SubBytesInput[117]) );
  XOR2_X1 U1529 ( .A(key_shifted[126]), .B(state_shifted[126]), .Z(
        SubBytesInput[118]) );
  XOR2_X1 U1530 ( .A(key_shifted[127]), .B(state_shifted[127]), .Z(
        SubBytesInput[119]) );
  XOR2_X1 U1531 ( .A(key_shifted[19]), .B(state_shifted[19]), .Z(
        SubBytesInput[11]) );
  XOR2_X1 U1532 ( .A(key_shifted[20]), .B(state_shifted[20]), .Z(
        SubBytesInput[12]) );
  XOR2_X1 U1533 ( .A(key_shifted[21]), .B(state_shifted[21]), .Z(
        SubBytesInput[13]) );
  XOR2_X1 U1534 ( .A(key_shifted[22]), .B(state_shifted[22]), .Z(
        SubBytesInput[14]) );
  XOR2_X1 U1535 ( .A(key_shifted[23]), .B(state_shifted[23]), .Z(
        SubBytesInput[15]) );
  XOR2_X1 U1536 ( .A(key_shifted[24]), .B(state_shifted[24]), .Z(
        SubBytesInput[16]) );
  XOR2_X1 U1537 ( .A(key_shifted[25]), .B(state_shifted[25]), .Z(
        SubBytesInput[17]) );
  XOR2_X1 U1538 ( .A(key_shifted[26]), .B(state_shifted[26]), .Z(
        SubBytesInput[18]) );
  XOR2_X1 U1539 ( .A(key_shifted[27]), .B(state_shifted[27]), .Z(
        SubBytesInput[19]) );
  XOR2_X1 U1540 ( .A(key_shifted[9]), .B(state_shifted[9]), .Z(
        SubBytesInput[1]) );
  XOR2_X1 U1541 ( .A(key_shifted[28]), .B(state_shifted[28]), .Z(
        SubBytesInput[20]) );
  XOR2_X1 U1542 ( .A(key_shifted[29]), .B(state_shifted[29]), .Z(
        SubBytesInput[21]) );
  XOR2_X1 U1543 ( .A(key_shifted[30]), .B(state_shifted[30]), .Z(
        SubBytesInput[22]) );
  XOR2_X1 U1544 ( .A(key_shifted[31]), .B(state_shifted[31]), .Z(
        SubBytesInput[23]) );
  XOR2_X1 U1545 ( .A(key_shifted[32]), .B(state_shifted[32]), .Z(
        SubBytesInput[24]) );
  XOR2_X1 U1546 ( .A(key_shifted[33]), .B(state_shifted[33]), .Z(
        SubBytesInput[25]) );
  XOR2_X1 U1547 ( .A(key_shifted[34]), .B(state_shifted[34]), .Z(
        SubBytesInput[26]) );
  XOR2_X1 U1548 ( .A(key_shifted[35]), .B(state_shifted[35]), .Z(
        SubBytesInput[27]) );
  XOR2_X1 U1549 ( .A(key_shifted[36]), .B(state_shifted[36]), .Z(
        SubBytesInput[28]) );
  XOR2_X1 U1550 ( .A(key_shifted[37]), .B(state_shifted[37]), .Z(
        SubBytesInput[29]) );
  XOR2_X1 U1551 ( .A(key_shifted[10]), .B(state_shifted[10]), .Z(
        SubBytesInput[2]) );
  XOR2_X1 U1552 ( .A(key_shifted[38]), .B(state_shifted[38]), .Z(
        SubBytesInput[30]) );
  XOR2_X1 U1553 ( .A(key_shifted[39]), .B(state_shifted[39]), .Z(
        SubBytesInput[31]) );
  XOR2_X1 U1554 ( .A(key_shifted[40]), .B(state_shifted[40]), .Z(
        SubBytesInput[32]) );
  XOR2_X1 U1555 ( .A(key_shifted[41]), .B(state_shifted[41]), .Z(
        SubBytesInput[33]) );
  XOR2_X1 U1556 ( .A(key_shifted[42]), .B(state_shifted[42]), .Z(
        SubBytesInput[34]) );
  XOR2_X1 U1557 ( .A(key_shifted[43]), .B(state_shifted[43]), .Z(
        SubBytesInput[35]) );
  XOR2_X1 U1558 ( .A(key_shifted[44]), .B(state_shifted[44]), .Z(
        SubBytesInput[36]) );
  XOR2_X1 U1559 ( .A(key_shifted[45]), .B(state_shifted[45]), .Z(
        SubBytesInput[37]) );
  XOR2_X1 U1560 ( .A(key_shifted[46]), .B(state_shifted[46]), .Z(
        SubBytesInput[38]) );
  XOR2_X1 U1561 ( .A(key_shifted[47]), .B(state_shifted[47]), .Z(
        SubBytesInput[39]) );
  XOR2_X1 U1562 ( .A(key_shifted[11]), .B(state_shifted[11]), .Z(
        SubBytesInput[3]) );
  XOR2_X1 U1563 ( .A(key_shifted[48]), .B(state_shifted[48]), .Z(
        SubBytesInput[40]) );
  XOR2_X1 U1564 ( .A(key_shifted[49]), .B(state_shifted[49]), .Z(
        SubBytesInput[41]) );
  XOR2_X1 U1565 ( .A(key_shifted[50]), .B(state_shifted[50]), .Z(
        SubBytesInput[42]) );
  XOR2_X1 U1566 ( .A(key_shifted[51]), .B(state_shifted[51]), .Z(
        SubBytesInput[43]) );
  XOR2_X1 U1567 ( .A(key_shifted[52]), .B(state_shifted[52]), .Z(
        SubBytesInput[44]) );
  XOR2_X1 U1568 ( .A(key_shifted[53]), .B(state_shifted[53]), .Z(
        SubBytesInput[45]) );
  XOR2_X1 U1569 ( .A(key_shifted[54]), .B(state_shifted[54]), .Z(
        SubBytesInput[46]) );
  XOR2_X1 U1570 ( .A(key_shifted[55]), .B(state_shifted[55]), .Z(
        SubBytesInput[47]) );
  XOR2_X1 U1571 ( .A(key_shifted[56]), .B(state_shifted[56]), .Z(
        SubBytesInput[48]) );
  XOR2_X1 U1572 ( .A(key_shifted[57]), .B(state_shifted[57]), .Z(
        SubBytesInput[49]) );
  XOR2_X1 U1573 ( .A(key_shifted[12]), .B(state_shifted[12]), .Z(
        SubBytesInput[4]) );
  XOR2_X1 U1574 ( .A(key_shifted[58]), .B(state_shifted[58]), .Z(
        SubBytesInput[50]) );
  XOR2_X1 U1575 ( .A(key_shifted[59]), .B(state_shifted[59]), .Z(
        SubBytesInput[51]) );
  XOR2_X1 U1576 ( .A(key_shifted[60]), .B(state_shifted[60]), .Z(
        SubBytesInput[52]) );
  XOR2_X1 U1577 ( .A(key_shifted[61]), .B(state_shifted[61]), .Z(
        SubBytesInput[53]) );
  XOR2_X1 U1578 ( .A(key_shifted[62]), .B(state_shifted[62]), .Z(
        SubBytesInput[54]) );
  XOR2_X1 U1579 ( .A(key_shifted[63]), .B(state_shifted[63]), .Z(
        SubBytesInput[55]) );
  XOR2_X1 U1580 ( .A(key_shifted[64]), .B(state_shifted[64]), .Z(
        SubBytesInput[56]) );
  XOR2_X1 U1581 ( .A(key_shifted[65]), .B(state_shifted[65]), .Z(
        SubBytesInput[57]) );
  XOR2_X1 U1582 ( .A(key_shifted[66]), .B(state_shifted[66]), .Z(
        SubBytesInput[58]) );
  XOR2_X1 U1583 ( .A(key_shifted[67]), .B(state_shifted[67]), .Z(
        SubBytesInput[59]) );
  XOR2_X1 U1584 ( .A(key_shifted[13]), .B(state_shifted[13]), .Z(
        SubBytesInput[5]) );
  XOR2_X1 U1585 ( .A(key_shifted[68]), .B(state_shifted[68]), .Z(
        SubBytesInput[60]) );
  XOR2_X1 U1586 ( .A(key_shifted[69]), .B(state_shifted[69]), .Z(
        SubBytesInput[61]) );
  XOR2_X1 U1587 ( .A(key_shifted[70]), .B(state_shifted[70]), .Z(
        SubBytesInput[62]) );
  XOR2_X1 U1588 ( .A(key_shifted[71]), .B(state_shifted[71]), .Z(
        SubBytesInput[63]) );
  XOR2_X1 U1589 ( .A(key_shifted[72]), .B(state_shifted[72]), .Z(
        SubBytesInput[64]) );
  XOR2_X1 U1590 ( .A(key_shifted[73]), .B(state_shifted[73]), .Z(
        SubBytesInput[65]) );
  XOR2_X1 U1591 ( .A(key_shifted[74]), .B(state_shifted[74]), .Z(
        SubBytesInput[66]) );
  XOR2_X1 U1592 ( .A(key_shifted[75]), .B(state_shifted[75]), .Z(
        SubBytesInput[67]) );
  XOR2_X1 U1593 ( .A(key_shifted[76]), .B(state_shifted[76]), .Z(
        SubBytesInput[68]) );
  XOR2_X1 U1594 ( .A(key_shifted[77]), .B(state_shifted[77]), .Z(
        SubBytesInput[69]) );
  XOR2_X1 U1595 ( .A(key_shifted[14]), .B(state_shifted[14]), .Z(
        SubBytesInput[6]) );
  XOR2_X1 U1596 ( .A(key_shifted[78]), .B(state_shifted[78]), .Z(
        SubBytesInput[70]) );
  XOR2_X1 U1597 ( .A(key_shifted[79]), .B(state_shifted[79]), .Z(
        SubBytesInput[71]) );
  XOR2_X1 U1598 ( .A(key_shifted[80]), .B(state_shifted[80]), .Z(
        SubBytesInput[72]) );
  XOR2_X1 U1599 ( .A(key_shifted[81]), .B(state_shifted[81]), .Z(
        SubBytesInput[73]) );
  XOR2_X1 U1600 ( .A(key_shifted[82]), .B(state_shifted[82]), .Z(
        SubBytesInput[74]) );
  XOR2_X1 U1601 ( .A(key_shifted[83]), .B(state_shifted[83]), .Z(
        SubBytesInput[75]) );
  XOR2_X1 U1602 ( .A(key_shifted[84]), .B(state_shifted[84]), .Z(
        SubBytesInput[76]) );
  XOR2_X1 U1603 ( .A(key_shifted[85]), .B(state_shifted[85]), .Z(
        SubBytesInput[77]) );
  XOR2_X1 U1604 ( .A(key_shifted[86]), .B(state_shifted[86]), .Z(
        SubBytesInput[78]) );
  XOR2_X1 U1605 ( .A(key_shifted[87]), .B(state_shifted[87]), .Z(
        SubBytesInput[79]) );
  XOR2_X1 U1606 ( .A(key_shifted[15]), .B(state_shifted[15]), .Z(
        SubBytesInput[7]) );
  XOR2_X1 U1607 ( .A(key_shifted[88]), .B(state_shifted[88]), .Z(
        SubBytesInput[80]) );
  XOR2_X1 U1608 ( .A(key_shifted[89]), .B(state_shifted[89]), .Z(
        SubBytesInput[81]) );
  XOR2_X1 U1609 ( .A(key_shifted[90]), .B(state_shifted[90]), .Z(
        SubBytesInput[82]) );
  XOR2_X1 U1610 ( .A(key_shifted[91]), .B(state_shifted[91]), .Z(
        SubBytesInput[83]) );
  XOR2_X1 U1611 ( .A(key_shifted[92]), .B(state_shifted[92]), .Z(
        SubBytesInput[84]) );
  XOR2_X1 U1612 ( .A(key_shifted[93]), .B(state_shifted[93]), .Z(
        SubBytesInput[85]) );
  XOR2_X1 U1613 ( .A(key_shifted[94]), .B(state_shifted[94]), .Z(
        SubBytesInput[86]) );
  XOR2_X1 U1614 ( .A(key_shifted[95]), .B(state_shifted[95]), .Z(
        SubBytesInput[87]) );
  XOR2_X1 U1615 ( .A(key_shifted[96]), .B(state_shifted[96]), .Z(
        SubBytesInput[88]) );
  XOR2_X1 U1616 ( .A(key_shifted[97]), .B(state_shifted[97]), .Z(
        SubBytesInput[89]) );
  XOR2_X1 U1617 ( .A(key_shifted[16]), .B(state_shifted[16]), .Z(
        SubBytesInput[8]) );
  XOR2_X1 U1618 ( .A(key_shifted[98]), .B(state_shifted[98]), .Z(
        SubBytesInput[90]) );
  XOR2_X1 U1619 ( .A(key_shifted[99]), .B(state_shifted[99]), .Z(
        SubBytesInput[91]) );
  XOR2_X1 U1620 ( .A(key_shifted[100]), .B(state_shifted[100]), .Z(
        SubBytesInput[92]) );
  XOR2_X1 U1621 ( .A(key_shifted[101]), .B(state_shifted[101]), .Z(
        SubBytesInput[93]) );
  XOR2_X1 U1622 ( .A(key_shifted[102]), .B(state_shifted[102]), .Z(
        SubBytesInput[94]) );
  XOR2_X1 U1623 ( .A(key_shifted[103]), .B(state_shifted[103]), .Z(
        SubBytesInput[95]) );
  XOR2_X1 U1624 ( .A(key_shifted[104]), .B(state_shifted[104]), .Z(
        SubBytesInput[96]) );
  XOR2_X1 U1625 ( .A(key_shifted[105]), .B(state_shifted[105]), .Z(
        SubBytesInput[97]) );
  XOR2_X1 U1626 ( .A(key_shifted[106]), .B(state_shifted[106]), .Z(
        SubBytesInput[98]) );
  XOR2_X1 U1627 ( .A(key_shifted[107]), .B(state_shifted[107]), .Z(
        SubBytesInput[99]) );
  XOR2_X1 U1628 ( .A(key_shifted[17]), .B(state_shifted[17]), .Z(
        SubBytesInput[9]) );
  AND2_X1 U1629 ( .A1(RoundCounter[2]), .A2(n848), .ZN(n286) );
  NAND2_X1 U1630 ( .A1(RoundCounter[1]), .A2(n849), .ZN(n850) );
  NOR2_X1 U1631 ( .A1(n851), .A2(n850), .ZN(n287) );
  XOR2_X1 U1632 ( .A(RoundInput[120]), .B(RoundKey[120]), .Z(port_out[0]) );
  XOR2_X1 U1633 ( .A(RoundInput[121]), .B(RoundKey[121]), .Z(port_out[1]) );
  XOR2_X1 U1634 ( .A(RoundInput[122]), .B(RoundKey[122]), .Z(port_out[2]) );
  XOR2_X1 U1635 ( .A(RoundInput[123]), .B(RoundKey[123]), .Z(port_out[3]) );
  XOR2_X1 U1636 ( .A(RoundInput[124]), .B(RoundKey[124]), .Z(port_out[4]) );
  XOR2_X1 U1637 ( .A(RoundInput[125]), .B(RoundKey[125]), .Z(port_out[5]) );
  XOR2_X1 U1638 ( .A(RoundInput[126]), .B(RoundKey[126]), .Z(port_out[6]) );
  XOR2_X1 U1639 ( .A(RoundInput[127]), .B(RoundKey[127]), .Z(port_out[7]) );
endmodule

