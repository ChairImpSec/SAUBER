/* modified netlist. Source: module SkinnyTop in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/9-Skinny64_64_round_based_encryption_PortParallel/4-AGEMA/SkinnyTop.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module SkinnyTop_SAUBER_Pipeline_d1 (Plaintext_s0_t, Key_s0_t, rst_t, Key_s0_f, Key_s1_t, Key_s1_f, rst_f, Plaintext_s0_f, Plaintext_s1_t, Plaintext_s1_f, Ciphertext_s0_t, done_t, Ciphertext_s0_f, Ciphertext_s1_t, Ciphertext_s1_f, done_f);
    input [63:0] Plaintext_s0_t ;
    input [63:0] Key_s0_t ;
    input rst_t ;
    input [63:0] Key_s0_f ;
    input [63:0] Key_s1_t ;
    input [63:0] Key_s1_f ;
    input rst_f ;
    input [63:0] Plaintext_s0_f ;
    input [63:0] Plaintext_s1_t ;
    input [63:0] Plaintext_s1_f ;
    output [63:0] Ciphertext_s0_t ;
    output done_t ;
    output [63:0] Ciphertext_s0_f ;
    output [63:0] Ciphertext_s1_t ;
    output [63:0] Ciphertext_s1_f ;
    output done_f ;
    wire PlaintextMUX_MUXInst_0_U1_Y ;
    wire PlaintextMUX_MUXInst_0_U1_X ;
    wire PlaintextMUX_MUXInst_1_U1_Y ;
    wire PlaintextMUX_MUXInst_1_U1_X ;
    wire PlaintextMUX_MUXInst_2_U1_Y ;
    wire PlaintextMUX_MUXInst_2_U1_X ;
    wire PlaintextMUX_MUXInst_3_U1_Y ;
    wire PlaintextMUX_MUXInst_3_U1_X ;
    wire PlaintextMUX_MUXInst_4_U1_Y ;
    wire PlaintextMUX_MUXInst_4_U1_X ;
    wire PlaintextMUX_MUXInst_5_U1_Y ;
    wire PlaintextMUX_MUXInst_5_U1_X ;
    wire PlaintextMUX_MUXInst_6_U1_Y ;
    wire PlaintextMUX_MUXInst_6_U1_X ;
    wire PlaintextMUX_MUXInst_7_U1_Y ;
    wire PlaintextMUX_MUXInst_7_U1_X ;
    wire PlaintextMUX_MUXInst_8_U1_Y ;
    wire PlaintextMUX_MUXInst_8_U1_X ;
    wire PlaintextMUX_MUXInst_9_U1_Y ;
    wire PlaintextMUX_MUXInst_9_U1_X ;
    wire PlaintextMUX_MUXInst_10_U1_Y ;
    wire PlaintextMUX_MUXInst_10_U1_X ;
    wire PlaintextMUX_MUXInst_11_U1_Y ;
    wire PlaintextMUX_MUXInst_11_U1_X ;
    wire PlaintextMUX_MUXInst_12_U1_Y ;
    wire PlaintextMUX_MUXInst_12_U1_X ;
    wire PlaintextMUX_MUXInst_13_U1_Y ;
    wire PlaintextMUX_MUXInst_13_U1_X ;
    wire PlaintextMUX_MUXInst_14_U1_Y ;
    wire PlaintextMUX_MUXInst_14_U1_X ;
    wire PlaintextMUX_MUXInst_15_U1_Y ;
    wire PlaintextMUX_MUXInst_15_U1_X ;
    wire PlaintextMUX_MUXInst_16_U1_Y ;
    wire PlaintextMUX_MUXInst_16_U1_X ;
    wire PlaintextMUX_MUXInst_17_U1_Y ;
    wire PlaintextMUX_MUXInst_17_U1_X ;
    wire PlaintextMUX_MUXInst_18_U1_Y ;
    wire PlaintextMUX_MUXInst_18_U1_X ;
    wire PlaintextMUX_MUXInst_19_U1_Y ;
    wire PlaintextMUX_MUXInst_19_U1_X ;
    wire PlaintextMUX_MUXInst_20_U1_Y ;
    wire PlaintextMUX_MUXInst_20_U1_X ;
    wire PlaintextMUX_MUXInst_21_U1_Y ;
    wire PlaintextMUX_MUXInst_21_U1_X ;
    wire PlaintextMUX_MUXInst_22_U1_Y ;
    wire PlaintextMUX_MUXInst_22_U1_X ;
    wire PlaintextMUX_MUXInst_23_U1_Y ;
    wire PlaintextMUX_MUXInst_23_U1_X ;
    wire PlaintextMUX_MUXInst_24_U1_Y ;
    wire PlaintextMUX_MUXInst_24_U1_X ;
    wire PlaintextMUX_MUXInst_25_U1_Y ;
    wire PlaintextMUX_MUXInst_25_U1_X ;
    wire PlaintextMUX_MUXInst_26_U1_Y ;
    wire PlaintextMUX_MUXInst_26_U1_X ;
    wire PlaintextMUX_MUXInst_27_U1_Y ;
    wire PlaintextMUX_MUXInst_27_U1_X ;
    wire PlaintextMUX_MUXInst_28_U1_Y ;
    wire PlaintextMUX_MUXInst_28_U1_X ;
    wire PlaintextMUX_MUXInst_29_U1_Y ;
    wire PlaintextMUX_MUXInst_29_U1_X ;
    wire PlaintextMUX_MUXInst_30_U1_Y ;
    wire PlaintextMUX_MUXInst_30_U1_X ;
    wire PlaintextMUX_MUXInst_31_U1_Y ;
    wire PlaintextMUX_MUXInst_31_U1_X ;
    wire PlaintextMUX_MUXInst_32_U1_Y ;
    wire PlaintextMUX_MUXInst_32_U1_X ;
    wire PlaintextMUX_MUXInst_33_U1_Y ;
    wire PlaintextMUX_MUXInst_33_U1_X ;
    wire PlaintextMUX_MUXInst_34_U1_Y ;
    wire PlaintextMUX_MUXInst_34_U1_X ;
    wire PlaintextMUX_MUXInst_35_U1_Y ;
    wire PlaintextMUX_MUXInst_35_U1_X ;
    wire PlaintextMUX_MUXInst_36_U1_Y ;
    wire PlaintextMUX_MUXInst_36_U1_X ;
    wire PlaintextMUX_MUXInst_37_U1_Y ;
    wire PlaintextMUX_MUXInst_37_U1_X ;
    wire PlaintextMUX_MUXInst_38_U1_Y ;
    wire PlaintextMUX_MUXInst_38_U1_X ;
    wire PlaintextMUX_MUXInst_39_U1_Y ;
    wire PlaintextMUX_MUXInst_39_U1_X ;
    wire PlaintextMUX_MUXInst_40_U1_Y ;
    wire PlaintextMUX_MUXInst_40_U1_X ;
    wire PlaintextMUX_MUXInst_41_U1_Y ;
    wire PlaintextMUX_MUXInst_41_U1_X ;
    wire PlaintextMUX_MUXInst_42_U1_Y ;
    wire PlaintextMUX_MUXInst_42_U1_X ;
    wire PlaintextMUX_MUXInst_43_U1_Y ;
    wire PlaintextMUX_MUXInst_43_U1_X ;
    wire PlaintextMUX_MUXInst_44_U1_Y ;
    wire PlaintextMUX_MUXInst_44_U1_X ;
    wire PlaintextMUX_MUXInst_45_U1_Y ;
    wire PlaintextMUX_MUXInst_45_U1_X ;
    wire PlaintextMUX_MUXInst_46_U1_Y ;
    wire PlaintextMUX_MUXInst_46_U1_X ;
    wire PlaintextMUX_MUXInst_47_U1_Y ;
    wire PlaintextMUX_MUXInst_47_U1_X ;
    wire PlaintextMUX_MUXInst_48_U1_Y ;
    wire PlaintextMUX_MUXInst_48_U1_X ;
    wire PlaintextMUX_MUXInst_49_U1_Y ;
    wire PlaintextMUX_MUXInst_49_U1_X ;
    wire PlaintextMUX_MUXInst_50_U1_Y ;
    wire PlaintextMUX_MUXInst_50_U1_X ;
    wire PlaintextMUX_MUXInst_51_U1_Y ;
    wire PlaintextMUX_MUXInst_51_U1_X ;
    wire PlaintextMUX_MUXInst_52_U1_Y ;
    wire PlaintextMUX_MUXInst_52_U1_X ;
    wire PlaintextMUX_MUXInst_53_U1_Y ;
    wire PlaintextMUX_MUXInst_53_U1_X ;
    wire PlaintextMUX_MUXInst_54_U1_Y ;
    wire PlaintextMUX_MUXInst_54_U1_X ;
    wire PlaintextMUX_MUXInst_55_U1_Y ;
    wire PlaintextMUX_MUXInst_55_U1_X ;
    wire PlaintextMUX_MUXInst_56_U1_Y ;
    wire PlaintextMUX_MUXInst_56_U1_X ;
    wire PlaintextMUX_MUXInst_57_U1_Y ;
    wire PlaintextMUX_MUXInst_57_U1_X ;
    wire PlaintextMUX_MUXInst_58_U1_Y ;
    wire PlaintextMUX_MUXInst_58_U1_X ;
    wire PlaintextMUX_MUXInst_59_U1_Y ;
    wire PlaintextMUX_MUXInst_59_U1_X ;
    wire PlaintextMUX_MUXInst_60_U1_Y ;
    wire PlaintextMUX_MUXInst_60_U1_X ;
    wire PlaintextMUX_MUXInst_61_U1_Y ;
    wire PlaintextMUX_MUXInst_61_U1_X ;
    wire PlaintextMUX_MUXInst_62_U1_Y ;
    wire PlaintextMUX_MUXInst_62_U1_X ;
    wire PlaintextMUX_MUXInst_63_U1_Y ;
    wire PlaintextMUX_MUXInst_63_U1_X ;
    wire SubCellInst_SboxInst_0_L3 ;
    wire SubCellInst_SboxInst_0_YY_3 ;
    wire SubCellInst_SboxInst_0_L2 ;
    wire SubCellInst_SboxInst_0_T3 ;
    wire SubCellInst_SboxInst_0_Q7 ;
    wire SubCellInst_SboxInst_0_L1 ;
    wire SubCellInst_SboxInst_0_Q6 ;
    wire SubCellInst_SboxInst_0_L0 ;
    wire SubCellInst_SboxInst_0_T2 ;
    wire SubCellInst_SboxInst_0_Q4 ;
    wire SubCellInst_SboxInst_0_T1 ;
    wire SubCellInst_SboxInst_0_Q2 ;
    wire SubCellInst_SboxInst_0_T0 ;
    wire SubCellInst_SboxInst_0_Q1 ;
    wire SubCellInst_SboxInst_0_Q0 ;
    wire SubCellInst_SboxInst_1_L3 ;
    wire SubCellInst_SboxInst_1_YY_3 ;
    wire SubCellInst_SboxInst_1_L2 ;
    wire SubCellInst_SboxInst_1_T3 ;
    wire SubCellInst_SboxInst_1_Q7 ;
    wire SubCellInst_SboxInst_1_L1 ;
    wire SubCellInst_SboxInst_1_Q6 ;
    wire SubCellInst_SboxInst_1_L0 ;
    wire SubCellInst_SboxInst_1_T2 ;
    wire SubCellInst_SboxInst_1_Q4 ;
    wire SubCellInst_SboxInst_1_T1 ;
    wire SubCellInst_SboxInst_1_Q2 ;
    wire SubCellInst_SboxInst_1_T0 ;
    wire SubCellInst_SboxInst_1_Q1 ;
    wire SubCellInst_SboxInst_1_Q0 ;
    wire SubCellInst_SboxInst_2_L3 ;
    wire SubCellInst_SboxInst_2_YY_3 ;
    wire SubCellInst_SboxInst_2_L2 ;
    wire SubCellInst_SboxInst_2_T3 ;
    wire SubCellInst_SboxInst_2_Q7 ;
    wire SubCellInst_SboxInst_2_L1 ;
    wire SubCellInst_SboxInst_2_Q6 ;
    wire SubCellInst_SboxInst_2_L0 ;
    wire SubCellInst_SboxInst_2_T2 ;
    wire SubCellInst_SboxInst_2_Q4 ;
    wire SubCellInst_SboxInst_2_T1 ;
    wire SubCellInst_SboxInst_2_Q2 ;
    wire SubCellInst_SboxInst_2_T0 ;
    wire SubCellInst_SboxInst_2_Q1 ;
    wire SubCellInst_SboxInst_2_Q0 ;
    wire SubCellInst_SboxInst_3_L3 ;
    wire SubCellInst_SboxInst_3_YY_3 ;
    wire SubCellInst_SboxInst_3_L2 ;
    wire SubCellInst_SboxInst_3_T3 ;
    wire SubCellInst_SboxInst_3_Q7 ;
    wire SubCellInst_SboxInst_3_L1 ;
    wire SubCellInst_SboxInst_3_Q6 ;
    wire SubCellInst_SboxInst_3_L0 ;
    wire SubCellInst_SboxInst_3_T2 ;
    wire SubCellInst_SboxInst_3_Q4 ;
    wire SubCellInst_SboxInst_3_T1 ;
    wire SubCellInst_SboxInst_3_Q2 ;
    wire SubCellInst_SboxInst_3_T0 ;
    wire SubCellInst_SboxInst_3_Q1 ;
    wire SubCellInst_SboxInst_3_Q0 ;
    wire SubCellInst_SboxInst_4_L3 ;
    wire SubCellInst_SboxInst_4_YY_3 ;
    wire SubCellInst_SboxInst_4_L2 ;
    wire SubCellInst_SboxInst_4_T3 ;
    wire SubCellInst_SboxInst_4_Q7 ;
    wire SubCellInst_SboxInst_4_L1 ;
    wire SubCellInst_SboxInst_4_Q6 ;
    wire SubCellInst_SboxInst_4_L0 ;
    wire SubCellInst_SboxInst_4_T2 ;
    wire SubCellInst_SboxInst_4_Q4 ;
    wire SubCellInst_SboxInst_4_T1 ;
    wire SubCellInst_SboxInst_4_Q2 ;
    wire SubCellInst_SboxInst_4_T0 ;
    wire SubCellInst_SboxInst_4_Q1 ;
    wire SubCellInst_SboxInst_4_Q0 ;
    wire SubCellInst_SboxInst_5_L3 ;
    wire SubCellInst_SboxInst_5_YY_3 ;
    wire SubCellInst_SboxInst_5_L2 ;
    wire SubCellInst_SboxInst_5_T3 ;
    wire SubCellInst_SboxInst_5_Q7 ;
    wire SubCellInst_SboxInst_5_L1 ;
    wire SubCellInst_SboxInst_5_Q6 ;
    wire SubCellInst_SboxInst_5_L0 ;
    wire SubCellInst_SboxInst_5_T2 ;
    wire SubCellInst_SboxInst_5_Q4 ;
    wire SubCellInst_SboxInst_5_T1 ;
    wire SubCellInst_SboxInst_5_Q2 ;
    wire SubCellInst_SboxInst_5_T0 ;
    wire SubCellInst_SboxInst_5_Q1 ;
    wire SubCellInst_SboxInst_5_Q0 ;
    wire SubCellInst_SboxInst_6_L3 ;
    wire SubCellInst_SboxInst_6_YY_3 ;
    wire SubCellInst_SboxInst_6_L2 ;
    wire SubCellInst_SboxInst_6_T3 ;
    wire SubCellInst_SboxInst_6_Q7 ;
    wire SubCellInst_SboxInst_6_L1 ;
    wire SubCellInst_SboxInst_6_Q6 ;
    wire SubCellInst_SboxInst_6_L0 ;
    wire SubCellInst_SboxInst_6_T2 ;
    wire SubCellInst_SboxInst_6_Q4 ;
    wire SubCellInst_SboxInst_6_T1 ;
    wire SubCellInst_SboxInst_6_Q2 ;
    wire SubCellInst_SboxInst_6_T0 ;
    wire SubCellInst_SboxInst_6_Q1 ;
    wire SubCellInst_SboxInst_6_Q0 ;
    wire SubCellInst_SboxInst_7_L3 ;
    wire SubCellInst_SboxInst_7_YY_3 ;
    wire SubCellInst_SboxInst_7_L2 ;
    wire SubCellInst_SboxInst_7_T3 ;
    wire SubCellInst_SboxInst_7_Q7 ;
    wire SubCellInst_SboxInst_7_L1 ;
    wire SubCellInst_SboxInst_7_Q6 ;
    wire SubCellInst_SboxInst_7_L0 ;
    wire SubCellInst_SboxInst_7_T2 ;
    wire SubCellInst_SboxInst_7_Q4 ;
    wire SubCellInst_SboxInst_7_T1 ;
    wire SubCellInst_SboxInst_7_Q2 ;
    wire SubCellInst_SboxInst_7_T0 ;
    wire SubCellInst_SboxInst_7_Q1 ;
    wire SubCellInst_SboxInst_7_Q0 ;
    wire SubCellInst_SboxInst_8_L3 ;
    wire SubCellInst_SboxInst_8_YY_3 ;
    wire SubCellInst_SboxInst_8_L2 ;
    wire SubCellInst_SboxInst_8_T3 ;
    wire SubCellInst_SboxInst_8_Q7 ;
    wire SubCellInst_SboxInst_8_L1 ;
    wire SubCellInst_SboxInst_8_Q6 ;
    wire SubCellInst_SboxInst_8_L0 ;
    wire SubCellInst_SboxInst_8_T2 ;
    wire SubCellInst_SboxInst_8_Q4 ;
    wire SubCellInst_SboxInst_8_T1 ;
    wire SubCellInst_SboxInst_8_Q2 ;
    wire SubCellInst_SboxInst_8_T0 ;
    wire SubCellInst_SboxInst_8_Q1 ;
    wire SubCellInst_SboxInst_8_Q0 ;
    wire SubCellInst_SboxInst_9_L3 ;
    wire SubCellInst_SboxInst_9_YY_3 ;
    wire SubCellInst_SboxInst_9_L2 ;
    wire SubCellInst_SboxInst_9_T3 ;
    wire SubCellInst_SboxInst_9_Q7 ;
    wire SubCellInst_SboxInst_9_L1 ;
    wire SubCellInst_SboxInst_9_Q6 ;
    wire SubCellInst_SboxInst_9_L0 ;
    wire SubCellInst_SboxInst_9_T2 ;
    wire SubCellInst_SboxInst_9_Q4 ;
    wire SubCellInst_SboxInst_9_T1 ;
    wire SubCellInst_SboxInst_9_Q2 ;
    wire SubCellInst_SboxInst_9_T0 ;
    wire SubCellInst_SboxInst_9_Q1 ;
    wire SubCellInst_SboxInst_9_Q0 ;
    wire SubCellInst_SboxInst_10_L3 ;
    wire SubCellInst_SboxInst_10_YY_3 ;
    wire SubCellInst_SboxInst_10_L2 ;
    wire SubCellInst_SboxInst_10_T3 ;
    wire SubCellInst_SboxInst_10_Q7 ;
    wire SubCellInst_SboxInst_10_L1 ;
    wire SubCellInst_SboxInst_10_Q6 ;
    wire SubCellInst_SboxInst_10_L0 ;
    wire SubCellInst_SboxInst_10_T2 ;
    wire SubCellInst_SboxInst_10_Q4 ;
    wire SubCellInst_SboxInst_10_T1 ;
    wire SubCellInst_SboxInst_10_Q2 ;
    wire SubCellInst_SboxInst_10_T0 ;
    wire SubCellInst_SboxInst_10_Q1 ;
    wire SubCellInst_SboxInst_10_Q0 ;
    wire SubCellInst_SboxInst_11_L3 ;
    wire SubCellInst_SboxInst_11_YY_3 ;
    wire SubCellInst_SboxInst_11_L2 ;
    wire SubCellInst_SboxInst_11_T3 ;
    wire SubCellInst_SboxInst_11_Q7 ;
    wire SubCellInst_SboxInst_11_L1 ;
    wire SubCellInst_SboxInst_11_Q6 ;
    wire SubCellInst_SboxInst_11_L0 ;
    wire SubCellInst_SboxInst_11_T2 ;
    wire SubCellInst_SboxInst_11_Q4 ;
    wire SubCellInst_SboxInst_11_T1 ;
    wire SubCellInst_SboxInst_11_Q2 ;
    wire SubCellInst_SboxInst_11_T0 ;
    wire SubCellInst_SboxInst_11_Q1 ;
    wire SubCellInst_SboxInst_11_Q0 ;
    wire SubCellInst_SboxInst_12_L3 ;
    wire SubCellInst_SboxInst_12_YY_3 ;
    wire SubCellInst_SboxInst_12_L2 ;
    wire SubCellInst_SboxInst_12_T3 ;
    wire SubCellInst_SboxInst_12_Q7 ;
    wire SubCellInst_SboxInst_12_L1 ;
    wire SubCellInst_SboxInst_12_Q6 ;
    wire SubCellInst_SboxInst_12_L0 ;
    wire SubCellInst_SboxInst_12_T2 ;
    wire SubCellInst_SboxInst_12_Q4 ;
    wire SubCellInst_SboxInst_12_T1 ;
    wire SubCellInst_SboxInst_12_Q2 ;
    wire SubCellInst_SboxInst_12_T0 ;
    wire SubCellInst_SboxInst_12_Q1 ;
    wire SubCellInst_SboxInst_12_Q0 ;
    wire SubCellInst_SboxInst_13_L3 ;
    wire SubCellInst_SboxInst_13_YY_3 ;
    wire SubCellInst_SboxInst_13_L2 ;
    wire SubCellInst_SboxInst_13_T3 ;
    wire SubCellInst_SboxInst_13_Q7 ;
    wire SubCellInst_SboxInst_13_L1 ;
    wire SubCellInst_SboxInst_13_Q6 ;
    wire SubCellInst_SboxInst_13_L0 ;
    wire SubCellInst_SboxInst_13_T2 ;
    wire SubCellInst_SboxInst_13_Q4 ;
    wire SubCellInst_SboxInst_13_T1 ;
    wire SubCellInst_SboxInst_13_Q2 ;
    wire SubCellInst_SboxInst_13_T0 ;
    wire SubCellInst_SboxInst_13_Q1 ;
    wire SubCellInst_SboxInst_13_Q0 ;
    wire SubCellInst_SboxInst_14_L3 ;
    wire SubCellInst_SboxInst_14_YY_3 ;
    wire SubCellInst_SboxInst_14_L2 ;
    wire SubCellInst_SboxInst_14_T3 ;
    wire SubCellInst_SboxInst_14_Q7 ;
    wire SubCellInst_SboxInst_14_L1 ;
    wire SubCellInst_SboxInst_14_Q6 ;
    wire SubCellInst_SboxInst_14_L0 ;
    wire SubCellInst_SboxInst_14_T2 ;
    wire SubCellInst_SboxInst_14_Q4 ;
    wire SubCellInst_SboxInst_14_T1 ;
    wire SubCellInst_SboxInst_14_Q2 ;
    wire SubCellInst_SboxInst_14_T0 ;
    wire SubCellInst_SboxInst_14_Q1 ;
    wire SubCellInst_SboxInst_14_Q0 ;
    wire SubCellInst_SboxInst_15_L3 ;
    wire SubCellInst_SboxInst_15_YY_3 ;
    wire SubCellInst_SboxInst_15_L2 ;
    wire SubCellInst_SboxInst_15_T3 ;
    wire SubCellInst_SboxInst_15_Q7 ;
    wire SubCellInst_SboxInst_15_L1 ;
    wire SubCellInst_SboxInst_15_Q6 ;
    wire SubCellInst_SboxInst_15_L0 ;
    wire SubCellInst_SboxInst_15_T2 ;
    wire SubCellInst_SboxInst_15_Q4 ;
    wire SubCellInst_SboxInst_15_T1 ;
    wire SubCellInst_SboxInst_15_Q2 ;
    wire SubCellInst_SboxInst_15_T0 ;
    wire SubCellInst_SboxInst_15_Q1 ;
    wire SubCellInst_SboxInst_15_Q0 ;
    wire MCInst_MCR0_XORInst_0_0_n1 ;
    wire MCInst_MCR0_XORInst_0_1_n1 ;
    wire MCInst_MCR0_XORInst_0_2_n1 ;
    wire MCInst_MCR0_XORInst_0_3_n1 ;
    wire MCInst_MCR0_XORInst_1_0_n1 ;
    wire MCInst_MCR0_XORInst_1_1_n1 ;
    wire MCInst_MCR0_XORInst_1_2_n1 ;
    wire MCInst_MCR0_XORInst_1_3_n1 ;
    wire MCInst_MCR0_XORInst_2_0_n1 ;
    wire MCInst_MCR0_XORInst_2_1_n1 ;
    wire MCInst_MCR0_XORInst_2_2_n1 ;
    wire MCInst_MCR0_XORInst_2_3_n1 ;
    wire MCInst_MCR0_XORInst_3_0_n1 ;
    wire MCInst_MCR0_XORInst_3_1_n1 ;
    wire MCInst_MCR0_XORInst_3_2_n1 ;
    wire MCInst_MCR0_XORInst_3_3_n1 ;
    wire TweakeyGeneration_KEYMUX_MUXInst_0_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_0_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_1_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_1_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_2_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_2_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_3_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_3_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_4_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_4_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_5_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_5_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_6_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_6_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_7_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_7_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_8_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_8_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_9_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_9_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_10_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_10_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_11_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_11_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_12_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_12_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_13_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_13_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_14_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_14_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_15_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_15_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_16_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_16_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_17_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_17_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_18_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_18_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_19_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_19_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_20_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_20_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_21_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_21_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_22_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_22_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_23_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_23_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_24_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_24_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_25_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_25_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_26_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_26_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_27_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_27_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_28_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_28_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_29_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_29_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_30_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_30_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_31_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_31_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_32_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_32_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_33_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_33_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_34_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_34_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_35_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_35_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_36_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_36_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_37_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_37_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_38_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_38_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_39_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_39_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_40_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_40_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_41_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_41_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_42_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_42_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_43_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_43_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_44_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_44_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_45_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_45_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_46_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_46_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_47_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_47_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_48_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_48_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_49_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_49_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_50_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_50_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_51_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_51_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_52_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_52_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_53_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_53_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_54_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_54_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_55_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_55_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_56_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_56_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_57_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_57_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_58_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_58_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_59_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_59_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_60_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_60_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_61_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_61_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_62_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_62_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_63_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_63_U1_X ;
    wire FSMUpdateInst_StateUpdateInst_0_n3 ;
    wire FSMUpdateInst_StateUpdateInst_0_n2 ;
    wire FSMUpdateInst_StateUpdateInst_0_n1 ;
    wire FSMUpdateInst_StateUpdateInst_0_n4 ;
    wire FSMUpdateInst_StateUpdateInst_0_U7_Y ;
    wire FSMUpdateInst_StateUpdateInst_0_U7_X ;
    wire FSMUpdateInst_StateUpdateInst_2_n4 ;
    wire FSMUpdateInst_StateUpdateInst_2_n3 ;
    wire FSMUpdateInst_StateUpdateInst_2_n2 ;
    wire FSMUpdateInst_StateUpdateInst_2_n1 ;
    wire FSMUpdateInst_StateUpdateInst_5_n4 ;
    wire FSMUpdateInst_StateUpdateInst_5_n3 ;
    wire FSMUpdateInst_StateUpdateInst_5_n2 ;
    wire FSMUpdateInst_StateUpdateInst_5_n1 ;
    wire FSMSignalsInst_doneInst_n5 ;
    wire FSMSignalsInst_doneInst_n4 ;
    wire FSMSignalsInst_doneInst_n3 ;
    wire FSMSignalsInst_doneInst_n2 ;
    wire [63:0] MCOutput ;
    wire [61:29] SubCellOutput ;
    wire [5:1] FSM ;
    wire [63:32] AddRoundConstantOutput ;
    wire [47:0] ShiftRowsOutput ;
    wire [5:0] FSMUpdate ;
    wire [1:0] SubCellInst_SboxInst_0_YY ;
    wire [2:1] SubCellInst_SboxInst_0_XX ;
    wire [1:0] SubCellInst_SboxInst_1_YY ;
    wire [2:1] SubCellInst_SboxInst_1_XX ;
    wire [1:0] SubCellInst_SboxInst_2_YY ;
    wire [2:1] SubCellInst_SboxInst_2_XX ;
    wire [1:0] SubCellInst_SboxInst_3_YY ;
    wire [2:1] SubCellInst_SboxInst_3_XX ;
    wire [1:0] SubCellInst_SboxInst_4_YY ;
    wire [2:1] SubCellInst_SboxInst_4_XX ;
    wire [1:0] SubCellInst_SboxInst_5_YY ;
    wire [2:1] SubCellInst_SboxInst_5_XX ;
    wire [1:0] SubCellInst_SboxInst_6_YY ;
    wire [2:1] SubCellInst_SboxInst_6_XX ;
    wire [1:0] SubCellInst_SboxInst_7_YY ;
    wire [2:1] SubCellInst_SboxInst_7_XX ;
    wire [1:0] SubCellInst_SboxInst_8_YY ;
    wire [2:1] SubCellInst_SboxInst_8_XX ;
    wire [1:0] SubCellInst_SboxInst_9_YY ;
    wire [2:1] SubCellInst_SboxInst_9_XX ;
    wire [1:0] SubCellInst_SboxInst_10_YY ;
    wire [2:1] SubCellInst_SboxInst_10_XX ;
    wire [1:0] SubCellInst_SboxInst_11_YY ;
    wire [2:1] SubCellInst_SboxInst_11_XX ;
    wire [1:0] SubCellInst_SboxInst_12_YY ;
    wire [2:1] SubCellInst_SboxInst_12_XX ;
    wire [1:0] SubCellInst_SboxInst_13_YY ;
    wire [2:1] SubCellInst_SboxInst_13_XX ;
    wire [1:0] SubCellInst_SboxInst_14_YY ;
    wire [2:1] SubCellInst_SboxInst_14_XX ;
    wire [1:0] SubCellInst_SboxInst_15_YY ;
    wire [2:1] SubCellInst_SboxInst_15_XX ;
    wire [63:0] TweakeyGeneration_key_Feedback ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;

    /* cells in depth 0 */
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_0_U1_XOR1_U1 ( .A0_t (MCOutput[0]), .A0_f (new_AGEMA_signal_3843), .A1_t (new_AGEMA_signal_3844), .A1_f (new_AGEMA_signal_3845), .B0_t (Plaintext_s0_t[0]), .B0_f (Plaintext_s0_f[0]), .B1_t (Plaintext_s1_t[0]), .B1_f (Plaintext_s1_f[0]), .Z0_t (PlaintextMUX_MUXInst_0_U1_X), .Z0_f (new_AGEMA_signal_3855), .Z1_t (new_AGEMA_signal_3856), .Z1_f (new_AGEMA_signal_3857) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_0_U1_X), .B0_f (new_AGEMA_signal_3855), .B1_t (new_AGEMA_signal_3856), .B1_f (new_AGEMA_signal_3857), .Z0_t (PlaintextMUX_MUXInst_0_U1_Y), .Z0_f (new_AGEMA_signal_3990), .Z1_t (new_AGEMA_signal_3991), .Z1_f (new_AGEMA_signal_3992) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_0_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_0_U1_Y), .A0_f (new_AGEMA_signal_3990), .A1_t (new_AGEMA_signal_3991), .A1_f (new_AGEMA_signal_3992), .B0_t (MCOutput[0]), .B0_f (new_AGEMA_signal_3843), .B1_t (new_AGEMA_signal_3844), .B1_f (new_AGEMA_signal_3845), .Z0_t (Ciphertext_s0_t[0]), .Z0_f (Ciphertext_s0_f[0]), .Z1_t (Ciphertext_s1_t[0]), .Z1_f (Ciphertext_s1_f[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_1_U1_XOR1_U1 ( .A0_t (MCOutput[1]), .A0_f (new_AGEMA_signal_3978), .A1_t (new_AGEMA_signal_3979), .A1_f (new_AGEMA_signal_3980), .B0_t (Plaintext_s0_t[1]), .B0_f (Plaintext_s0_f[1]), .B1_t (Plaintext_s1_t[1]), .B1_f (Plaintext_s1_f[1]), .Z0_t (PlaintextMUX_MUXInst_1_U1_X), .Z0_f (new_AGEMA_signal_3996), .Z1_t (new_AGEMA_signal_3997), .Z1_f (new_AGEMA_signal_3998) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_1_U1_X), .B0_f (new_AGEMA_signal_3996), .B1_t (new_AGEMA_signal_3997), .B1_f (new_AGEMA_signal_3998), .Z0_t (PlaintextMUX_MUXInst_1_U1_Y), .Z0_f (new_AGEMA_signal_4116), .Z1_t (new_AGEMA_signal_4117), .Z1_f (new_AGEMA_signal_4118) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_1_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_1_U1_Y), .A0_f (new_AGEMA_signal_4116), .A1_t (new_AGEMA_signal_4117), .A1_f (new_AGEMA_signal_4118), .B0_t (MCOutput[1]), .B0_f (new_AGEMA_signal_3978), .B1_t (new_AGEMA_signal_3979), .B1_f (new_AGEMA_signal_3980), .Z0_t (Ciphertext_s0_t[1]), .Z0_f (Ciphertext_s0_f[1]), .Z1_t (Ciphertext_s1_t[1]), .Z1_f (Ciphertext_s1_f[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_2_U1_XOR1_U1 ( .A0_t (MCOutput[2]), .A0_f (new_AGEMA_signal_3206), .A1_t (new_AGEMA_signal_3207), .A1_f (new_AGEMA_signal_3208), .B0_t (Plaintext_s0_t[2]), .B0_f (Plaintext_s0_f[2]), .B1_t (Plaintext_s1_t[2]), .B1_f (Plaintext_s1_f[2]), .Z0_t (PlaintextMUX_MUXInst_2_U1_X), .Z0_f (new_AGEMA_signal_3221), .Z1_t (new_AGEMA_signal_3222), .Z1_f (new_AGEMA_signal_3223) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_2_U1_X), .B0_f (new_AGEMA_signal_3221), .B1_t (new_AGEMA_signal_3222), .B1_f (new_AGEMA_signal_3223), .Z0_t (PlaintextMUX_MUXInst_2_U1_Y), .Z0_f (new_AGEMA_signal_3363), .Z1_t (new_AGEMA_signal_3364), .Z1_f (new_AGEMA_signal_3365) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_2_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_2_U1_Y), .A0_f (new_AGEMA_signal_3363), .A1_t (new_AGEMA_signal_3364), .A1_f (new_AGEMA_signal_3365), .B0_t (MCOutput[2]), .B0_f (new_AGEMA_signal_3206), .B1_t (new_AGEMA_signal_3207), .B1_f (new_AGEMA_signal_3208), .Z0_t (Ciphertext_s0_t[2]), .Z0_f (Ciphertext_s0_f[2]), .Z1_t (Ciphertext_s1_t[2]), .Z1_f (Ciphertext_s1_f[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_3_U1_XOR1_U1 ( .A0_t (MCOutput[3]), .A0_f (new_AGEMA_signal_3552), .A1_t (new_AGEMA_signal_3553), .A1_f (new_AGEMA_signal_3554), .B0_t (Plaintext_s0_t[3]), .B0_f (Plaintext_s0_f[3]), .B1_t (Plaintext_s1_t[3]), .B1_f (Plaintext_s1_f[3]), .Z0_t (PlaintextMUX_MUXInst_3_U1_X), .Z0_f (new_AGEMA_signal_3564), .Z1_t (new_AGEMA_signal_3565), .Z1_f (new_AGEMA_signal_3566) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_3_U1_X), .B0_f (new_AGEMA_signal_3564), .B1_t (new_AGEMA_signal_3565), .B1_f (new_AGEMA_signal_3566), .Z0_t (PlaintextMUX_MUXInst_3_U1_Y), .Z0_f (new_AGEMA_signal_3723), .Z1_t (new_AGEMA_signal_3724), .Z1_f (new_AGEMA_signal_3725) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_3_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_3_U1_Y), .A0_f (new_AGEMA_signal_3723), .A1_t (new_AGEMA_signal_3724), .A1_f (new_AGEMA_signal_3725), .B0_t (MCOutput[3]), .B0_f (new_AGEMA_signal_3552), .B1_t (new_AGEMA_signal_3553), .B1_f (new_AGEMA_signal_3554), .Z0_t (Ciphertext_s0_t[3]), .Z0_f (Ciphertext_s0_f[3]), .Z1_t (Ciphertext_s1_t[3]), .Z1_f (Ciphertext_s1_f[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_4_U1_XOR1_U1 ( .A0_t (MCOutput[4]), .A0_f (new_AGEMA_signal_3846), .A1_t (new_AGEMA_signal_3847), .A1_f (new_AGEMA_signal_3848), .B0_t (Plaintext_s0_t[4]), .B0_f (Plaintext_s0_f[4]), .B1_t (Plaintext_s1_t[4]), .B1_f (Plaintext_s1_f[4]), .Z0_t (PlaintextMUX_MUXInst_4_U1_X), .Z0_f (new_AGEMA_signal_3861), .Z1_t (new_AGEMA_signal_3862), .Z1_f (new_AGEMA_signal_3863) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_4_U1_X), .B0_f (new_AGEMA_signal_3861), .B1_t (new_AGEMA_signal_3862), .B1_f (new_AGEMA_signal_3863), .Z0_t (PlaintextMUX_MUXInst_4_U1_Y), .Z0_f (new_AGEMA_signal_3999), .Z1_t (new_AGEMA_signal_4000), .Z1_f (new_AGEMA_signal_4001) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_4_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_4_U1_Y), .A0_f (new_AGEMA_signal_3999), .A1_t (new_AGEMA_signal_4000), .A1_f (new_AGEMA_signal_4001), .B0_t (MCOutput[4]), .B0_f (new_AGEMA_signal_3846), .B1_t (new_AGEMA_signal_3847), .B1_f (new_AGEMA_signal_3848), .Z0_t (Ciphertext_s0_t[4]), .Z0_f (Ciphertext_s0_f[4]), .Z1_t (Ciphertext_s1_t[4]), .Z1_f (Ciphertext_s1_f[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_5_U1_XOR1_U1 ( .A0_t (MCOutput[5]), .A0_f (new_AGEMA_signal_3981), .A1_t (new_AGEMA_signal_3982), .A1_f (new_AGEMA_signal_3983), .B0_t (Plaintext_s0_t[5]), .B0_f (Plaintext_s0_f[5]), .B1_t (Plaintext_s1_t[5]), .B1_f (Plaintext_s1_f[5]), .Z0_t (PlaintextMUX_MUXInst_5_U1_X), .Z0_f (new_AGEMA_signal_4005), .Z1_t (new_AGEMA_signal_4006), .Z1_f (new_AGEMA_signal_4007) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_5_U1_X), .B0_f (new_AGEMA_signal_4005), .B1_t (new_AGEMA_signal_4006), .B1_f (new_AGEMA_signal_4007), .Z0_t (PlaintextMUX_MUXInst_5_U1_Y), .Z0_f (new_AGEMA_signal_4119), .Z1_t (new_AGEMA_signal_4120), .Z1_f (new_AGEMA_signal_4121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_5_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_5_U1_Y), .A0_f (new_AGEMA_signal_4119), .A1_t (new_AGEMA_signal_4120), .A1_f (new_AGEMA_signal_4121), .B0_t (MCOutput[5]), .B0_f (new_AGEMA_signal_3981), .B1_t (new_AGEMA_signal_3982), .B1_f (new_AGEMA_signal_3983), .Z0_t (Ciphertext_s0_t[5]), .Z0_f (Ciphertext_s0_f[5]), .Z1_t (Ciphertext_s1_t[5]), .Z1_f (Ciphertext_s1_f[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_6_U1_XOR1_U1 ( .A0_t (MCOutput[6]), .A0_f (new_AGEMA_signal_3209), .A1_t (new_AGEMA_signal_3210), .A1_f (new_AGEMA_signal_3211), .B0_t (Plaintext_s0_t[6]), .B0_f (Plaintext_s0_f[6]), .B1_t (Plaintext_s1_t[6]), .B1_f (Plaintext_s1_f[6]), .Z0_t (PlaintextMUX_MUXInst_6_U1_X), .Z0_f (new_AGEMA_signal_3227), .Z1_t (new_AGEMA_signal_3228), .Z1_f (new_AGEMA_signal_3229) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_6_U1_X), .B0_f (new_AGEMA_signal_3227), .B1_t (new_AGEMA_signal_3228), .B1_f (new_AGEMA_signal_3229), .Z0_t (PlaintextMUX_MUXInst_6_U1_Y), .Z0_f (new_AGEMA_signal_3366), .Z1_t (new_AGEMA_signal_3367), .Z1_f (new_AGEMA_signal_3368) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_6_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_6_U1_Y), .A0_f (new_AGEMA_signal_3366), .A1_t (new_AGEMA_signal_3367), .A1_f (new_AGEMA_signal_3368), .B0_t (MCOutput[6]), .B0_f (new_AGEMA_signal_3209), .B1_t (new_AGEMA_signal_3210), .B1_f (new_AGEMA_signal_3211), .Z0_t (Ciphertext_s0_t[6]), .Z0_f (Ciphertext_s0_f[6]), .Z1_t (Ciphertext_s1_t[6]), .Z1_f (Ciphertext_s1_f[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_7_U1_XOR1_U1 ( .A0_t (MCOutput[7]), .A0_f (new_AGEMA_signal_3555), .A1_t (new_AGEMA_signal_3556), .A1_f (new_AGEMA_signal_3557), .B0_t (Plaintext_s0_t[7]), .B0_f (Plaintext_s0_f[7]), .B1_t (Plaintext_s1_t[7]), .B1_f (Plaintext_s1_f[7]), .Z0_t (PlaintextMUX_MUXInst_7_U1_X), .Z0_f (new_AGEMA_signal_3570), .Z1_t (new_AGEMA_signal_3571), .Z1_f (new_AGEMA_signal_3572) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_7_U1_X), .B0_f (new_AGEMA_signal_3570), .B1_t (new_AGEMA_signal_3571), .B1_f (new_AGEMA_signal_3572), .Z0_t (PlaintextMUX_MUXInst_7_U1_Y), .Z0_f (new_AGEMA_signal_3726), .Z1_t (new_AGEMA_signal_3727), .Z1_f (new_AGEMA_signal_3728) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_7_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_7_U1_Y), .A0_f (new_AGEMA_signal_3726), .A1_t (new_AGEMA_signal_3727), .A1_f (new_AGEMA_signal_3728), .B0_t (MCOutput[7]), .B0_f (new_AGEMA_signal_3555), .B1_t (new_AGEMA_signal_3556), .B1_f (new_AGEMA_signal_3557), .Z0_t (Ciphertext_s0_t[7]), .Z0_f (Ciphertext_s0_f[7]), .Z1_t (Ciphertext_s1_t[7]), .Z1_f (Ciphertext_s1_f[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_8_U1_XOR1_U1 ( .A0_t (MCOutput[8]), .A0_f (new_AGEMA_signal_3849), .A1_t (new_AGEMA_signal_3850), .A1_f (new_AGEMA_signal_3851), .B0_t (Plaintext_s0_t[8]), .B0_f (Plaintext_s0_f[8]), .B1_t (Plaintext_s1_t[8]), .B1_f (Plaintext_s1_f[8]), .Z0_t (PlaintextMUX_MUXInst_8_U1_X), .Z0_f (new_AGEMA_signal_3867), .Z1_t (new_AGEMA_signal_3868), .Z1_f (new_AGEMA_signal_3869) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_8_U1_X), .B0_f (new_AGEMA_signal_3867), .B1_t (new_AGEMA_signal_3868), .B1_f (new_AGEMA_signal_3869), .Z0_t (PlaintextMUX_MUXInst_8_U1_Y), .Z0_f (new_AGEMA_signal_4008), .Z1_t (new_AGEMA_signal_4009), .Z1_f (new_AGEMA_signal_4010) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_8_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_8_U1_Y), .A0_f (new_AGEMA_signal_4008), .A1_t (new_AGEMA_signal_4009), .A1_f (new_AGEMA_signal_4010), .B0_t (MCOutput[8]), .B0_f (new_AGEMA_signal_3849), .B1_t (new_AGEMA_signal_3850), .B1_f (new_AGEMA_signal_3851), .Z0_t (Ciphertext_s0_t[8]), .Z0_f (Ciphertext_s0_f[8]), .Z1_t (Ciphertext_s1_t[8]), .Z1_f (Ciphertext_s1_f[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_9_U1_XOR1_U1 ( .A0_t (MCOutput[9]), .A0_f (new_AGEMA_signal_3984), .A1_t (new_AGEMA_signal_3985), .A1_f (new_AGEMA_signal_3986), .B0_t (Plaintext_s0_t[9]), .B0_f (Plaintext_s0_f[9]), .B1_t (Plaintext_s1_t[9]), .B1_f (Plaintext_s1_f[9]), .Z0_t (PlaintextMUX_MUXInst_9_U1_X), .Z0_f (new_AGEMA_signal_4014), .Z1_t (new_AGEMA_signal_4015), .Z1_f (new_AGEMA_signal_4016) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_9_U1_X), .B0_f (new_AGEMA_signal_4014), .B1_t (new_AGEMA_signal_4015), .B1_f (new_AGEMA_signal_4016), .Z0_t (PlaintextMUX_MUXInst_9_U1_Y), .Z0_f (new_AGEMA_signal_4122), .Z1_t (new_AGEMA_signal_4123), .Z1_f (new_AGEMA_signal_4124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_9_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_9_U1_Y), .A0_f (new_AGEMA_signal_4122), .A1_t (new_AGEMA_signal_4123), .A1_f (new_AGEMA_signal_4124), .B0_t (MCOutput[9]), .B0_f (new_AGEMA_signal_3984), .B1_t (new_AGEMA_signal_3985), .B1_f (new_AGEMA_signal_3986), .Z0_t (Ciphertext_s0_t[9]), .Z0_f (Ciphertext_s0_f[9]), .Z1_t (Ciphertext_s1_t[9]), .Z1_f (Ciphertext_s1_f[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_10_U1_XOR1_U1 ( .A0_t (MCOutput[10]), .A0_f (new_AGEMA_signal_3212), .A1_t (new_AGEMA_signal_3213), .A1_f (new_AGEMA_signal_3214), .B0_t (Plaintext_s0_t[10]), .B0_f (Plaintext_s0_f[10]), .B1_t (Plaintext_s1_t[10]), .B1_f (Plaintext_s1_f[10]), .Z0_t (PlaintextMUX_MUXInst_10_U1_X), .Z0_f (new_AGEMA_signal_3233), .Z1_t (new_AGEMA_signal_3234), .Z1_f (new_AGEMA_signal_3235) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_10_U1_X), .B0_f (new_AGEMA_signal_3233), .B1_t (new_AGEMA_signal_3234), .B1_f (new_AGEMA_signal_3235), .Z0_t (PlaintextMUX_MUXInst_10_U1_Y), .Z0_f (new_AGEMA_signal_3369), .Z1_t (new_AGEMA_signal_3370), .Z1_f (new_AGEMA_signal_3371) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_10_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_10_U1_Y), .A0_f (new_AGEMA_signal_3369), .A1_t (new_AGEMA_signal_3370), .A1_f (new_AGEMA_signal_3371), .B0_t (MCOutput[10]), .B0_f (new_AGEMA_signal_3212), .B1_t (new_AGEMA_signal_3213), .B1_f (new_AGEMA_signal_3214), .Z0_t (Ciphertext_s0_t[10]), .Z0_f (Ciphertext_s0_f[10]), .Z1_t (Ciphertext_s1_t[10]), .Z1_f (Ciphertext_s1_f[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_11_U1_XOR1_U1 ( .A0_t (MCOutput[11]), .A0_f (new_AGEMA_signal_3558), .A1_t (new_AGEMA_signal_3559), .A1_f (new_AGEMA_signal_3560), .B0_t (Plaintext_s0_t[11]), .B0_f (Plaintext_s0_f[11]), .B1_t (Plaintext_s1_t[11]), .B1_f (Plaintext_s1_f[11]), .Z0_t (PlaintextMUX_MUXInst_11_U1_X), .Z0_f (new_AGEMA_signal_3576), .Z1_t (new_AGEMA_signal_3577), .Z1_f (new_AGEMA_signal_3578) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_11_U1_X), .B0_f (new_AGEMA_signal_3576), .B1_t (new_AGEMA_signal_3577), .B1_f (new_AGEMA_signal_3578), .Z0_t (PlaintextMUX_MUXInst_11_U1_Y), .Z0_f (new_AGEMA_signal_3729), .Z1_t (new_AGEMA_signal_3730), .Z1_f (new_AGEMA_signal_3731) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_11_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_11_U1_Y), .A0_f (new_AGEMA_signal_3729), .A1_t (new_AGEMA_signal_3730), .A1_f (new_AGEMA_signal_3731), .B0_t (MCOutput[11]), .B0_f (new_AGEMA_signal_3558), .B1_t (new_AGEMA_signal_3559), .B1_f (new_AGEMA_signal_3560), .Z0_t (Ciphertext_s0_t[11]), .Z0_f (Ciphertext_s0_f[11]), .Z1_t (Ciphertext_s1_t[11]), .Z1_f (Ciphertext_s1_f[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_12_U1_XOR1_U1 ( .A0_t (MCOutput[12]), .A0_f (new_AGEMA_signal_3987), .A1_t (new_AGEMA_signal_3988), .A1_f (new_AGEMA_signal_3989), .B0_t (Plaintext_s0_t[12]), .B0_f (Plaintext_s0_f[12]), .B1_t (Plaintext_s1_t[12]), .B1_f (Plaintext_s1_f[12]), .Z0_t (PlaintextMUX_MUXInst_12_U1_X), .Z0_f (new_AGEMA_signal_4020), .Z1_t (new_AGEMA_signal_4021), .Z1_f (new_AGEMA_signal_4022) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_12_U1_X), .B0_f (new_AGEMA_signal_4020), .B1_t (new_AGEMA_signal_4021), .B1_f (new_AGEMA_signal_4022), .Z0_t (PlaintextMUX_MUXInst_12_U1_Y), .Z0_f (new_AGEMA_signal_4125), .Z1_t (new_AGEMA_signal_4126), .Z1_f (new_AGEMA_signal_4127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_12_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_12_U1_Y), .A0_f (new_AGEMA_signal_4125), .A1_t (new_AGEMA_signal_4126), .A1_f (new_AGEMA_signal_4127), .B0_t (MCOutput[12]), .B0_f (new_AGEMA_signal_3987), .B1_t (new_AGEMA_signal_3988), .B1_f (new_AGEMA_signal_3989), .Z0_t (Ciphertext_s0_t[12]), .Z0_f (Ciphertext_s0_f[12]), .Z1_t (Ciphertext_s1_t[12]), .Z1_f (Ciphertext_s1_f[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_13_U1_XOR1_U1 ( .A0_t (MCOutput[13]), .A0_f (new_AGEMA_signal_4113), .A1_t (new_AGEMA_signal_4114), .A1_f (new_AGEMA_signal_4115), .B0_t (Plaintext_s0_t[13]), .B0_f (Plaintext_s0_f[13]), .B1_t (Plaintext_s1_t[13]), .B1_f (Plaintext_s1_f[13]), .Z0_t (PlaintextMUX_MUXInst_13_U1_X), .Z0_f (new_AGEMA_signal_4131), .Z1_t (new_AGEMA_signal_4132), .Z1_f (new_AGEMA_signal_4133) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_13_U1_X), .B0_f (new_AGEMA_signal_4131), .B1_t (new_AGEMA_signal_4132), .B1_f (new_AGEMA_signal_4133), .Z0_t (PlaintextMUX_MUXInst_13_U1_Y), .Z0_f (new_AGEMA_signal_4191), .Z1_t (new_AGEMA_signal_4192), .Z1_f (new_AGEMA_signal_4193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_13_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_13_U1_Y), .A0_f (new_AGEMA_signal_4191), .A1_t (new_AGEMA_signal_4192), .A1_f (new_AGEMA_signal_4193), .B0_t (MCOutput[13]), .B0_f (new_AGEMA_signal_4113), .B1_t (new_AGEMA_signal_4114), .B1_f (new_AGEMA_signal_4115), .Z0_t (Ciphertext_s0_t[13]), .Z0_f (Ciphertext_s0_f[13]), .Z1_t (Ciphertext_s1_t[13]), .Z1_f (Ciphertext_s1_f[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_14_U1_XOR1_U1 ( .A0_t (MCOutput[14]), .A0_f (new_AGEMA_signal_3359), .A1_t (new_AGEMA_signal_3360), .A1_f (new_AGEMA_signal_3361), .B0_t (Plaintext_s0_t[14]), .B0_f (Plaintext_s0_f[14]), .B1_t (Plaintext_s1_t[14]), .B1_f (Plaintext_s1_f[14]), .Z0_t (PlaintextMUX_MUXInst_14_U1_X), .Z0_f (new_AGEMA_signal_3375), .Z1_t (new_AGEMA_signal_3376), .Z1_f (new_AGEMA_signal_3377) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_14_U1_X), .B0_f (new_AGEMA_signal_3375), .B1_t (new_AGEMA_signal_3376), .B1_f (new_AGEMA_signal_3377), .Z0_t (PlaintextMUX_MUXInst_14_U1_Y), .Z0_f (new_AGEMA_signal_3579), .Z1_t (new_AGEMA_signal_3580), .Z1_f (new_AGEMA_signal_3581) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_14_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_14_U1_Y), .A0_f (new_AGEMA_signal_3579), .A1_t (new_AGEMA_signal_3580), .A1_f (new_AGEMA_signal_3581), .B0_t (MCOutput[14]), .B0_f (new_AGEMA_signal_3359), .B1_t (new_AGEMA_signal_3360), .B1_f (new_AGEMA_signal_3361), .Z0_t (Ciphertext_s0_t[14]), .Z0_f (Ciphertext_s0_f[14]), .Z1_t (Ciphertext_s1_t[14]), .Z1_f (Ciphertext_s1_f[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_15_U1_XOR1_U1 ( .A0_t (MCOutput[15]), .A0_f (new_AGEMA_signal_3720), .A1_t (new_AGEMA_signal_3721), .A1_f (new_AGEMA_signal_3722), .B0_t (Plaintext_s0_t[15]), .B0_f (Plaintext_s0_f[15]), .B1_t (Plaintext_s1_t[15]), .B1_f (Plaintext_s1_f[15]), .Z0_t (PlaintextMUX_MUXInst_15_U1_X), .Z0_f (new_AGEMA_signal_3735), .Z1_t (new_AGEMA_signal_3736), .Z1_f (new_AGEMA_signal_3737) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_15_U1_X), .B0_f (new_AGEMA_signal_3735), .B1_t (new_AGEMA_signal_3736), .B1_f (new_AGEMA_signal_3737), .Z0_t (PlaintextMUX_MUXInst_15_U1_Y), .Z0_f (new_AGEMA_signal_3870), .Z1_t (new_AGEMA_signal_3871), .Z1_f (new_AGEMA_signal_3872) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_15_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_15_U1_Y), .A0_f (new_AGEMA_signal_3870), .A1_t (new_AGEMA_signal_3871), .A1_f (new_AGEMA_signal_3872), .B0_t (MCOutput[15]), .B0_f (new_AGEMA_signal_3720), .B1_t (new_AGEMA_signal_3721), .B1_f (new_AGEMA_signal_3722), .Z0_t (Ciphertext_s0_t[15]), .Z0_f (Ciphertext_s0_f[15]), .Z1_t (Ciphertext_s1_t[15]), .Z1_f (Ciphertext_s1_f[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_16_U1_XOR1_U1 ( .A0_t (MCOutput[16]), .A0_f (new_AGEMA_signal_3834), .A1_t (new_AGEMA_signal_3835), .A1_f (new_AGEMA_signal_3836), .B0_t (Plaintext_s0_t[16]), .B0_f (Plaintext_s0_f[16]), .B1_t (Plaintext_s1_t[16]), .B1_f (Plaintext_s1_f[16]), .Z0_t (PlaintextMUX_MUXInst_16_U1_X), .Z0_f (new_AGEMA_signal_3876), .Z1_t (new_AGEMA_signal_3877), .Z1_f (new_AGEMA_signal_3878) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_16_U1_X), .B0_f (new_AGEMA_signal_3876), .B1_t (new_AGEMA_signal_3877), .B1_f (new_AGEMA_signal_3878), .Z0_t (PlaintextMUX_MUXInst_16_U1_Y), .Z0_f (new_AGEMA_signal_4023), .Z1_t (new_AGEMA_signal_4024), .Z1_f (new_AGEMA_signal_4025) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_16_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_16_U1_Y), .A0_f (new_AGEMA_signal_4023), .A1_t (new_AGEMA_signal_4024), .A1_f (new_AGEMA_signal_4025), .B0_t (MCOutput[16]), .B0_f (new_AGEMA_signal_3834), .B1_t (new_AGEMA_signal_3835), .B1_f (new_AGEMA_signal_3836), .Z0_t (Ciphertext_s0_t[16]), .Z0_f (Ciphertext_s0_f[16]), .Z1_t (Ciphertext_s1_t[16]), .Z1_f (Ciphertext_s1_f[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_17_U1_XOR1_U1 ( .A0_t (MCOutput[17]), .A0_f (new_AGEMA_signal_3966), .A1_t (new_AGEMA_signal_3967), .A1_f (new_AGEMA_signal_3968), .B0_t (Plaintext_s0_t[17]), .B0_f (Plaintext_s0_f[17]), .B1_t (Plaintext_s1_t[17]), .B1_f (Plaintext_s1_f[17]), .Z0_t (PlaintextMUX_MUXInst_17_U1_X), .Z0_f (new_AGEMA_signal_4029), .Z1_t (new_AGEMA_signal_4030), .Z1_f (new_AGEMA_signal_4031) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_17_U1_X), .B0_f (new_AGEMA_signal_4029), .B1_t (new_AGEMA_signal_4030), .B1_f (new_AGEMA_signal_4031), .Z0_t (PlaintextMUX_MUXInst_17_U1_Y), .Z0_f (new_AGEMA_signal_4134), .Z1_t (new_AGEMA_signal_4135), .Z1_f (new_AGEMA_signal_4136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_17_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_17_U1_Y), .A0_f (new_AGEMA_signal_4134), .A1_t (new_AGEMA_signal_4135), .A1_f (new_AGEMA_signal_4136), .B0_t (MCOutput[17]), .B0_f (new_AGEMA_signal_3966), .B1_t (new_AGEMA_signal_3967), .B1_f (new_AGEMA_signal_3968), .Z0_t (Ciphertext_s0_t[17]), .Z0_f (Ciphertext_s0_f[17]), .Z1_t (Ciphertext_s1_t[17]), .Z1_f (Ciphertext_s1_f[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_18_U1_XOR1_U1 ( .A0_t (MCOutput[18]), .A0_f (new_AGEMA_signal_3194), .A1_t (new_AGEMA_signal_3195), .A1_f (new_AGEMA_signal_3196), .B0_t (Plaintext_s0_t[18]), .B0_f (Plaintext_s0_f[18]), .B1_t (Plaintext_s1_t[18]), .B1_f (Plaintext_s1_f[18]), .Z0_t (PlaintextMUX_MUXInst_18_U1_X), .Z0_f (new_AGEMA_signal_3239), .Z1_t (new_AGEMA_signal_3240), .Z1_f (new_AGEMA_signal_3241) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_18_U1_X), .B0_f (new_AGEMA_signal_3239), .B1_t (new_AGEMA_signal_3240), .B1_f (new_AGEMA_signal_3241), .Z0_t (PlaintextMUX_MUXInst_18_U1_Y), .Z0_f (new_AGEMA_signal_3378), .Z1_t (new_AGEMA_signal_3379), .Z1_f (new_AGEMA_signal_3380) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_18_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_18_U1_Y), .A0_f (new_AGEMA_signal_3378), .A1_t (new_AGEMA_signal_3379), .A1_f (new_AGEMA_signal_3380), .B0_t (MCOutput[18]), .B0_f (new_AGEMA_signal_3194), .B1_t (new_AGEMA_signal_3195), .B1_f (new_AGEMA_signal_3196), .Z0_t (Ciphertext_s0_t[18]), .Z0_f (Ciphertext_s0_f[18]), .Z1_t (Ciphertext_s1_t[18]), .Z1_f (Ciphertext_s1_f[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_19_U1_XOR1_U1 ( .A0_t (MCOutput[19]), .A0_f (new_AGEMA_signal_3540), .A1_t (new_AGEMA_signal_3541), .A1_f (new_AGEMA_signal_3542), .B0_t (Plaintext_s0_t[19]), .B0_f (Plaintext_s0_f[19]), .B1_t (Plaintext_s1_t[19]), .B1_f (Plaintext_s1_f[19]), .Z0_t (PlaintextMUX_MUXInst_19_U1_X), .Z0_f (new_AGEMA_signal_3585), .Z1_t (new_AGEMA_signal_3586), .Z1_f (new_AGEMA_signal_3587) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_19_U1_X), .B0_f (new_AGEMA_signal_3585), .B1_t (new_AGEMA_signal_3586), .B1_f (new_AGEMA_signal_3587), .Z0_t (PlaintextMUX_MUXInst_19_U1_Y), .Z0_f (new_AGEMA_signal_3738), .Z1_t (new_AGEMA_signal_3739), .Z1_f (new_AGEMA_signal_3740) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_19_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_19_U1_Y), .A0_f (new_AGEMA_signal_3738), .A1_t (new_AGEMA_signal_3739), .A1_f (new_AGEMA_signal_3740), .B0_t (MCOutput[19]), .B0_f (new_AGEMA_signal_3540), .B1_t (new_AGEMA_signal_3541), .B1_f (new_AGEMA_signal_3542), .Z0_t (Ciphertext_s0_t[19]), .Z0_f (Ciphertext_s0_f[19]), .Z1_t (Ciphertext_s1_t[19]), .Z1_f (Ciphertext_s1_f[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_20_U1_XOR1_U1 ( .A0_t (MCOutput[20]), .A0_f (new_AGEMA_signal_3837), .A1_t (new_AGEMA_signal_3838), .A1_f (new_AGEMA_signal_3839), .B0_t (Plaintext_s0_t[20]), .B0_f (Plaintext_s0_f[20]), .B1_t (Plaintext_s1_t[20]), .B1_f (Plaintext_s1_f[20]), .Z0_t (PlaintextMUX_MUXInst_20_U1_X), .Z0_f (new_AGEMA_signal_3882), .Z1_t (new_AGEMA_signal_3883), .Z1_f (new_AGEMA_signal_3884) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_20_U1_X), .B0_f (new_AGEMA_signal_3882), .B1_t (new_AGEMA_signal_3883), .B1_f (new_AGEMA_signal_3884), .Z0_t (PlaintextMUX_MUXInst_20_U1_Y), .Z0_f (new_AGEMA_signal_4032), .Z1_t (new_AGEMA_signal_4033), .Z1_f (new_AGEMA_signal_4034) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_20_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_20_U1_Y), .A0_f (new_AGEMA_signal_4032), .A1_t (new_AGEMA_signal_4033), .A1_f (new_AGEMA_signal_4034), .B0_t (MCOutput[20]), .B0_f (new_AGEMA_signal_3837), .B1_t (new_AGEMA_signal_3838), .B1_f (new_AGEMA_signal_3839), .Z0_t (Ciphertext_s0_t[20]), .Z0_f (Ciphertext_s0_f[20]), .Z1_t (Ciphertext_s1_t[20]), .Z1_f (Ciphertext_s1_f[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_21_U1_XOR1_U1 ( .A0_t (MCOutput[21]), .A0_f (new_AGEMA_signal_3969), .A1_t (new_AGEMA_signal_3970), .A1_f (new_AGEMA_signal_3971), .B0_t (Plaintext_s0_t[21]), .B0_f (Plaintext_s0_f[21]), .B1_t (Plaintext_s1_t[21]), .B1_f (Plaintext_s1_f[21]), .Z0_t (PlaintextMUX_MUXInst_21_U1_X), .Z0_f (new_AGEMA_signal_4038), .Z1_t (new_AGEMA_signal_4039), .Z1_f (new_AGEMA_signal_4040) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_21_U1_X), .B0_f (new_AGEMA_signal_4038), .B1_t (new_AGEMA_signal_4039), .B1_f (new_AGEMA_signal_4040), .Z0_t (PlaintextMUX_MUXInst_21_U1_Y), .Z0_f (new_AGEMA_signal_4137), .Z1_t (new_AGEMA_signal_4138), .Z1_f (new_AGEMA_signal_4139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_21_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_21_U1_Y), .A0_f (new_AGEMA_signal_4137), .A1_t (new_AGEMA_signal_4138), .A1_f (new_AGEMA_signal_4139), .B0_t (MCOutput[21]), .B0_f (new_AGEMA_signal_3969), .B1_t (new_AGEMA_signal_3970), .B1_f (new_AGEMA_signal_3971), .Z0_t (Ciphertext_s0_t[21]), .Z0_f (Ciphertext_s0_f[21]), .Z1_t (Ciphertext_s1_t[21]), .Z1_f (Ciphertext_s1_f[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_22_U1_XOR1_U1 ( .A0_t (MCOutput[22]), .A0_f (new_AGEMA_signal_3197), .A1_t (new_AGEMA_signal_3198), .A1_f (new_AGEMA_signal_3199), .B0_t (Plaintext_s0_t[22]), .B0_f (Plaintext_s0_f[22]), .B1_t (Plaintext_s1_t[22]), .B1_f (Plaintext_s1_f[22]), .Z0_t (PlaintextMUX_MUXInst_22_U1_X), .Z0_f (new_AGEMA_signal_3245), .Z1_t (new_AGEMA_signal_3246), .Z1_f (new_AGEMA_signal_3247) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_22_U1_X), .B0_f (new_AGEMA_signal_3245), .B1_t (new_AGEMA_signal_3246), .B1_f (new_AGEMA_signal_3247), .Z0_t (PlaintextMUX_MUXInst_22_U1_Y), .Z0_f (new_AGEMA_signal_3381), .Z1_t (new_AGEMA_signal_3382), .Z1_f (new_AGEMA_signal_3383) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_22_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_22_U1_Y), .A0_f (new_AGEMA_signal_3381), .A1_t (new_AGEMA_signal_3382), .A1_f (new_AGEMA_signal_3383), .B0_t (MCOutput[22]), .B0_f (new_AGEMA_signal_3197), .B1_t (new_AGEMA_signal_3198), .B1_f (new_AGEMA_signal_3199), .Z0_t (Ciphertext_s0_t[22]), .Z0_f (Ciphertext_s0_f[22]), .Z1_t (Ciphertext_s1_t[22]), .Z1_f (Ciphertext_s1_f[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_23_U1_XOR1_U1 ( .A0_t (MCOutput[23]), .A0_f (new_AGEMA_signal_3543), .A1_t (new_AGEMA_signal_3544), .A1_f (new_AGEMA_signal_3545), .B0_t (Plaintext_s0_t[23]), .B0_f (Plaintext_s0_f[23]), .B1_t (Plaintext_s1_t[23]), .B1_f (Plaintext_s1_f[23]), .Z0_t (PlaintextMUX_MUXInst_23_U1_X), .Z0_f (new_AGEMA_signal_3591), .Z1_t (new_AGEMA_signal_3592), .Z1_f (new_AGEMA_signal_3593) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_23_U1_X), .B0_f (new_AGEMA_signal_3591), .B1_t (new_AGEMA_signal_3592), .B1_f (new_AGEMA_signal_3593), .Z0_t (PlaintextMUX_MUXInst_23_U1_Y), .Z0_f (new_AGEMA_signal_3741), .Z1_t (new_AGEMA_signal_3742), .Z1_f (new_AGEMA_signal_3743) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_23_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_23_U1_Y), .A0_f (new_AGEMA_signal_3741), .A1_t (new_AGEMA_signal_3742), .A1_f (new_AGEMA_signal_3743), .B0_t (MCOutput[23]), .B0_f (new_AGEMA_signal_3543), .B1_t (new_AGEMA_signal_3544), .B1_f (new_AGEMA_signal_3545), .Z0_t (Ciphertext_s0_t[23]), .Z0_f (Ciphertext_s0_f[23]), .Z1_t (Ciphertext_s1_t[23]), .Z1_f (Ciphertext_s1_f[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_24_U1_XOR1_U1 ( .A0_t (MCOutput[24]), .A0_f (new_AGEMA_signal_3972), .A1_t (new_AGEMA_signal_3973), .A1_f (new_AGEMA_signal_3974), .B0_t (Plaintext_s0_t[24]), .B0_f (Plaintext_s0_f[24]), .B1_t (Plaintext_s1_t[24]), .B1_f (Plaintext_s1_f[24]), .Z0_t (PlaintextMUX_MUXInst_24_U1_X), .Z0_f (new_AGEMA_signal_4044), .Z1_t (new_AGEMA_signal_4045), .Z1_f (new_AGEMA_signal_4046) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_24_U1_X), .B0_f (new_AGEMA_signal_4044), .B1_t (new_AGEMA_signal_4045), .B1_f (new_AGEMA_signal_4046), .Z0_t (PlaintextMUX_MUXInst_24_U1_Y), .Z0_f (new_AGEMA_signal_4140), .Z1_t (new_AGEMA_signal_4141), .Z1_f (new_AGEMA_signal_4142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_24_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_24_U1_Y), .A0_f (new_AGEMA_signal_4140), .A1_t (new_AGEMA_signal_4141), .A1_f (new_AGEMA_signal_4142), .B0_t (MCOutput[24]), .B0_f (new_AGEMA_signal_3972), .B1_t (new_AGEMA_signal_3973), .B1_f (new_AGEMA_signal_3974), .Z0_t (Ciphertext_s0_t[24]), .Z0_f (Ciphertext_s0_f[24]), .Z1_t (Ciphertext_s1_t[24]), .Z1_f (Ciphertext_s1_f[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_25_U1_XOR1_U1 ( .A0_t (MCOutput[25]), .A0_f (new_AGEMA_signal_4110), .A1_t (new_AGEMA_signal_4111), .A1_f (new_AGEMA_signal_4112), .B0_t (Plaintext_s0_t[25]), .B0_f (Plaintext_s0_f[25]), .B1_t (Plaintext_s1_t[25]), .B1_f (Plaintext_s1_f[25]), .Z0_t (PlaintextMUX_MUXInst_25_U1_X), .Z0_f (new_AGEMA_signal_4146), .Z1_t (new_AGEMA_signal_4147), .Z1_f (new_AGEMA_signal_4148) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_25_U1_X), .B0_f (new_AGEMA_signal_4146), .B1_t (new_AGEMA_signal_4147), .B1_f (new_AGEMA_signal_4148), .Z0_t (PlaintextMUX_MUXInst_25_U1_Y), .Z0_f (new_AGEMA_signal_4194), .Z1_t (new_AGEMA_signal_4195), .Z1_f (new_AGEMA_signal_4196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_25_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_25_U1_Y), .A0_f (new_AGEMA_signal_4194), .A1_t (new_AGEMA_signal_4195), .A1_f (new_AGEMA_signal_4196), .B0_t (MCOutput[25]), .B0_f (new_AGEMA_signal_4110), .B1_t (new_AGEMA_signal_4111), .B1_f (new_AGEMA_signal_4112), .Z0_t (Ciphertext_s0_t[25]), .Z0_f (Ciphertext_s0_f[25]), .Z1_t (Ciphertext_s1_t[25]), .Z1_f (Ciphertext_s1_f[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_26_U1_XOR1_U1 ( .A0_t (MCOutput[26]), .A0_f (new_AGEMA_signal_3200), .A1_t (new_AGEMA_signal_3201), .A1_f (new_AGEMA_signal_3202), .B0_t (Plaintext_s0_t[26]), .B0_f (Plaintext_s0_f[26]), .B1_t (Plaintext_s1_t[26]), .B1_f (Plaintext_s1_f[26]), .Z0_t (PlaintextMUX_MUXInst_26_U1_X), .Z0_f (new_AGEMA_signal_3251), .Z1_t (new_AGEMA_signal_3252), .Z1_f (new_AGEMA_signal_3253) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_26_U1_X), .B0_f (new_AGEMA_signal_3251), .B1_t (new_AGEMA_signal_3252), .B1_f (new_AGEMA_signal_3253), .Z0_t (PlaintextMUX_MUXInst_26_U1_Y), .Z0_f (new_AGEMA_signal_3384), .Z1_t (new_AGEMA_signal_3385), .Z1_f (new_AGEMA_signal_3386) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_26_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_26_U1_Y), .A0_f (new_AGEMA_signal_3384), .A1_t (new_AGEMA_signal_3385), .A1_f (new_AGEMA_signal_3386), .B0_t (MCOutput[26]), .B0_f (new_AGEMA_signal_3200), .B1_t (new_AGEMA_signal_3201), .B1_f (new_AGEMA_signal_3202), .Z0_t (Ciphertext_s0_t[26]), .Z0_f (Ciphertext_s0_f[26]), .Z1_t (Ciphertext_s1_t[26]), .Z1_f (Ciphertext_s1_f[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_27_U1_XOR1_U1 ( .A0_t (MCOutput[27]), .A0_f (new_AGEMA_signal_3546), .A1_t (new_AGEMA_signal_3547), .A1_f (new_AGEMA_signal_3548), .B0_t (Plaintext_s0_t[27]), .B0_f (Plaintext_s0_f[27]), .B1_t (Plaintext_s1_t[27]), .B1_f (Plaintext_s1_f[27]), .Z0_t (PlaintextMUX_MUXInst_27_U1_X), .Z0_f (new_AGEMA_signal_3597), .Z1_t (new_AGEMA_signal_3598), .Z1_f (new_AGEMA_signal_3599) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_27_U1_X), .B0_f (new_AGEMA_signal_3597), .B1_t (new_AGEMA_signal_3598), .B1_f (new_AGEMA_signal_3599), .Z0_t (PlaintextMUX_MUXInst_27_U1_Y), .Z0_f (new_AGEMA_signal_3744), .Z1_t (new_AGEMA_signal_3745), .Z1_f (new_AGEMA_signal_3746) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_27_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_27_U1_Y), .A0_f (new_AGEMA_signal_3744), .A1_t (new_AGEMA_signal_3745), .A1_f (new_AGEMA_signal_3746), .B0_t (MCOutput[27]), .B0_f (new_AGEMA_signal_3546), .B1_t (new_AGEMA_signal_3547), .B1_f (new_AGEMA_signal_3548), .Z0_t (Ciphertext_s0_t[27]), .Z0_f (Ciphertext_s0_f[27]), .Z1_t (Ciphertext_s1_t[27]), .Z1_f (Ciphertext_s1_f[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_28_U1_XOR1_U1 ( .A0_t (MCOutput[28]), .A0_f (new_AGEMA_signal_3840), .A1_t (new_AGEMA_signal_3841), .A1_f (new_AGEMA_signal_3842), .B0_t (Plaintext_s0_t[28]), .B0_f (Plaintext_s0_f[28]), .B1_t (Plaintext_s1_t[28]), .B1_f (Plaintext_s1_f[28]), .Z0_t (PlaintextMUX_MUXInst_28_U1_X), .Z0_f (new_AGEMA_signal_3888), .Z1_t (new_AGEMA_signal_3889), .Z1_f (new_AGEMA_signal_3890) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_28_U1_X), .B0_f (new_AGEMA_signal_3888), .B1_t (new_AGEMA_signal_3889), .B1_f (new_AGEMA_signal_3890), .Z0_t (PlaintextMUX_MUXInst_28_U1_Y), .Z0_f (new_AGEMA_signal_4047), .Z1_t (new_AGEMA_signal_4048), .Z1_f (new_AGEMA_signal_4049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_28_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_28_U1_Y), .A0_f (new_AGEMA_signal_4047), .A1_t (new_AGEMA_signal_4048), .A1_f (new_AGEMA_signal_4049), .B0_t (MCOutput[28]), .B0_f (new_AGEMA_signal_3840), .B1_t (new_AGEMA_signal_3841), .B1_f (new_AGEMA_signal_3842), .Z0_t (Ciphertext_s0_t[28]), .Z0_f (Ciphertext_s0_f[28]), .Z1_t (Ciphertext_s1_t[28]), .Z1_f (Ciphertext_s1_f[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_29_U1_XOR1_U1 ( .A0_t (MCOutput[29]), .A0_f (new_AGEMA_signal_3975), .A1_t (new_AGEMA_signal_3976), .A1_f (new_AGEMA_signal_3977), .B0_t (Plaintext_s0_t[29]), .B0_f (Plaintext_s0_f[29]), .B1_t (Plaintext_s1_t[29]), .B1_f (Plaintext_s1_f[29]), .Z0_t (PlaintextMUX_MUXInst_29_U1_X), .Z0_f (new_AGEMA_signal_4053), .Z1_t (new_AGEMA_signal_4054), .Z1_f (new_AGEMA_signal_4055) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_29_U1_X), .B0_f (new_AGEMA_signal_4053), .B1_t (new_AGEMA_signal_4054), .B1_f (new_AGEMA_signal_4055), .Z0_t (PlaintextMUX_MUXInst_29_U1_Y), .Z0_f (new_AGEMA_signal_4149), .Z1_t (new_AGEMA_signal_4150), .Z1_f (new_AGEMA_signal_4151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_29_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_29_U1_Y), .A0_f (new_AGEMA_signal_4149), .A1_t (new_AGEMA_signal_4150), .A1_f (new_AGEMA_signal_4151), .B0_t (MCOutput[29]), .B0_f (new_AGEMA_signal_3975), .B1_t (new_AGEMA_signal_3976), .B1_f (new_AGEMA_signal_3977), .Z0_t (Ciphertext_s0_t[29]), .Z0_f (Ciphertext_s0_f[29]), .Z1_t (Ciphertext_s1_t[29]), .Z1_f (Ciphertext_s1_f[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_30_U1_XOR1_U1 ( .A0_t (MCOutput[30]), .A0_f (new_AGEMA_signal_3203), .A1_t (new_AGEMA_signal_3204), .A1_f (new_AGEMA_signal_3205), .B0_t (Plaintext_s0_t[30]), .B0_f (Plaintext_s0_f[30]), .B1_t (Plaintext_s1_t[30]), .B1_f (Plaintext_s1_f[30]), .Z0_t (PlaintextMUX_MUXInst_30_U1_X), .Z0_f (new_AGEMA_signal_3257), .Z1_t (new_AGEMA_signal_3258), .Z1_f (new_AGEMA_signal_3259) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_30_U1_X), .B0_f (new_AGEMA_signal_3257), .B1_t (new_AGEMA_signal_3258), .B1_f (new_AGEMA_signal_3259), .Z0_t (PlaintextMUX_MUXInst_30_U1_Y), .Z0_f (new_AGEMA_signal_3387), .Z1_t (new_AGEMA_signal_3388), .Z1_f (new_AGEMA_signal_3389) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_30_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_30_U1_Y), .A0_f (new_AGEMA_signal_3387), .A1_t (new_AGEMA_signal_3388), .A1_f (new_AGEMA_signal_3389), .B0_t (MCOutput[30]), .B0_f (new_AGEMA_signal_3203), .B1_t (new_AGEMA_signal_3204), .B1_f (new_AGEMA_signal_3205), .Z0_t (Ciphertext_s0_t[30]), .Z0_f (Ciphertext_s0_f[30]), .Z1_t (Ciphertext_s1_t[30]), .Z1_f (Ciphertext_s1_f[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_31_U1_XOR1_U1 ( .A0_t (MCOutput[31]), .A0_f (new_AGEMA_signal_3549), .A1_t (new_AGEMA_signal_3550), .A1_f (new_AGEMA_signal_3551), .B0_t (Plaintext_s0_t[31]), .B0_f (Plaintext_s0_f[31]), .B1_t (Plaintext_s1_t[31]), .B1_f (Plaintext_s1_f[31]), .Z0_t (PlaintextMUX_MUXInst_31_U1_X), .Z0_f (new_AGEMA_signal_3603), .Z1_t (new_AGEMA_signal_3604), .Z1_f (new_AGEMA_signal_3605) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_31_U1_X), .B0_f (new_AGEMA_signal_3603), .B1_t (new_AGEMA_signal_3604), .B1_f (new_AGEMA_signal_3605), .Z0_t (PlaintextMUX_MUXInst_31_U1_Y), .Z0_f (new_AGEMA_signal_3747), .Z1_t (new_AGEMA_signal_3748), .Z1_f (new_AGEMA_signal_3749) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_31_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_31_U1_Y), .A0_f (new_AGEMA_signal_3747), .A1_t (new_AGEMA_signal_3748), .A1_f (new_AGEMA_signal_3749), .B0_t (MCOutput[31]), .B0_f (new_AGEMA_signal_3549), .B1_t (new_AGEMA_signal_3550), .B1_f (new_AGEMA_signal_3551), .Z0_t (Ciphertext_s0_t[31]), .Z0_f (Ciphertext_s0_f[31]), .Z1_t (Ciphertext_s1_t[31]), .Z1_f (Ciphertext_s1_f[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_32_U1_XOR1_U1 ( .A0_t (MCOutput[32]), .A0_f (new_AGEMA_signal_3699), .A1_t (new_AGEMA_signal_3700), .A1_f (new_AGEMA_signal_3701), .B0_t (Plaintext_s0_t[32]), .B0_f (Plaintext_s0_f[32]), .B1_t (Plaintext_s1_t[32]), .B1_f (Plaintext_s1_f[32]), .Z0_t (PlaintextMUX_MUXInst_32_U1_X), .Z0_f (new_AGEMA_signal_3753), .Z1_t (new_AGEMA_signal_3754), .Z1_f (new_AGEMA_signal_3755) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_32_U1_X), .B0_f (new_AGEMA_signal_3753), .B1_t (new_AGEMA_signal_3754), .B1_f (new_AGEMA_signal_3755), .Z0_t (PlaintextMUX_MUXInst_32_U1_Y), .Z0_f (new_AGEMA_signal_3891), .Z1_t (new_AGEMA_signal_3892), .Z1_f (new_AGEMA_signal_3893) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_32_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_32_U1_Y), .A0_f (new_AGEMA_signal_3891), .A1_t (new_AGEMA_signal_3892), .A1_f (new_AGEMA_signal_3893), .B0_t (MCOutput[32]), .B0_f (new_AGEMA_signal_3699), .B1_t (new_AGEMA_signal_3700), .B1_f (new_AGEMA_signal_3701), .Z0_t (Ciphertext_s0_t[32]), .Z0_f (Ciphertext_s0_f[32]), .Z1_t (Ciphertext_s1_t[32]), .Z1_f (Ciphertext_s1_f[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_33_U1_XOR1_U1 ( .A0_t (MCOutput[33]), .A0_f (new_AGEMA_signal_3810), .A1_t (new_AGEMA_signal_3811), .A1_f (new_AGEMA_signal_3812), .B0_t (Plaintext_s0_t[33]), .B0_f (Plaintext_s0_f[33]), .B1_t (Plaintext_s1_t[33]), .B1_f (Plaintext_s1_f[33]), .Z0_t (PlaintextMUX_MUXInst_33_U1_X), .Z0_f (new_AGEMA_signal_3897), .Z1_t (new_AGEMA_signal_3898), .Z1_f (new_AGEMA_signal_3899) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_33_U1_X), .B0_f (new_AGEMA_signal_3897), .B1_t (new_AGEMA_signal_3898), .B1_f (new_AGEMA_signal_3899), .Z0_t (PlaintextMUX_MUXInst_33_U1_Y), .Z0_f (new_AGEMA_signal_4056), .Z1_t (new_AGEMA_signal_4057), .Z1_f (new_AGEMA_signal_4058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_33_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_33_U1_Y), .A0_f (new_AGEMA_signal_4056), .A1_t (new_AGEMA_signal_4057), .A1_f (new_AGEMA_signal_4058), .B0_t (MCOutput[33]), .B0_f (new_AGEMA_signal_3810), .B1_t (new_AGEMA_signal_3811), .B1_f (new_AGEMA_signal_3812), .Z0_t (Ciphertext_s0_t[33]), .Z0_f (Ciphertext_s0_f[33]), .Z1_t (Ciphertext_s1_t[33]), .Z1_f (Ciphertext_s1_f[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_34_U1_XOR1_U1 ( .A0_t (MCOutput[34]), .A0_f (new_AGEMA_signal_3008), .A1_t (new_AGEMA_signal_3009), .A1_f (new_AGEMA_signal_3010), .B0_t (Plaintext_s0_t[34]), .B0_f (Plaintext_s0_f[34]), .B1_t (Plaintext_s1_t[34]), .B1_f (Plaintext_s1_f[34]), .Z0_t (PlaintextMUX_MUXInst_34_U1_X), .Z0_f (new_AGEMA_signal_3023), .Z1_t (new_AGEMA_signal_3024), .Z1_f (new_AGEMA_signal_3025) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_34_U1_X), .B0_f (new_AGEMA_signal_3023), .B1_t (new_AGEMA_signal_3024), .B1_f (new_AGEMA_signal_3025), .Z0_t (PlaintextMUX_MUXInst_34_U1_Y), .Z0_f (new_AGEMA_signal_3260), .Z1_t (new_AGEMA_signal_3261), .Z1_f (new_AGEMA_signal_3262) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_34_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_34_U1_Y), .A0_f (new_AGEMA_signal_3260), .A1_t (new_AGEMA_signal_3261), .A1_f (new_AGEMA_signal_3262), .B0_t (MCOutput[34]), .B0_f (new_AGEMA_signal_3008), .B1_t (new_AGEMA_signal_3009), .B1_f (new_AGEMA_signal_3010), .Z0_t (Ciphertext_s0_t[34]), .Z0_f (Ciphertext_s0_f[34]), .Z1_t (Ciphertext_s1_t[34]), .Z1_f (Ciphertext_s1_f[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_35_U1_XOR1_U1 ( .A0_t (MCOutput[35]), .A0_f (new_AGEMA_signal_3338), .A1_t (new_AGEMA_signal_3339), .A1_f (new_AGEMA_signal_3340), .B0_t (Plaintext_s0_t[35]), .B0_f (Plaintext_s0_f[35]), .B1_t (Plaintext_s1_t[35]), .B1_f (Plaintext_s1_f[35]), .Z0_t (PlaintextMUX_MUXInst_35_U1_X), .Z0_f (new_AGEMA_signal_3393), .Z1_t (new_AGEMA_signal_3394), .Z1_f (new_AGEMA_signal_3395) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_35_U1_X), .B0_f (new_AGEMA_signal_3393), .B1_t (new_AGEMA_signal_3394), .B1_f (new_AGEMA_signal_3395), .Z0_t (PlaintextMUX_MUXInst_35_U1_Y), .Z0_f (new_AGEMA_signal_3606), .Z1_t (new_AGEMA_signal_3607), .Z1_f (new_AGEMA_signal_3608) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_35_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_35_U1_Y), .A0_f (new_AGEMA_signal_3606), .A1_t (new_AGEMA_signal_3607), .A1_f (new_AGEMA_signal_3608), .B0_t (MCOutput[35]), .B0_f (new_AGEMA_signal_3338), .B1_t (new_AGEMA_signal_3339), .B1_f (new_AGEMA_signal_3340), .Z0_t (Ciphertext_s0_t[35]), .Z0_f (Ciphertext_s0_f[35]), .Z1_t (Ciphertext_s1_t[35]), .Z1_f (Ciphertext_s1_f[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_36_U1_XOR1_U1 ( .A0_t (MCOutput[36]), .A0_f (new_AGEMA_signal_3702), .A1_t (new_AGEMA_signal_3703), .A1_f (new_AGEMA_signal_3704), .B0_t (Plaintext_s0_t[36]), .B0_f (Plaintext_s0_f[36]), .B1_t (Plaintext_s1_t[36]), .B1_f (Plaintext_s1_f[36]), .Z0_t (PlaintextMUX_MUXInst_36_U1_X), .Z0_f (new_AGEMA_signal_3759), .Z1_t (new_AGEMA_signal_3760), .Z1_f (new_AGEMA_signal_3761) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_36_U1_X), .B0_f (new_AGEMA_signal_3759), .B1_t (new_AGEMA_signal_3760), .B1_f (new_AGEMA_signal_3761), .Z0_t (PlaintextMUX_MUXInst_36_U1_Y), .Z0_f (new_AGEMA_signal_3900), .Z1_t (new_AGEMA_signal_3901), .Z1_f (new_AGEMA_signal_3902) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_36_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_36_U1_Y), .A0_f (new_AGEMA_signal_3900), .A1_t (new_AGEMA_signal_3901), .A1_f (new_AGEMA_signal_3902), .B0_t (MCOutput[36]), .B0_f (new_AGEMA_signal_3702), .B1_t (new_AGEMA_signal_3703), .B1_f (new_AGEMA_signal_3704), .Z0_t (Ciphertext_s0_t[36]), .Z0_f (Ciphertext_s0_f[36]), .Z1_t (Ciphertext_s1_t[36]), .Z1_f (Ciphertext_s1_f[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_37_U1_XOR1_U1 ( .A0_t (MCOutput[37]), .A0_f (new_AGEMA_signal_3813), .A1_t (new_AGEMA_signal_3814), .A1_f (new_AGEMA_signal_3815), .B0_t (Plaintext_s0_t[37]), .B0_f (Plaintext_s0_f[37]), .B1_t (Plaintext_s1_t[37]), .B1_f (Plaintext_s1_f[37]), .Z0_t (PlaintextMUX_MUXInst_37_U1_X), .Z0_f (new_AGEMA_signal_3906), .Z1_t (new_AGEMA_signal_3907), .Z1_f (new_AGEMA_signal_3908) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_37_U1_X), .B0_f (new_AGEMA_signal_3906), .B1_t (new_AGEMA_signal_3907), .B1_f (new_AGEMA_signal_3908), .Z0_t (PlaintextMUX_MUXInst_37_U1_Y), .Z0_f (new_AGEMA_signal_4059), .Z1_t (new_AGEMA_signal_4060), .Z1_f (new_AGEMA_signal_4061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_37_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_37_U1_Y), .A0_f (new_AGEMA_signal_4059), .A1_t (new_AGEMA_signal_4060), .A1_f (new_AGEMA_signal_4061), .B0_t (MCOutput[37]), .B0_f (new_AGEMA_signal_3813), .B1_t (new_AGEMA_signal_3814), .B1_f (new_AGEMA_signal_3815), .Z0_t (Ciphertext_s0_t[37]), .Z0_f (Ciphertext_s0_f[37]), .Z1_t (Ciphertext_s1_t[37]), .Z1_f (Ciphertext_s1_f[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_38_U1_XOR1_U1 ( .A0_t (MCOutput[38]), .A0_f (new_AGEMA_signal_3011), .A1_t (new_AGEMA_signal_3012), .A1_f (new_AGEMA_signal_3013), .B0_t (Plaintext_s0_t[38]), .B0_f (Plaintext_s0_f[38]), .B1_t (Plaintext_s1_t[38]), .B1_f (Plaintext_s1_f[38]), .Z0_t (PlaintextMUX_MUXInst_38_U1_X), .Z0_f (new_AGEMA_signal_3029), .Z1_t (new_AGEMA_signal_3030), .Z1_f (new_AGEMA_signal_3031) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_38_U1_X), .B0_f (new_AGEMA_signal_3029), .B1_t (new_AGEMA_signal_3030), .B1_f (new_AGEMA_signal_3031), .Z0_t (PlaintextMUX_MUXInst_38_U1_Y), .Z0_f (new_AGEMA_signal_3263), .Z1_t (new_AGEMA_signal_3264), .Z1_f (new_AGEMA_signal_3265) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_38_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_38_U1_Y), .A0_f (new_AGEMA_signal_3263), .A1_t (new_AGEMA_signal_3264), .A1_f (new_AGEMA_signal_3265), .B0_t (MCOutput[38]), .B0_f (new_AGEMA_signal_3011), .B1_t (new_AGEMA_signal_3012), .B1_f (new_AGEMA_signal_3013), .Z0_t (Ciphertext_s0_t[38]), .Z0_f (Ciphertext_s0_f[38]), .Z1_t (Ciphertext_s1_t[38]), .Z1_f (Ciphertext_s1_f[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_39_U1_XOR1_U1 ( .A0_t (MCOutput[39]), .A0_f (new_AGEMA_signal_3341), .A1_t (new_AGEMA_signal_3342), .A1_f (new_AGEMA_signal_3343), .B0_t (Plaintext_s0_t[39]), .B0_f (Plaintext_s0_f[39]), .B1_t (Plaintext_s1_t[39]), .B1_f (Plaintext_s1_f[39]), .Z0_t (PlaintextMUX_MUXInst_39_U1_X), .Z0_f (new_AGEMA_signal_3399), .Z1_t (new_AGEMA_signal_3400), .Z1_f (new_AGEMA_signal_3401) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_39_U1_X), .B0_f (new_AGEMA_signal_3399), .B1_t (new_AGEMA_signal_3400), .B1_f (new_AGEMA_signal_3401), .Z0_t (PlaintextMUX_MUXInst_39_U1_Y), .Z0_f (new_AGEMA_signal_3609), .Z1_t (new_AGEMA_signal_3610), .Z1_f (new_AGEMA_signal_3611) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_39_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_39_U1_Y), .A0_f (new_AGEMA_signal_3609), .A1_t (new_AGEMA_signal_3610), .A1_f (new_AGEMA_signal_3611), .B0_t (MCOutput[39]), .B0_f (new_AGEMA_signal_3341), .B1_t (new_AGEMA_signal_3342), .B1_f (new_AGEMA_signal_3343), .Z0_t (Ciphertext_s0_t[39]), .Z0_f (Ciphertext_s0_f[39]), .Z1_t (Ciphertext_s1_t[39]), .Z1_f (Ciphertext_s1_f[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_40_U1_XOR1_U1 ( .A0_t (MCOutput[40]), .A0_f (new_AGEMA_signal_3705), .A1_t (new_AGEMA_signal_3706), .A1_f (new_AGEMA_signal_3707), .B0_t (Plaintext_s0_t[40]), .B0_f (Plaintext_s0_f[40]), .B1_t (Plaintext_s1_t[40]), .B1_f (Plaintext_s1_f[40]), .Z0_t (PlaintextMUX_MUXInst_40_U1_X), .Z0_f (new_AGEMA_signal_3765), .Z1_t (new_AGEMA_signal_3766), .Z1_f (new_AGEMA_signal_3767) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_40_U1_X), .B0_f (new_AGEMA_signal_3765), .B1_t (new_AGEMA_signal_3766), .B1_f (new_AGEMA_signal_3767), .Z0_t (PlaintextMUX_MUXInst_40_U1_Y), .Z0_f (new_AGEMA_signal_3909), .Z1_t (new_AGEMA_signal_3910), .Z1_f (new_AGEMA_signal_3911) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_40_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_40_U1_Y), .A0_f (new_AGEMA_signal_3909), .A1_t (new_AGEMA_signal_3910), .A1_f (new_AGEMA_signal_3911), .B0_t (MCOutput[40]), .B0_f (new_AGEMA_signal_3705), .B1_t (new_AGEMA_signal_3706), .B1_f (new_AGEMA_signal_3707), .Z0_t (Ciphertext_s0_t[40]), .Z0_f (Ciphertext_s0_f[40]), .Z1_t (Ciphertext_s1_t[40]), .Z1_f (Ciphertext_s1_f[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_41_U1_XOR1_U1 ( .A0_t (MCOutput[41]), .A0_f (new_AGEMA_signal_3816), .A1_t (new_AGEMA_signal_3817), .A1_f (new_AGEMA_signal_3818), .B0_t (Plaintext_s0_t[41]), .B0_f (Plaintext_s0_f[41]), .B1_t (Plaintext_s1_t[41]), .B1_f (Plaintext_s1_f[41]), .Z0_t (PlaintextMUX_MUXInst_41_U1_X), .Z0_f (new_AGEMA_signal_3915), .Z1_t (new_AGEMA_signal_3916), .Z1_f (new_AGEMA_signal_3917) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_41_U1_X), .B0_f (new_AGEMA_signal_3915), .B1_t (new_AGEMA_signal_3916), .B1_f (new_AGEMA_signal_3917), .Z0_t (PlaintextMUX_MUXInst_41_U1_Y), .Z0_f (new_AGEMA_signal_4062), .Z1_t (new_AGEMA_signal_4063), .Z1_f (new_AGEMA_signal_4064) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_41_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_41_U1_Y), .A0_f (new_AGEMA_signal_4062), .A1_t (new_AGEMA_signal_4063), .A1_f (new_AGEMA_signal_4064), .B0_t (MCOutput[41]), .B0_f (new_AGEMA_signal_3816), .B1_t (new_AGEMA_signal_3817), .B1_f (new_AGEMA_signal_3818), .Z0_t (Ciphertext_s0_t[41]), .Z0_f (Ciphertext_s0_f[41]), .Z1_t (Ciphertext_s1_t[41]), .Z1_f (Ciphertext_s1_f[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_42_U1_XOR1_U1 ( .A0_t (MCOutput[42]), .A0_f (new_AGEMA_signal_3014), .A1_t (new_AGEMA_signal_3015), .A1_f (new_AGEMA_signal_3016), .B0_t (Plaintext_s0_t[42]), .B0_f (Plaintext_s0_f[42]), .B1_t (Plaintext_s1_t[42]), .B1_f (Plaintext_s1_f[42]), .Z0_t (PlaintextMUX_MUXInst_42_U1_X), .Z0_f (new_AGEMA_signal_3035), .Z1_t (new_AGEMA_signal_3036), .Z1_f (new_AGEMA_signal_3037) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_42_U1_X), .B0_f (new_AGEMA_signal_3035), .B1_t (new_AGEMA_signal_3036), .B1_f (new_AGEMA_signal_3037), .Z0_t (PlaintextMUX_MUXInst_42_U1_Y), .Z0_f (new_AGEMA_signal_3266), .Z1_t (new_AGEMA_signal_3267), .Z1_f (new_AGEMA_signal_3268) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_42_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_42_U1_Y), .A0_f (new_AGEMA_signal_3266), .A1_t (new_AGEMA_signal_3267), .A1_f (new_AGEMA_signal_3268), .B0_t (MCOutput[42]), .B0_f (new_AGEMA_signal_3014), .B1_t (new_AGEMA_signal_3015), .B1_f (new_AGEMA_signal_3016), .Z0_t (Ciphertext_s0_t[42]), .Z0_f (Ciphertext_s0_f[42]), .Z1_t (Ciphertext_s1_t[42]), .Z1_f (Ciphertext_s1_f[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_43_U1_XOR1_U1 ( .A0_t (MCOutput[43]), .A0_f (new_AGEMA_signal_3344), .A1_t (new_AGEMA_signal_3345), .A1_f (new_AGEMA_signal_3346), .B0_t (Plaintext_s0_t[43]), .B0_f (Plaintext_s0_f[43]), .B1_t (Plaintext_s1_t[43]), .B1_f (Plaintext_s1_f[43]), .Z0_t (PlaintextMUX_MUXInst_43_U1_X), .Z0_f (new_AGEMA_signal_3405), .Z1_t (new_AGEMA_signal_3406), .Z1_f (new_AGEMA_signal_3407) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_43_U1_X), .B0_f (new_AGEMA_signal_3405), .B1_t (new_AGEMA_signal_3406), .B1_f (new_AGEMA_signal_3407), .Z0_t (PlaintextMUX_MUXInst_43_U1_Y), .Z0_f (new_AGEMA_signal_3612), .Z1_t (new_AGEMA_signal_3613), .Z1_f (new_AGEMA_signal_3614) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_43_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_43_U1_Y), .A0_f (new_AGEMA_signal_3612), .A1_t (new_AGEMA_signal_3613), .A1_f (new_AGEMA_signal_3614), .B0_t (MCOutput[43]), .B0_f (new_AGEMA_signal_3344), .B1_t (new_AGEMA_signal_3345), .B1_f (new_AGEMA_signal_3346), .Z0_t (Ciphertext_s0_t[43]), .Z0_f (Ciphertext_s0_f[43]), .Z1_t (Ciphertext_s1_t[43]), .Z1_f (Ciphertext_s1_f[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_44_U1_XOR1_U1 ( .A0_t (MCOutput[44]), .A0_f (new_AGEMA_signal_3819), .A1_t (new_AGEMA_signal_3820), .A1_f (new_AGEMA_signal_3821), .B0_t (Plaintext_s0_t[44]), .B0_f (Plaintext_s0_f[44]), .B1_t (Plaintext_s1_t[44]), .B1_f (Plaintext_s1_f[44]), .Z0_t (PlaintextMUX_MUXInst_44_U1_X), .Z0_f (new_AGEMA_signal_3921), .Z1_t (new_AGEMA_signal_3922), .Z1_f (new_AGEMA_signal_3923) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_44_U1_X), .B0_f (new_AGEMA_signal_3921), .B1_t (new_AGEMA_signal_3922), .B1_f (new_AGEMA_signal_3923), .Z0_t (PlaintextMUX_MUXInst_44_U1_Y), .Z0_f (new_AGEMA_signal_4065), .Z1_t (new_AGEMA_signal_4066), .Z1_f (new_AGEMA_signal_4067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_44_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_44_U1_Y), .A0_f (new_AGEMA_signal_4065), .A1_t (new_AGEMA_signal_4066), .A1_f (new_AGEMA_signal_4067), .B0_t (MCOutput[44]), .B0_f (new_AGEMA_signal_3819), .B1_t (new_AGEMA_signal_3820), .B1_f (new_AGEMA_signal_3821), .Z0_t (Ciphertext_s0_t[44]), .Z0_f (Ciphertext_s0_f[44]), .Z1_t (Ciphertext_s1_t[44]), .Z1_f (Ciphertext_s1_f[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_45_U1_XOR1_U1 ( .A0_t (MCOutput[45]), .A0_f (new_AGEMA_signal_3942), .A1_t (new_AGEMA_signal_3943), .A1_f (new_AGEMA_signal_3944), .B0_t (Plaintext_s0_t[45]), .B0_f (Plaintext_s0_f[45]), .B1_t (Plaintext_s1_t[45]), .B1_f (Plaintext_s1_f[45]), .Z0_t (PlaintextMUX_MUXInst_45_U1_X), .Z0_f (new_AGEMA_signal_4071), .Z1_t (new_AGEMA_signal_4072), .Z1_f (new_AGEMA_signal_4073) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_45_U1_X), .B0_f (new_AGEMA_signal_4071), .B1_t (new_AGEMA_signal_4072), .B1_f (new_AGEMA_signal_4073), .Z0_t (PlaintextMUX_MUXInst_45_U1_Y), .Z0_f (new_AGEMA_signal_4152), .Z1_t (new_AGEMA_signal_4153), .Z1_f (new_AGEMA_signal_4154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_45_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_45_U1_Y), .A0_f (new_AGEMA_signal_4152), .A1_t (new_AGEMA_signal_4153), .A1_f (new_AGEMA_signal_4154), .B0_t (MCOutput[45]), .B0_f (new_AGEMA_signal_3942), .B1_t (new_AGEMA_signal_3943), .B1_f (new_AGEMA_signal_3944), .Z0_t (Ciphertext_s0_t[45]), .Z0_f (Ciphertext_s0_f[45]), .Z1_t (Ciphertext_s1_t[45]), .Z1_f (Ciphertext_s1_f[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_46_U1_XOR1_U1 ( .A0_t (MCOutput[46]), .A0_f (new_AGEMA_signal_3182), .A1_t (new_AGEMA_signal_3183), .A1_f (new_AGEMA_signal_3184), .B0_t (Plaintext_s0_t[46]), .B0_f (Plaintext_s0_f[46]), .B1_t (Plaintext_s1_t[46]), .B1_f (Plaintext_s1_f[46]), .Z0_t (PlaintextMUX_MUXInst_46_U1_X), .Z0_f (new_AGEMA_signal_3272), .Z1_t (new_AGEMA_signal_3273), .Z1_f (new_AGEMA_signal_3274) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_46_U1_X), .B0_f (new_AGEMA_signal_3272), .B1_t (new_AGEMA_signal_3273), .B1_f (new_AGEMA_signal_3274), .Z0_t (PlaintextMUX_MUXInst_46_U1_Y), .Z0_f (new_AGEMA_signal_3408), .Z1_t (new_AGEMA_signal_3409), .Z1_f (new_AGEMA_signal_3410) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_46_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_46_U1_Y), .A0_f (new_AGEMA_signal_3408), .A1_t (new_AGEMA_signal_3409), .A1_f (new_AGEMA_signal_3410), .B0_t (MCOutput[46]), .B0_f (new_AGEMA_signal_3182), .B1_t (new_AGEMA_signal_3183), .B1_f (new_AGEMA_signal_3184), .Z0_t (Ciphertext_s0_t[46]), .Z0_f (Ciphertext_s0_f[46]), .Z1_t (Ciphertext_s1_t[46]), .Z1_f (Ciphertext_s1_f[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_47_U1_XOR1_U1 ( .A0_t (MCOutput[47]), .A0_f (new_AGEMA_signal_3525), .A1_t (new_AGEMA_signal_3526), .A1_f (new_AGEMA_signal_3527), .B0_t (Plaintext_s0_t[47]), .B0_f (Plaintext_s0_f[47]), .B1_t (Plaintext_s1_t[47]), .B1_f (Plaintext_s1_f[47]), .Z0_t (PlaintextMUX_MUXInst_47_U1_X), .Z0_f (new_AGEMA_signal_3618), .Z1_t (new_AGEMA_signal_3619), .Z1_f (new_AGEMA_signal_3620) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_47_U1_X), .B0_f (new_AGEMA_signal_3618), .B1_t (new_AGEMA_signal_3619), .B1_f (new_AGEMA_signal_3620), .Z0_t (PlaintextMUX_MUXInst_47_U1_Y), .Z0_f (new_AGEMA_signal_3768), .Z1_t (new_AGEMA_signal_3769), .Z1_f (new_AGEMA_signal_3770) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_47_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_47_U1_Y), .A0_f (new_AGEMA_signal_3768), .A1_t (new_AGEMA_signal_3769), .A1_f (new_AGEMA_signal_3770), .B0_t (MCOutput[47]), .B0_f (new_AGEMA_signal_3525), .B1_t (new_AGEMA_signal_3526), .B1_f (new_AGEMA_signal_3527), .Z0_t (Ciphertext_s0_t[47]), .Z0_f (Ciphertext_s0_f[47]), .Z1_t (Ciphertext_s1_t[47]), .Z1_f (Ciphertext_s1_f[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_48_U1_XOR1_U1 ( .A0_t (MCOutput[48]), .A0_f (new_AGEMA_signal_3945), .A1_t (new_AGEMA_signal_3946), .A1_f (new_AGEMA_signal_3947), .B0_t (Plaintext_s0_t[48]), .B0_f (Plaintext_s0_f[48]), .B1_t (Plaintext_s1_t[48]), .B1_f (Plaintext_s1_f[48]), .Z0_t (PlaintextMUX_MUXInst_48_U1_X), .Z0_f (new_AGEMA_signal_4077), .Z1_t (new_AGEMA_signal_4078), .Z1_f (new_AGEMA_signal_4079) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_48_U1_X), .B0_f (new_AGEMA_signal_4077), .B1_t (new_AGEMA_signal_4078), .B1_f (new_AGEMA_signal_4079), .Z0_t (PlaintextMUX_MUXInst_48_U1_Y), .Z0_f (new_AGEMA_signal_4155), .Z1_t (new_AGEMA_signal_4156), .Z1_f (new_AGEMA_signal_4157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_48_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_48_U1_Y), .A0_f (new_AGEMA_signal_4155), .A1_t (new_AGEMA_signal_4156), .A1_f (new_AGEMA_signal_4157), .B0_t (MCOutput[48]), .B0_f (new_AGEMA_signal_3945), .B1_t (new_AGEMA_signal_3946), .B1_f (new_AGEMA_signal_3947), .Z0_t (Ciphertext_s0_t[48]), .Z0_f (Ciphertext_s0_f[48]), .Z1_t (Ciphertext_s1_t[48]), .Z1_f (Ciphertext_s1_f[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_49_U1_XOR1_U1 ( .A0_t (MCOutput[49]), .A0_f (new_AGEMA_signal_4095), .A1_t (new_AGEMA_signal_4096), .A1_f (new_AGEMA_signal_4097), .B0_t (Plaintext_s0_t[49]), .B0_f (Plaintext_s0_f[49]), .B1_t (Plaintext_s1_t[49]), .B1_f (Plaintext_s1_f[49]), .Z0_t (PlaintextMUX_MUXInst_49_U1_X), .Z0_f (new_AGEMA_signal_4161), .Z1_t (new_AGEMA_signal_4162), .Z1_f (new_AGEMA_signal_4163) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_49_U1_X), .B0_f (new_AGEMA_signal_4161), .B1_t (new_AGEMA_signal_4162), .B1_f (new_AGEMA_signal_4163), .Z0_t (PlaintextMUX_MUXInst_49_U1_Y), .Z0_f (new_AGEMA_signal_4197), .Z1_t (new_AGEMA_signal_4198), .Z1_f (new_AGEMA_signal_4199) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_49_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_49_U1_Y), .A0_f (new_AGEMA_signal_4197), .A1_t (new_AGEMA_signal_4198), .A1_f (new_AGEMA_signal_4199), .B0_t (MCOutput[49]), .B0_f (new_AGEMA_signal_4095), .B1_t (new_AGEMA_signal_4096), .B1_f (new_AGEMA_signal_4097), .Z0_t (Ciphertext_s0_t[49]), .Z0_f (Ciphertext_s0_f[49]), .Z1_t (Ciphertext_s1_t[49]), .Z1_f (Ciphertext_s1_f[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_50_U1_XOR1_U1 ( .A0_t (MCOutput[50]), .A0_f (new_AGEMA_signal_3347), .A1_t (new_AGEMA_signal_3348), .A1_f (new_AGEMA_signal_3349), .B0_t (Plaintext_s0_t[50]), .B0_f (Plaintext_s0_f[50]), .B1_t (Plaintext_s1_t[50]), .B1_f (Plaintext_s1_f[50]), .Z0_t (PlaintextMUX_MUXInst_50_U1_X), .Z0_f (new_AGEMA_signal_3414), .Z1_t (new_AGEMA_signal_3415), .Z1_f (new_AGEMA_signal_3416) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_50_U1_X), .B0_f (new_AGEMA_signal_3414), .B1_t (new_AGEMA_signal_3415), .B1_f (new_AGEMA_signal_3416), .Z0_t (PlaintextMUX_MUXInst_50_U1_Y), .Z0_f (new_AGEMA_signal_3621), .Z1_t (new_AGEMA_signal_3622), .Z1_f (new_AGEMA_signal_3623) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_50_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_50_U1_Y), .A0_f (new_AGEMA_signal_3621), .A1_t (new_AGEMA_signal_3622), .A1_f (new_AGEMA_signal_3623), .B0_t (MCOutput[50]), .B0_f (new_AGEMA_signal_3347), .B1_t (new_AGEMA_signal_3348), .B1_f (new_AGEMA_signal_3349), .Z0_t (Ciphertext_s0_t[50]), .Z0_f (Ciphertext_s0_f[50]), .Z1_t (Ciphertext_s1_t[50]), .Z1_f (Ciphertext_s1_f[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_51_U1_XOR1_U1 ( .A0_t (MCOutput[51]), .A0_f (new_AGEMA_signal_3708), .A1_t (new_AGEMA_signal_3709), .A1_f (new_AGEMA_signal_3710), .B0_t (Plaintext_s0_t[51]), .B0_f (Plaintext_s0_f[51]), .B1_t (Plaintext_s1_t[51]), .B1_f (Plaintext_s1_f[51]), .Z0_t (PlaintextMUX_MUXInst_51_U1_X), .Z0_f (new_AGEMA_signal_3774), .Z1_t (new_AGEMA_signal_3775), .Z1_f (new_AGEMA_signal_3776) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_51_U1_X), .B0_f (new_AGEMA_signal_3774), .B1_t (new_AGEMA_signal_3775), .B1_f (new_AGEMA_signal_3776), .Z0_t (PlaintextMUX_MUXInst_51_U1_Y), .Z0_f (new_AGEMA_signal_3924), .Z1_t (new_AGEMA_signal_3925), .Z1_f (new_AGEMA_signal_3926) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_51_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_51_U1_Y), .A0_f (new_AGEMA_signal_3924), .A1_t (new_AGEMA_signal_3925), .A1_f (new_AGEMA_signal_3926), .B0_t (MCOutput[51]), .B0_f (new_AGEMA_signal_3708), .B1_t (new_AGEMA_signal_3709), .B1_f (new_AGEMA_signal_3710), .Z0_t (Ciphertext_s0_t[51]), .Z0_f (Ciphertext_s0_f[51]), .Z1_t (Ciphertext_s1_t[51]), .Z1_f (Ciphertext_s1_f[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_52_U1_XOR1_U1 ( .A0_t (MCOutput[52]), .A0_f (new_AGEMA_signal_3951), .A1_t (new_AGEMA_signal_3952), .A1_f (new_AGEMA_signal_3953), .B0_t (Plaintext_s0_t[52]), .B0_f (Plaintext_s0_f[52]), .B1_t (Plaintext_s1_t[52]), .B1_f (Plaintext_s1_f[52]), .Z0_t (PlaintextMUX_MUXInst_52_U1_X), .Z0_f (new_AGEMA_signal_4083), .Z1_t (new_AGEMA_signal_4084), .Z1_f (new_AGEMA_signal_4085) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_52_U1_X), .B0_f (new_AGEMA_signal_4083), .B1_t (new_AGEMA_signal_4084), .B1_f (new_AGEMA_signal_4085), .Z0_t (PlaintextMUX_MUXInst_52_U1_Y), .Z0_f (new_AGEMA_signal_4164), .Z1_t (new_AGEMA_signal_4165), .Z1_f (new_AGEMA_signal_4166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_52_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_52_U1_Y), .A0_f (new_AGEMA_signal_4164), .A1_t (new_AGEMA_signal_4165), .A1_f (new_AGEMA_signal_4166), .B0_t (MCOutput[52]), .B0_f (new_AGEMA_signal_3951), .B1_t (new_AGEMA_signal_3952), .B1_f (new_AGEMA_signal_3953), .Z0_t (Ciphertext_s0_t[52]), .Z0_f (Ciphertext_s0_f[52]), .Z1_t (Ciphertext_s1_t[52]), .Z1_f (Ciphertext_s1_f[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_53_U1_XOR1_U1 ( .A0_t (MCOutput[53]), .A0_f (new_AGEMA_signal_4098), .A1_t (new_AGEMA_signal_4099), .A1_f (new_AGEMA_signal_4100), .B0_t (Plaintext_s0_t[53]), .B0_f (Plaintext_s0_f[53]), .B1_t (Plaintext_s1_t[53]), .B1_f (Plaintext_s1_f[53]), .Z0_t (PlaintextMUX_MUXInst_53_U1_X), .Z0_f (new_AGEMA_signal_4170), .Z1_t (new_AGEMA_signal_4171), .Z1_f (new_AGEMA_signal_4172) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_53_U1_X), .B0_f (new_AGEMA_signal_4170), .B1_t (new_AGEMA_signal_4171), .B1_f (new_AGEMA_signal_4172), .Z0_t (PlaintextMUX_MUXInst_53_U1_Y), .Z0_f (new_AGEMA_signal_4200), .Z1_t (new_AGEMA_signal_4201), .Z1_f (new_AGEMA_signal_4202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_53_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_53_U1_Y), .A0_f (new_AGEMA_signal_4200), .A1_t (new_AGEMA_signal_4201), .A1_f (new_AGEMA_signal_4202), .B0_t (MCOutput[53]), .B0_f (new_AGEMA_signal_4098), .B1_t (new_AGEMA_signal_4099), .B1_f (new_AGEMA_signal_4100), .Z0_t (Ciphertext_s0_t[53]), .Z0_f (Ciphertext_s0_f[53]), .Z1_t (Ciphertext_s1_t[53]), .Z1_f (Ciphertext_s1_f[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_54_U1_XOR1_U1 ( .A0_t (MCOutput[54]), .A0_f (new_AGEMA_signal_3350), .A1_t (new_AGEMA_signal_3351), .A1_f (new_AGEMA_signal_3352), .B0_t (Plaintext_s0_t[54]), .B0_f (Plaintext_s0_f[54]), .B1_t (Plaintext_s1_t[54]), .B1_f (Plaintext_s1_f[54]), .Z0_t (PlaintextMUX_MUXInst_54_U1_X), .Z0_f (new_AGEMA_signal_3420), .Z1_t (new_AGEMA_signal_3421), .Z1_f (new_AGEMA_signal_3422) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_54_U1_X), .B0_f (new_AGEMA_signal_3420), .B1_t (new_AGEMA_signal_3421), .B1_f (new_AGEMA_signal_3422), .Z0_t (PlaintextMUX_MUXInst_54_U1_Y), .Z0_f (new_AGEMA_signal_3624), .Z1_t (new_AGEMA_signal_3625), .Z1_f (new_AGEMA_signal_3626) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_54_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_54_U1_Y), .A0_f (new_AGEMA_signal_3624), .A1_t (new_AGEMA_signal_3625), .A1_f (new_AGEMA_signal_3626), .B0_t (MCOutput[54]), .B0_f (new_AGEMA_signal_3350), .B1_t (new_AGEMA_signal_3351), .B1_f (new_AGEMA_signal_3352), .Z0_t (Ciphertext_s0_t[54]), .Z0_f (Ciphertext_s0_f[54]), .Z1_t (Ciphertext_s1_t[54]), .Z1_f (Ciphertext_s1_f[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_55_U1_XOR1_U1 ( .A0_t (MCOutput[55]), .A0_f (new_AGEMA_signal_3711), .A1_t (new_AGEMA_signal_3712), .A1_f (new_AGEMA_signal_3713), .B0_t (Plaintext_s0_t[55]), .B0_f (Plaintext_s0_f[55]), .B1_t (Plaintext_s1_t[55]), .B1_f (Plaintext_s1_f[55]), .Z0_t (PlaintextMUX_MUXInst_55_U1_X), .Z0_f (new_AGEMA_signal_3780), .Z1_t (new_AGEMA_signal_3781), .Z1_f (new_AGEMA_signal_3782) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_55_U1_X), .B0_f (new_AGEMA_signal_3780), .B1_t (new_AGEMA_signal_3781), .B1_f (new_AGEMA_signal_3782), .Z0_t (PlaintextMUX_MUXInst_55_U1_Y), .Z0_f (new_AGEMA_signal_3927), .Z1_t (new_AGEMA_signal_3928), .Z1_f (new_AGEMA_signal_3929) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_55_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_55_U1_Y), .A0_f (new_AGEMA_signal_3927), .A1_t (new_AGEMA_signal_3928), .A1_f (new_AGEMA_signal_3929), .B0_t (MCOutput[55]), .B0_f (new_AGEMA_signal_3711), .B1_t (new_AGEMA_signal_3712), .B1_f (new_AGEMA_signal_3713), .Z0_t (Ciphertext_s0_t[55]), .Z0_f (Ciphertext_s0_f[55]), .Z1_t (Ciphertext_s1_t[55]), .Z1_f (Ciphertext_s1_f[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_56_U1_XOR1_U1 ( .A0_t (MCOutput[56]), .A0_f (new_AGEMA_signal_3957), .A1_t (new_AGEMA_signal_3958), .A1_f (new_AGEMA_signal_3959), .B0_t (Plaintext_s0_t[56]), .B0_f (Plaintext_s0_f[56]), .B1_t (Plaintext_s1_t[56]), .B1_f (Plaintext_s1_f[56]), .Z0_t (PlaintextMUX_MUXInst_56_U1_X), .Z0_f (new_AGEMA_signal_4089), .Z1_t (new_AGEMA_signal_4090), .Z1_f (new_AGEMA_signal_4091) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_56_U1_X), .B0_f (new_AGEMA_signal_4089), .B1_t (new_AGEMA_signal_4090), .B1_f (new_AGEMA_signal_4091), .Z0_t (PlaintextMUX_MUXInst_56_U1_Y), .Z0_f (new_AGEMA_signal_4173), .Z1_t (new_AGEMA_signal_4174), .Z1_f (new_AGEMA_signal_4175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_56_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_56_U1_Y), .A0_f (new_AGEMA_signal_4173), .A1_t (new_AGEMA_signal_4174), .A1_f (new_AGEMA_signal_4175), .B0_t (MCOutput[56]), .B0_f (new_AGEMA_signal_3957), .B1_t (new_AGEMA_signal_3958), .B1_f (new_AGEMA_signal_3959), .Z0_t (Ciphertext_s0_t[56]), .Z0_f (Ciphertext_s0_f[56]), .Z1_t (Ciphertext_s1_t[56]), .Z1_f (Ciphertext_s1_f[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_57_U1_XOR1_U1 ( .A0_t (MCOutput[57]), .A0_f (new_AGEMA_signal_4101), .A1_t (new_AGEMA_signal_4102), .A1_f (new_AGEMA_signal_4103), .B0_t (Plaintext_s0_t[57]), .B0_f (Plaintext_s0_f[57]), .B1_t (Plaintext_s1_t[57]), .B1_f (Plaintext_s1_f[57]), .Z0_t (PlaintextMUX_MUXInst_57_U1_X), .Z0_f (new_AGEMA_signal_4179), .Z1_t (new_AGEMA_signal_4180), .Z1_f (new_AGEMA_signal_4181) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_57_U1_X), .B0_f (new_AGEMA_signal_4179), .B1_t (new_AGEMA_signal_4180), .B1_f (new_AGEMA_signal_4181), .Z0_t (PlaintextMUX_MUXInst_57_U1_Y), .Z0_f (new_AGEMA_signal_4203), .Z1_t (new_AGEMA_signal_4204), .Z1_f (new_AGEMA_signal_4205) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_57_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_57_U1_Y), .A0_f (new_AGEMA_signal_4203), .A1_t (new_AGEMA_signal_4204), .A1_f (new_AGEMA_signal_4205), .B0_t (MCOutput[57]), .B0_f (new_AGEMA_signal_4101), .B1_t (new_AGEMA_signal_4102), .B1_f (new_AGEMA_signal_4103), .Z0_t (Ciphertext_s0_t[57]), .Z0_f (Ciphertext_s0_f[57]), .Z1_t (Ciphertext_s1_t[57]), .Z1_f (Ciphertext_s1_f[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_58_U1_XOR1_U1 ( .A0_t (MCOutput[58]), .A0_f (new_AGEMA_signal_3353), .A1_t (new_AGEMA_signal_3354), .A1_f (new_AGEMA_signal_3355), .B0_t (Plaintext_s0_t[58]), .B0_f (Plaintext_s0_f[58]), .B1_t (Plaintext_s1_t[58]), .B1_f (Plaintext_s1_f[58]), .Z0_t (PlaintextMUX_MUXInst_58_U1_X), .Z0_f (new_AGEMA_signal_3426), .Z1_t (new_AGEMA_signal_3427), .Z1_f (new_AGEMA_signal_3428) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_58_U1_X), .B0_f (new_AGEMA_signal_3426), .B1_t (new_AGEMA_signal_3427), .B1_f (new_AGEMA_signal_3428), .Z0_t (PlaintextMUX_MUXInst_58_U1_Y), .Z0_f (new_AGEMA_signal_3627), .Z1_t (new_AGEMA_signal_3628), .Z1_f (new_AGEMA_signal_3629) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_58_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_58_U1_Y), .A0_f (new_AGEMA_signal_3627), .A1_t (new_AGEMA_signal_3628), .A1_f (new_AGEMA_signal_3629), .B0_t (MCOutput[58]), .B0_f (new_AGEMA_signal_3353), .B1_t (new_AGEMA_signal_3354), .B1_f (new_AGEMA_signal_3355), .Z0_t (Ciphertext_s0_t[58]), .Z0_f (Ciphertext_s0_f[58]), .Z1_t (Ciphertext_s1_t[58]), .Z1_f (Ciphertext_s1_f[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_59_U1_XOR1_U1 ( .A0_t (MCOutput[59]), .A0_f (new_AGEMA_signal_3714), .A1_t (new_AGEMA_signal_3715), .A1_f (new_AGEMA_signal_3716), .B0_t (Plaintext_s0_t[59]), .B0_f (Plaintext_s0_f[59]), .B1_t (Plaintext_s1_t[59]), .B1_f (Plaintext_s1_f[59]), .Z0_t (PlaintextMUX_MUXInst_59_U1_X), .Z0_f (new_AGEMA_signal_3786), .Z1_t (new_AGEMA_signal_3787), .Z1_f (new_AGEMA_signal_3788) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_59_U1_X), .B0_f (new_AGEMA_signal_3786), .B1_t (new_AGEMA_signal_3787), .B1_f (new_AGEMA_signal_3788), .Z0_t (PlaintextMUX_MUXInst_59_U1_Y), .Z0_f (new_AGEMA_signal_3930), .Z1_t (new_AGEMA_signal_3931), .Z1_f (new_AGEMA_signal_3932) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_59_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_59_U1_Y), .A0_f (new_AGEMA_signal_3930), .A1_t (new_AGEMA_signal_3931), .A1_f (new_AGEMA_signal_3932), .B0_t (MCOutput[59]), .B0_f (new_AGEMA_signal_3714), .B1_t (new_AGEMA_signal_3715), .B1_f (new_AGEMA_signal_3716), .Z0_t (Ciphertext_s0_t[59]), .Z0_f (Ciphertext_s0_f[59]), .Z1_t (Ciphertext_s1_t[59]), .Z1_f (Ciphertext_s1_f[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_60_U1_XOR1_U1 ( .A0_t (MCOutput[60]), .A0_f (new_AGEMA_signal_4104), .A1_t (new_AGEMA_signal_4105), .A1_f (new_AGEMA_signal_4106), .B0_t (Plaintext_s0_t[60]), .B0_f (Plaintext_s0_f[60]), .B1_t (Plaintext_s1_t[60]), .B1_f (Plaintext_s1_f[60]), .Z0_t (PlaintextMUX_MUXInst_60_U1_X), .Z0_f (new_AGEMA_signal_4185), .Z1_t (new_AGEMA_signal_4186), .Z1_f (new_AGEMA_signal_4187) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_60_U1_X), .B0_f (new_AGEMA_signal_4185), .B1_t (new_AGEMA_signal_4186), .B1_f (new_AGEMA_signal_4187), .Z0_t (PlaintextMUX_MUXInst_60_U1_Y), .Z0_f (new_AGEMA_signal_4206), .Z1_t (new_AGEMA_signal_4207), .Z1_f (new_AGEMA_signal_4208) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_60_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_60_U1_Y), .A0_f (new_AGEMA_signal_4206), .A1_t (new_AGEMA_signal_4207), .A1_f (new_AGEMA_signal_4208), .B0_t (MCOutput[60]), .B0_f (new_AGEMA_signal_4104), .B1_t (new_AGEMA_signal_4105), .B1_f (new_AGEMA_signal_4106), .Z0_t (Ciphertext_s0_t[60]), .Z0_f (Ciphertext_s0_f[60]), .Z1_t (Ciphertext_s1_t[60]), .Z1_f (Ciphertext_s1_f[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_61_U1_XOR1_U1 ( .A0_t (MCOutput[61]), .A0_f (new_AGEMA_signal_4188), .A1_t (new_AGEMA_signal_4189), .A1_f (new_AGEMA_signal_4190), .B0_t (Plaintext_s0_t[61]), .B0_f (Plaintext_s0_f[61]), .B1_t (Plaintext_s1_t[61]), .B1_f (Plaintext_s1_f[61]), .Z0_t (PlaintextMUX_MUXInst_61_U1_X), .Z0_f (new_AGEMA_signal_4212), .Z1_t (new_AGEMA_signal_4213), .Z1_f (new_AGEMA_signal_4214) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_61_U1_X), .B0_f (new_AGEMA_signal_4212), .B1_t (new_AGEMA_signal_4213), .B1_f (new_AGEMA_signal_4214), .Z0_t (PlaintextMUX_MUXInst_61_U1_Y), .Z0_f (new_AGEMA_signal_4215), .Z1_t (new_AGEMA_signal_4216), .Z1_f (new_AGEMA_signal_4217) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_61_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_61_U1_Y), .A0_f (new_AGEMA_signal_4215), .A1_t (new_AGEMA_signal_4216), .A1_f (new_AGEMA_signal_4217), .B0_t (MCOutput[61]), .B0_f (new_AGEMA_signal_4188), .B1_t (new_AGEMA_signal_4189), .B1_f (new_AGEMA_signal_4190), .Z0_t (Ciphertext_s0_t[61]), .Z0_f (Ciphertext_s0_f[61]), .Z1_t (Ciphertext_s1_t[61]), .Z1_f (Ciphertext_s1_f[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_62_U1_XOR1_U1 ( .A0_t (MCOutput[62]), .A0_f (new_AGEMA_signal_3537), .A1_t (new_AGEMA_signal_3538), .A1_f (new_AGEMA_signal_3539), .B0_t (Plaintext_s0_t[62]), .B0_f (Plaintext_s0_f[62]), .B1_t (Plaintext_s1_t[62]), .B1_f (Plaintext_s1_f[62]), .Z0_t (PlaintextMUX_MUXInst_62_U1_X), .Z0_f (new_AGEMA_signal_3633), .Z1_t (new_AGEMA_signal_3634), .Z1_f (new_AGEMA_signal_3635) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_62_U1_X), .B0_f (new_AGEMA_signal_3633), .B1_t (new_AGEMA_signal_3634), .B1_f (new_AGEMA_signal_3635), .Z0_t (PlaintextMUX_MUXInst_62_U1_Y), .Z0_f (new_AGEMA_signal_3789), .Z1_t (new_AGEMA_signal_3790), .Z1_f (new_AGEMA_signal_3791) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_62_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_62_U1_Y), .A0_f (new_AGEMA_signal_3789), .A1_t (new_AGEMA_signal_3790), .A1_f (new_AGEMA_signal_3791), .B0_t (MCOutput[62]), .B0_f (new_AGEMA_signal_3537), .B1_t (new_AGEMA_signal_3538), .B1_f (new_AGEMA_signal_3539), .Z0_t (Ciphertext_s0_t[62]), .Z0_f (Ciphertext_s0_f[62]), .Z1_t (Ciphertext_s1_t[62]), .Z1_f (Ciphertext_s1_f[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_63_U1_XOR1_U1 ( .A0_t (MCOutput[63]), .A0_f (new_AGEMA_signal_3831), .A1_t (new_AGEMA_signal_3832), .A1_f (new_AGEMA_signal_3833), .B0_t (Plaintext_s0_t[63]), .B0_f (Plaintext_s0_f[63]), .B1_t (Plaintext_s1_t[63]), .B1_f (Plaintext_s1_f[63]), .Z0_t (PlaintextMUX_MUXInst_63_U1_X), .Z0_f (new_AGEMA_signal_3936), .Z1_t (new_AGEMA_signal_3937), .Z1_f (new_AGEMA_signal_3938) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (PlaintextMUX_MUXInst_63_U1_X), .B0_f (new_AGEMA_signal_3936), .B1_t (new_AGEMA_signal_3937), .B1_f (new_AGEMA_signal_3938), .Z0_t (PlaintextMUX_MUXInst_63_U1_Y), .Z0_f (new_AGEMA_signal_4092), .Z1_t (new_AGEMA_signal_4093), .Z1_f (new_AGEMA_signal_4094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_63_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_63_U1_Y), .A0_f (new_AGEMA_signal_4092), .A1_t (new_AGEMA_signal_4093), .A1_f (new_AGEMA_signal_4094), .B0_t (MCOutput[63]), .B0_f (new_AGEMA_signal_3831), .B1_t (new_AGEMA_signal_3832), .B1_f (new_AGEMA_signal_3833), .Z0_t (Ciphertext_s0_t[63]), .Z0_f (Ciphertext_s0_f[63]), .Z1_t (Ciphertext_s1_t[63]), .Z1_f (Ciphertext_s1_f[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[2]), .A0_f (Ciphertext_s0_f[2]), .A1_t (Ciphertext_s1_t[2]), .A1_f (Ciphertext_s1_f[2]), .B0_t (Ciphertext_s0_t[3]), .B0_f (Ciphertext_s0_f[3]), .B1_t (Ciphertext_s1_t[3]), .B1_f (Ciphertext_s1_f[3]), .Z0_t (SubCellInst_SboxInst_0_XX[1]), .Z0_f (new_AGEMA_signal_1345), .Z1_t (new_AGEMA_signal_1346), .Z1_f (new_AGEMA_signal_1347) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[0]), .A0_f (Ciphertext_s0_f[0]), .A1_t (Ciphertext_s1_t[0]), .A1_f (Ciphertext_s1_f[0]), .B0_t (Ciphertext_s0_t[2]), .B0_f (Ciphertext_s0_f[2]), .B1_t (Ciphertext_s1_t[2]), .B1_f (Ciphertext_s1_f[2]), .Z0_t (SubCellInst_SboxInst_0_XX[2]), .Z0_f (new_AGEMA_signal_1351), .Z1_t (new_AGEMA_signal_1352), .Z1_f (new_AGEMA_signal_1353) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR0_U1 ( .A0_t (Ciphertext_s0_t[1]), .A0_f (Ciphertext_s0_f[1]), .A1_t (Ciphertext_s1_t[1]), .A1_f (Ciphertext_s1_f[1]), .B0_t (SubCellInst_SboxInst_0_XX[2]), .B0_f (new_AGEMA_signal_1351), .B1_t (new_AGEMA_signal_1352), .B1_f (new_AGEMA_signal_1353), .Z0_t (SubCellInst_SboxInst_0_Q0), .Z0_f (new_AGEMA_signal_2313), .Z1_t (new_AGEMA_signal_2314), .Z1_f (new_AGEMA_signal_2315) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR1_U1 ( .A0_t (Ciphertext_s0_t[1]), .A0_f (Ciphertext_s0_f[1]), .A1_t (Ciphertext_s1_t[1]), .A1_f (Ciphertext_s1_f[1]), .B0_t (SubCellInst_SboxInst_0_XX[1]), .B0_f (new_AGEMA_signal_1345), .B1_t (new_AGEMA_signal_1346), .B1_f (new_AGEMA_signal_1347), .Z0_t (SubCellInst_SboxInst_0_Q1), .Z0_f (new_AGEMA_signal_2316), .Z1_t (new_AGEMA_signal_2317), .Z1_f (new_AGEMA_signal_2318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_AND1_U1 ( .A0_t (Ciphertext_s0_t[2]), .A0_f (Ciphertext_s0_f[2]), .A1_t (Ciphertext_s1_t[2]), .A1_f (Ciphertext_s1_f[2]), .B0_t (SubCellInst_SboxInst_0_Q1), .B0_f (new_AGEMA_signal_2316), .B1_t (new_AGEMA_signal_2317), .B1_f (new_AGEMA_signal_2318), .Z0_t (SubCellInst_SboxInst_0_T0), .Z0_f (new_AGEMA_signal_2701), .Z1_t (new_AGEMA_signal_2702), .Z1_f (new_AGEMA_signal_2703) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_0_Q0), .A0_f (new_AGEMA_signal_2313), .A1_t (new_AGEMA_signal_2314), .A1_f (new_AGEMA_signal_2315), .B0_t (SubCellInst_SboxInst_0_T0), .B0_f (new_AGEMA_signal_2701), .B1_t (new_AGEMA_signal_2702), .B1_f (new_AGEMA_signal_2703), .Z0_t (SubCellInst_SboxInst_0_Q2), .Z0_f (new_AGEMA_signal_2849), .Z1_t (new_AGEMA_signal_2850), .Z1_f (new_AGEMA_signal_2851) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_AND2_U1 ( .A0_t (Ciphertext_s0_t[1]), .A0_f (Ciphertext_s0_f[1]), .A1_t (Ciphertext_s1_t[1]), .A1_f (Ciphertext_s1_f[1]), .B0_t (SubCellInst_SboxInst_0_Q2), .B0_f (new_AGEMA_signal_2849), .B1_t (new_AGEMA_signal_2850), .B1_f (new_AGEMA_signal_2851), .Z0_t (SubCellInst_SboxInst_0_T1), .Z0_f (new_AGEMA_signal_3038), .Z1_t (new_AGEMA_signal_3039), .Z1_f (new_AGEMA_signal_3040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_XOR3_U1 ( .A0_t (Ciphertext_s0_t[1]), .A0_f (Ciphertext_s0_f[1]), .A1_t (Ciphertext_s1_t[1]), .A1_f (Ciphertext_s1_f[1]), .B0_t (Ciphertext_s0_t[2]), .B0_f (Ciphertext_s0_f[2]), .B1_t (Ciphertext_s1_t[2]), .B1_f (Ciphertext_s1_f[2]), .Z0_t (SubCellInst_SboxInst_0_Q4), .Z0_f (new_AGEMA_signal_1357), .Z1_t (new_AGEMA_signal_1358), .Z1_f (new_AGEMA_signal_1359) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_AND3_U1 ( .A0_t (Ciphertext_s0_t[2]), .A0_f (Ciphertext_s0_f[2]), .A1_t (Ciphertext_s1_t[2]), .A1_f (Ciphertext_s1_f[2]), .B0_t (SubCellInst_SboxInst_0_Q4), .B0_f (new_AGEMA_signal_1357), .B1_t (new_AGEMA_signal_1358), .B1_f (new_AGEMA_signal_1359), .Z0_t (SubCellInst_SboxInst_0_T2), .Z0_f (new_AGEMA_signal_2319), .Z1_t (new_AGEMA_signal_2320), .Z1_f (new_AGEMA_signal_2321) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_0_T1), .A0_f (new_AGEMA_signal_3038), .A1_t (new_AGEMA_signal_3039), .A1_f (new_AGEMA_signal_3040), .B0_t (SubCellInst_SboxInst_0_T2), .B0_f (new_AGEMA_signal_2319), .B1_t (new_AGEMA_signal_2320), .B1_f (new_AGEMA_signal_2321), .Z0_t (SubCellInst_SboxInst_0_L0), .Z0_f (new_AGEMA_signal_3275), .Z1_t (new_AGEMA_signal_3276), .Z1_f (new_AGEMA_signal_3277) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_0_XX[2]), .A0_f (new_AGEMA_signal_1351), .A1_t (new_AGEMA_signal_1352), .A1_f (new_AGEMA_signal_1353), .B0_t (Ciphertext_s0_t[2]), .B0_f (Ciphertext_s0_f[2]), .B1_t (Ciphertext_s1_t[2]), .B1_f (Ciphertext_s1_f[2]), .Z0_t (SubCellInst_SboxInst_0_Q6), .Z0_f (new_AGEMA_signal_2322), .Z1_t (new_AGEMA_signal_2323), .Z1_f (new_AGEMA_signal_2324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_0_Q1), .A0_f (new_AGEMA_signal_2316), .A1_t (new_AGEMA_signal_2317), .A1_f (new_AGEMA_signal_2318), .B0_t (SubCellInst_SboxInst_0_Q6), .B0_f (new_AGEMA_signal_2322), .B1_t (new_AGEMA_signal_2323), .B1_f (new_AGEMA_signal_2324), .Z0_t (SubCellInst_SboxInst_0_L1), .Z0_f (new_AGEMA_signal_2704), .Z1_t (new_AGEMA_signal_2705), .Z1_f (new_AGEMA_signal_2706) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_0_L1), .A0_f (new_AGEMA_signal_2704), .A1_t (new_AGEMA_signal_2705), .A1_f (new_AGEMA_signal_2706), .B0_t (SubCellInst_SboxInst_0_T2), .B0_f (new_AGEMA_signal_2319), .B1_t (new_AGEMA_signal_2320), .B1_f (new_AGEMA_signal_2321), .Z0_t (SubCellInst_SboxInst_0_Q7), .Z0_f (new_AGEMA_signal_2852), .Z1_t (new_AGEMA_signal_2853), .Z1_f (new_AGEMA_signal_2854) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_AND4_U1 ( .A0_t (SubCellInst_SboxInst_0_Q6), .A0_f (new_AGEMA_signal_2322), .A1_t (new_AGEMA_signal_2323), .A1_f (new_AGEMA_signal_2324), .B0_t (SubCellInst_SboxInst_0_Q7), .B0_f (new_AGEMA_signal_2852), .B1_t (new_AGEMA_signal_2853), .B1_f (new_AGEMA_signal_2854), .Z0_t (SubCellInst_SboxInst_0_T3), .Z0_f (new_AGEMA_signal_3041), .Z1_t (new_AGEMA_signal_3042), .Z1_f (new_AGEMA_signal_3043) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR8_U1 ( .A0_t (Ciphertext_s0_t[1]), .A0_f (Ciphertext_s0_f[1]), .A1_t (Ciphertext_s1_t[1]), .A1_f (Ciphertext_s1_f[1]), .B0_t (Ciphertext_s0_t[2]), .B0_f (Ciphertext_s0_f[2]), .B1_t (Ciphertext_s1_t[2]), .B1_f (Ciphertext_s1_f[2]), .Z0_t (SubCellInst_SboxInst_0_L2), .Z0_f (new_AGEMA_signal_1360), .Z1_t (new_AGEMA_signal_1361), .Z1_f (new_AGEMA_signal_1362) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_0_L0), .A0_f (new_AGEMA_signal_3275), .A1_t (new_AGEMA_signal_3276), .A1_f (new_AGEMA_signal_3277), .B0_t (SubCellInst_SboxInst_0_L2), .B0_f (new_AGEMA_signal_1360), .B1_t (new_AGEMA_signal_1361), .B1_f (new_AGEMA_signal_1362), .Z0_t (SubCellInst_SboxInst_0_YY_3), .Z0_f (new_AGEMA_signal_3429), .Z1_t (new_AGEMA_signal_3430), .Z1_f (new_AGEMA_signal_3431) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_0_L0), .A0_f (new_AGEMA_signal_3275), .A1_t (new_AGEMA_signal_3276), .A1_f (new_AGEMA_signal_3277), .B0_t (SubCellInst_SboxInst_0_T3), .B0_f (new_AGEMA_signal_3041), .B1_t (new_AGEMA_signal_3042), .B1_f (new_AGEMA_signal_3043), .Z0_t (ShiftRowsOutput[4]), .Z0_f (new_AGEMA_signal_3432), .Z1_t (new_AGEMA_signal_3433), .Z1_f (new_AGEMA_signal_3434) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_0_XX[2]), .A0_f (new_AGEMA_signal_1351), .A1_t (new_AGEMA_signal_1352), .A1_f (new_AGEMA_signal_1353), .B0_t (SubCellInst_SboxInst_0_T0), .B0_f (new_AGEMA_signal_2701), .B1_t (new_AGEMA_signal_2702), .B1_f (new_AGEMA_signal_2703), .Z0_t (SubCellInst_SboxInst_0_L3), .Z0_f (new_AGEMA_signal_2855), .Z1_t (new_AGEMA_signal_2856), .Z1_f (new_AGEMA_signal_2857) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_0_L3), .A0_f (new_AGEMA_signal_2855), .A1_t (new_AGEMA_signal_2856), .A1_f (new_AGEMA_signal_2857), .B0_t (SubCellInst_SboxInst_0_T2), .B0_f (new_AGEMA_signal_2319), .B1_t (new_AGEMA_signal_2320), .B1_f (new_AGEMA_signal_2321), .Z0_t (SubCellInst_SboxInst_0_YY[1]), .Z0_f (new_AGEMA_signal_3044), .Z1_t (new_AGEMA_signal_3045), .Z1_f (new_AGEMA_signal_3046) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_0_XX[1]), .A0_f (new_AGEMA_signal_1345), .A1_t (new_AGEMA_signal_1346), .A1_f (new_AGEMA_signal_1347), .B0_t (SubCellInst_SboxInst_0_T2), .B0_f (new_AGEMA_signal_2319), .B1_t (new_AGEMA_signal_2320), .B1_f (new_AGEMA_signal_2321), .Z0_t (SubCellInst_SboxInst_0_YY[0]), .Z0_f (new_AGEMA_signal_2707), .Z1_t (new_AGEMA_signal_2708), .Z1_f (new_AGEMA_signal_2709) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_0_YY[1]), .A0_f (new_AGEMA_signal_3044), .A1_t (new_AGEMA_signal_3045), .A1_f (new_AGEMA_signal_3046), .B0_t (SubCellInst_SboxInst_0_YY_3), .B0_f (new_AGEMA_signal_3429), .B1_t (new_AGEMA_signal_3430), .B1_f (new_AGEMA_signal_3431), .Z0_t (ShiftRowsOutput[5]), .Z0_f (new_AGEMA_signal_3636), .Z1_t (new_AGEMA_signal_3637), .Z1_f (new_AGEMA_signal_3638) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[6]), .A0_f (Ciphertext_s0_f[6]), .A1_t (Ciphertext_s1_t[6]), .A1_f (Ciphertext_s1_f[6]), .B0_t (Ciphertext_s0_t[7]), .B0_f (Ciphertext_s0_f[7]), .B1_t (Ciphertext_s1_t[7]), .B1_f (Ciphertext_s1_f[7]), .Z0_t (SubCellInst_SboxInst_1_XX[1]), .Z0_f (new_AGEMA_signal_1369), .Z1_t (new_AGEMA_signal_1370), .Z1_f (new_AGEMA_signal_1371) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[4]), .A0_f (Ciphertext_s0_f[4]), .A1_t (Ciphertext_s1_t[4]), .A1_f (Ciphertext_s1_f[4]), .B0_t (Ciphertext_s0_t[6]), .B0_f (Ciphertext_s0_f[6]), .B1_t (Ciphertext_s1_t[6]), .B1_f (Ciphertext_s1_f[6]), .Z0_t (SubCellInst_SboxInst_1_XX[2]), .Z0_f (new_AGEMA_signal_1375), .Z1_t (new_AGEMA_signal_1376), .Z1_f (new_AGEMA_signal_1377) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR0_U1 ( .A0_t (Ciphertext_s0_t[5]), .A0_f (Ciphertext_s0_f[5]), .A1_t (Ciphertext_s1_t[5]), .A1_f (Ciphertext_s1_f[5]), .B0_t (SubCellInst_SboxInst_1_XX[2]), .B0_f (new_AGEMA_signal_1375), .B1_t (new_AGEMA_signal_1376), .B1_f (new_AGEMA_signal_1377), .Z0_t (SubCellInst_SboxInst_1_Q0), .Z0_f (new_AGEMA_signal_2325), .Z1_t (new_AGEMA_signal_2326), .Z1_f (new_AGEMA_signal_2327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR1_U1 ( .A0_t (Ciphertext_s0_t[5]), .A0_f (Ciphertext_s0_f[5]), .A1_t (Ciphertext_s1_t[5]), .A1_f (Ciphertext_s1_f[5]), .B0_t (SubCellInst_SboxInst_1_XX[1]), .B0_f (new_AGEMA_signal_1369), .B1_t (new_AGEMA_signal_1370), .B1_f (new_AGEMA_signal_1371), .Z0_t (SubCellInst_SboxInst_1_Q1), .Z0_f (new_AGEMA_signal_2328), .Z1_t (new_AGEMA_signal_2329), .Z1_f (new_AGEMA_signal_2330) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_AND1_U1 ( .A0_t (Ciphertext_s0_t[6]), .A0_f (Ciphertext_s0_f[6]), .A1_t (Ciphertext_s1_t[6]), .A1_f (Ciphertext_s1_f[6]), .B0_t (SubCellInst_SboxInst_1_Q1), .B0_f (new_AGEMA_signal_2328), .B1_t (new_AGEMA_signal_2329), .B1_f (new_AGEMA_signal_2330), .Z0_t (SubCellInst_SboxInst_1_T0), .Z0_f (new_AGEMA_signal_2710), .Z1_t (new_AGEMA_signal_2711), .Z1_f (new_AGEMA_signal_2712) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_1_Q0), .A0_f (new_AGEMA_signal_2325), .A1_t (new_AGEMA_signal_2326), .A1_f (new_AGEMA_signal_2327), .B0_t (SubCellInst_SboxInst_1_T0), .B0_f (new_AGEMA_signal_2710), .B1_t (new_AGEMA_signal_2711), .B1_f (new_AGEMA_signal_2712), .Z0_t (SubCellInst_SboxInst_1_Q2), .Z0_f (new_AGEMA_signal_2858), .Z1_t (new_AGEMA_signal_2859), .Z1_f (new_AGEMA_signal_2860) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_AND2_U1 ( .A0_t (Ciphertext_s0_t[5]), .A0_f (Ciphertext_s0_f[5]), .A1_t (Ciphertext_s1_t[5]), .A1_f (Ciphertext_s1_f[5]), .B0_t (SubCellInst_SboxInst_1_Q2), .B0_f (new_AGEMA_signal_2858), .B1_t (new_AGEMA_signal_2859), .B1_f (new_AGEMA_signal_2860), .Z0_t (SubCellInst_SboxInst_1_T1), .Z0_f (new_AGEMA_signal_3047), .Z1_t (new_AGEMA_signal_3048), .Z1_f (new_AGEMA_signal_3049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_XOR3_U1 ( .A0_t (Ciphertext_s0_t[5]), .A0_f (Ciphertext_s0_f[5]), .A1_t (Ciphertext_s1_t[5]), .A1_f (Ciphertext_s1_f[5]), .B0_t (Ciphertext_s0_t[6]), .B0_f (Ciphertext_s0_f[6]), .B1_t (Ciphertext_s1_t[6]), .B1_f (Ciphertext_s1_f[6]), .Z0_t (SubCellInst_SboxInst_1_Q4), .Z0_f (new_AGEMA_signal_1381), .Z1_t (new_AGEMA_signal_1382), .Z1_f (new_AGEMA_signal_1383) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_AND3_U1 ( .A0_t (Ciphertext_s0_t[6]), .A0_f (Ciphertext_s0_f[6]), .A1_t (Ciphertext_s1_t[6]), .A1_f (Ciphertext_s1_f[6]), .B0_t (SubCellInst_SboxInst_1_Q4), .B0_f (new_AGEMA_signal_1381), .B1_t (new_AGEMA_signal_1382), .B1_f (new_AGEMA_signal_1383), .Z0_t (SubCellInst_SboxInst_1_T2), .Z0_f (new_AGEMA_signal_2331), .Z1_t (new_AGEMA_signal_2332), .Z1_f (new_AGEMA_signal_2333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_1_T1), .A0_f (new_AGEMA_signal_3047), .A1_t (new_AGEMA_signal_3048), .A1_f (new_AGEMA_signal_3049), .B0_t (SubCellInst_SboxInst_1_T2), .B0_f (new_AGEMA_signal_2331), .B1_t (new_AGEMA_signal_2332), .B1_f (new_AGEMA_signal_2333), .Z0_t (SubCellInst_SboxInst_1_L0), .Z0_f (new_AGEMA_signal_3278), .Z1_t (new_AGEMA_signal_3279), .Z1_f (new_AGEMA_signal_3280) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_1_XX[2]), .A0_f (new_AGEMA_signal_1375), .A1_t (new_AGEMA_signal_1376), .A1_f (new_AGEMA_signal_1377), .B0_t (Ciphertext_s0_t[6]), .B0_f (Ciphertext_s0_f[6]), .B1_t (Ciphertext_s1_t[6]), .B1_f (Ciphertext_s1_f[6]), .Z0_t (SubCellInst_SboxInst_1_Q6), .Z0_f (new_AGEMA_signal_2334), .Z1_t (new_AGEMA_signal_2335), .Z1_f (new_AGEMA_signal_2336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_1_Q1), .A0_f (new_AGEMA_signal_2328), .A1_t (new_AGEMA_signal_2329), .A1_f (new_AGEMA_signal_2330), .B0_t (SubCellInst_SboxInst_1_Q6), .B0_f (new_AGEMA_signal_2334), .B1_t (new_AGEMA_signal_2335), .B1_f (new_AGEMA_signal_2336), .Z0_t (SubCellInst_SboxInst_1_L1), .Z0_f (new_AGEMA_signal_2713), .Z1_t (new_AGEMA_signal_2714), .Z1_f (new_AGEMA_signal_2715) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_1_L1), .A0_f (new_AGEMA_signal_2713), .A1_t (new_AGEMA_signal_2714), .A1_f (new_AGEMA_signal_2715), .B0_t (SubCellInst_SboxInst_1_T2), .B0_f (new_AGEMA_signal_2331), .B1_t (new_AGEMA_signal_2332), .B1_f (new_AGEMA_signal_2333), .Z0_t (SubCellInst_SboxInst_1_Q7), .Z0_f (new_AGEMA_signal_2861), .Z1_t (new_AGEMA_signal_2862), .Z1_f (new_AGEMA_signal_2863) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_AND4_U1 ( .A0_t (SubCellInst_SboxInst_1_Q6), .A0_f (new_AGEMA_signal_2334), .A1_t (new_AGEMA_signal_2335), .A1_f (new_AGEMA_signal_2336), .B0_t (SubCellInst_SboxInst_1_Q7), .B0_f (new_AGEMA_signal_2861), .B1_t (new_AGEMA_signal_2862), .B1_f (new_AGEMA_signal_2863), .Z0_t (SubCellInst_SboxInst_1_T3), .Z0_f (new_AGEMA_signal_3050), .Z1_t (new_AGEMA_signal_3051), .Z1_f (new_AGEMA_signal_3052) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR8_U1 ( .A0_t (Ciphertext_s0_t[5]), .A0_f (Ciphertext_s0_f[5]), .A1_t (Ciphertext_s1_t[5]), .A1_f (Ciphertext_s1_f[5]), .B0_t (Ciphertext_s0_t[6]), .B0_f (Ciphertext_s0_f[6]), .B1_t (Ciphertext_s1_t[6]), .B1_f (Ciphertext_s1_f[6]), .Z0_t (SubCellInst_SboxInst_1_L2), .Z0_f (new_AGEMA_signal_1384), .Z1_t (new_AGEMA_signal_1385), .Z1_f (new_AGEMA_signal_1386) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_1_L0), .A0_f (new_AGEMA_signal_3278), .A1_t (new_AGEMA_signal_3279), .A1_f (new_AGEMA_signal_3280), .B0_t (SubCellInst_SboxInst_1_L2), .B0_f (new_AGEMA_signal_1384), .B1_t (new_AGEMA_signal_1385), .B1_f (new_AGEMA_signal_1386), .Z0_t (SubCellInst_SboxInst_1_YY_3), .Z0_f (new_AGEMA_signal_3435), .Z1_t (new_AGEMA_signal_3436), .Z1_f (new_AGEMA_signal_3437) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_1_L0), .A0_f (new_AGEMA_signal_3278), .A1_t (new_AGEMA_signal_3279), .A1_f (new_AGEMA_signal_3280), .B0_t (SubCellInst_SboxInst_1_T3), .B0_f (new_AGEMA_signal_3050), .B1_t (new_AGEMA_signal_3051), .B1_f (new_AGEMA_signal_3052), .Z0_t (ShiftRowsOutput[8]), .Z0_f (new_AGEMA_signal_3438), .Z1_t (new_AGEMA_signal_3439), .Z1_f (new_AGEMA_signal_3440) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_1_XX[2]), .A0_f (new_AGEMA_signal_1375), .A1_t (new_AGEMA_signal_1376), .A1_f (new_AGEMA_signal_1377), .B0_t (SubCellInst_SboxInst_1_T0), .B0_f (new_AGEMA_signal_2710), .B1_t (new_AGEMA_signal_2711), .B1_f (new_AGEMA_signal_2712), .Z0_t (SubCellInst_SboxInst_1_L3), .Z0_f (new_AGEMA_signal_2864), .Z1_t (new_AGEMA_signal_2865), .Z1_f (new_AGEMA_signal_2866) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_1_L3), .A0_f (new_AGEMA_signal_2864), .A1_t (new_AGEMA_signal_2865), .A1_f (new_AGEMA_signal_2866), .B0_t (SubCellInst_SboxInst_1_T2), .B0_f (new_AGEMA_signal_2331), .B1_t (new_AGEMA_signal_2332), .B1_f (new_AGEMA_signal_2333), .Z0_t (SubCellInst_SboxInst_1_YY[1]), .Z0_f (new_AGEMA_signal_3053), .Z1_t (new_AGEMA_signal_3054), .Z1_f (new_AGEMA_signal_3055) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_1_XX[1]), .A0_f (new_AGEMA_signal_1369), .A1_t (new_AGEMA_signal_1370), .A1_f (new_AGEMA_signal_1371), .B0_t (SubCellInst_SboxInst_1_T2), .B0_f (new_AGEMA_signal_2331), .B1_t (new_AGEMA_signal_2332), .B1_f (new_AGEMA_signal_2333), .Z0_t (SubCellInst_SboxInst_1_YY[0]), .Z0_f (new_AGEMA_signal_2716), .Z1_t (new_AGEMA_signal_2717), .Z1_f (new_AGEMA_signal_2718) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_1_YY[1]), .A0_f (new_AGEMA_signal_3053), .A1_t (new_AGEMA_signal_3054), .A1_f (new_AGEMA_signal_3055), .B0_t (SubCellInst_SboxInst_1_YY_3), .B0_f (new_AGEMA_signal_3435), .B1_t (new_AGEMA_signal_3436), .B1_f (new_AGEMA_signal_3437), .Z0_t (ShiftRowsOutput[9]), .Z0_f (new_AGEMA_signal_3639), .Z1_t (new_AGEMA_signal_3640), .Z1_f (new_AGEMA_signal_3641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[10]), .A0_f (Ciphertext_s0_f[10]), .A1_t (Ciphertext_s1_t[10]), .A1_f (Ciphertext_s1_f[10]), .B0_t (Ciphertext_s0_t[11]), .B0_f (Ciphertext_s0_f[11]), .B1_t (Ciphertext_s1_t[11]), .B1_f (Ciphertext_s1_f[11]), .Z0_t (SubCellInst_SboxInst_2_XX[1]), .Z0_f (new_AGEMA_signal_1393), .Z1_t (new_AGEMA_signal_1394), .Z1_f (new_AGEMA_signal_1395) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[8]), .A0_f (Ciphertext_s0_f[8]), .A1_t (Ciphertext_s1_t[8]), .A1_f (Ciphertext_s1_f[8]), .B0_t (Ciphertext_s0_t[10]), .B0_f (Ciphertext_s0_f[10]), .B1_t (Ciphertext_s1_t[10]), .B1_f (Ciphertext_s1_f[10]), .Z0_t (SubCellInst_SboxInst_2_XX[2]), .Z0_f (new_AGEMA_signal_1399), .Z1_t (new_AGEMA_signal_1400), .Z1_f (new_AGEMA_signal_1401) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR0_U1 ( .A0_t (Ciphertext_s0_t[9]), .A0_f (Ciphertext_s0_f[9]), .A1_t (Ciphertext_s1_t[9]), .A1_f (Ciphertext_s1_f[9]), .B0_t (SubCellInst_SboxInst_2_XX[2]), .B0_f (new_AGEMA_signal_1399), .B1_t (new_AGEMA_signal_1400), .B1_f (new_AGEMA_signal_1401), .Z0_t (SubCellInst_SboxInst_2_Q0), .Z0_f (new_AGEMA_signal_2337), .Z1_t (new_AGEMA_signal_2338), .Z1_f (new_AGEMA_signal_2339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR1_U1 ( .A0_t (Ciphertext_s0_t[9]), .A0_f (Ciphertext_s0_f[9]), .A1_t (Ciphertext_s1_t[9]), .A1_f (Ciphertext_s1_f[9]), .B0_t (SubCellInst_SboxInst_2_XX[1]), .B0_f (new_AGEMA_signal_1393), .B1_t (new_AGEMA_signal_1394), .B1_f (new_AGEMA_signal_1395), .Z0_t (SubCellInst_SboxInst_2_Q1), .Z0_f (new_AGEMA_signal_2340), .Z1_t (new_AGEMA_signal_2341), .Z1_f (new_AGEMA_signal_2342) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_AND1_U1 ( .A0_t (Ciphertext_s0_t[10]), .A0_f (Ciphertext_s0_f[10]), .A1_t (Ciphertext_s1_t[10]), .A1_f (Ciphertext_s1_f[10]), .B0_t (SubCellInst_SboxInst_2_Q1), .B0_f (new_AGEMA_signal_2340), .B1_t (new_AGEMA_signal_2341), .B1_f (new_AGEMA_signal_2342), .Z0_t (SubCellInst_SboxInst_2_T0), .Z0_f (new_AGEMA_signal_2719), .Z1_t (new_AGEMA_signal_2720), .Z1_f (new_AGEMA_signal_2721) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_2_Q0), .A0_f (new_AGEMA_signal_2337), .A1_t (new_AGEMA_signal_2338), .A1_f (new_AGEMA_signal_2339), .B0_t (SubCellInst_SboxInst_2_T0), .B0_f (new_AGEMA_signal_2719), .B1_t (new_AGEMA_signal_2720), .B1_f (new_AGEMA_signal_2721), .Z0_t (SubCellInst_SboxInst_2_Q2), .Z0_f (new_AGEMA_signal_2867), .Z1_t (new_AGEMA_signal_2868), .Z1_f (new_AGEMA_signal_2869) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_AND2_U1 ( .A0_t (Ciphertext_s0_t[9]), .A0_f (Ciphertext_s0_f[9]), .A1_t (Ciphertext_s1_t[9]), .A1_f (Ciphertext_s1_f[9]), .B0_t (SubCellInst_SboxInst_2_Q2), .B0_f (new_AGEMA_signal_2867), .B1_t (new_AGEMA_signal_2868), .B1_f (new_AGEMA_signal_2869), .Z0_t (SubCellInst_SboxInst_2_T1), .Z0_f (new_AGEMA_signal_3056), .Z1_t (new_AGEMA_signal_3057), .Z1_f (new_AGEMA_signal_3058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_XOR3_U1 ( .A0_t (Ciphertext_s0_t[9]), .A0_f (Ciphertext_s0_f[9]), .A1_t (Ciphertext_s1_t[9]), .A1_f (Ciphertext_s1_f[9]), .B0_t (Ciphertext_s0_t[10]), .B0_f (Ciphertext_s0_f[10]), .B1_t (Ciphertext_s1_t[10]), .B1_f (Ciphertext_s1_f[10]), .Z0_t (SubCellInst_SboxInst_2_Q4), .Z0_f (new_AGEMA_signal_1405), .Z1_t (new_AGEMA_signal_1406), .Z1_f (new_AGEMA_signal_1407) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_AND3_U1 ( .A0_t (Ciphertext_s0_t[10]), .A0_f (Ciphertext_s0_f[10]), .A1_t (Ciphertext_s1_t[10]), .A1_f (Ciphertext_s1_f[10]), .B0_t (SubCellInst_SboxInst_2_Q4), .B0_f (new_AGEMA_signal_1405), .B1_t (new_AGEMA_signal_1406), .B1_f (new_AGEMA_signal_1407), .Z0_t (SubCellInst_SboxInst_2_T2), .Z0_f (new_AGEMA_signal_2343), .Z1_t (new_AGEMA_signal_2344), .Z1_f (new_AGEMA_signal_2345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_2_T1), .A0_f (new_AGEMA_signal_3056), .A1_t (new_AGEMA_signal_3057), .A1_f (new_AGEMA_signal_3058), .B0_t (SubCellInst_SboxInst_2_T2), .B0_f (new_AGEMA_signal_2343), .B1_t (new_AGEMA_signal_2344), .B1_f (new_AGEMA_signal_2345), .Z0_t (SubCellInst_SboxInst_2_L0), .Z0_f (new_AGEMA_signal_3281), .Z1_t (new_AGEMA_signal_3282), .Z1_f (new_AGEMA_signal_3283) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_2_XX[2]), .A0_f (new_AGEMA_signal_1399), .A1_t (new_AGEMA_signal_1400), .A1_f (new_AGEMA_signal_1401), .B0_t (Ciphertext_s0_t[10]), .B0_f (Ciphertext_s0_f[10]), .B1_t (Ciphertext_s1_t[10]), .B1_f (Ciphertext_s1_f[10]), .Z0_t (SubCellInst_SboxInst_2_Q6), .Z0_f (new_AGEMA_signal_2346), .Z1_t (new_AGEMA_signal_2347), .Z1_f (new_AGEMA_signal_2348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_2_Q1), .A0_f (new_AGEMA_signal_2340), .A1_t (new_AGEMA_signal_2341), .A1_f (new_AGEMA_signal_2342), .B0_t (SubCellInst_SboxInst_2_Q6), .B0_f (new_AGEMA_signal_2346), .B1_t (new_AGEMA_signal_2347), .B1_f (new_AGEMA_signal_2348), .Z0_t (SubCellInst_SboxInst_2_L1), .Z0_f (new_AGEMA_signal_2722), .Z1_t (new_AGEMA_signal_2723), .Z1_f (new_AGEMA_signal_2724) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_2_L1), .A0_f (new_AGEMA_signal_2722), .A1_t (new_AGEMA_signal_2723), .A1_f (new_AGEMA_signal_2724), .B0_t (SubCellInst_SboxInst_2_T2), .B0_f (new_AGEMA_signal_2343), .B1_t (new_AGEMA_signal_2344), .B1_f (new_AGEMA_signal_2345), .Z0_t (SubCellInst_SboxInst_2_Q7), .Z0_f (new_AGEMA_signal_2870), .Z1_t (new_AGEMA_signal_2871), .Z1_f (new_AGEMA_signal_2872) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_AND4_U1 ( .A0_t (SubCellInst_SboxInst_2_Q6), .A0_f (new_AGEMA_signal_2346), .A1_t (new_AGEMA_signal_2347), .A1_f (new_AGEMA_signal_2348), .B0_t (SubCellInst_SboxInst_2_Q7), .B0_f (new_AGEMA_signal_2870), .B1_t (new_AGEMA_signal_2871), .B1_f (new_AGEMA_signal_2872), .Z0_t (SubCellInst_SboxInst_2_T3), .Z0_f (new_AGEMA_signal_3059), .Z1_t (new_AGEMA_signal_3060), .Z1_f (new_AGEMA_signal_3061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR8_U1 ( .A0_t (Ciphertext_s0_t[9]), .A0_f (Ciphertext_s0_f[9]), .A1_t (Ciphertext_s1_t[9]), .A1_f (Ciphertext_s1_f[9]), .B0_t (Ciphertext_s0_t[10]), .B0_f (Ciphertext_s0_f[10]), .B1_t (Ciphertext_s1_t[10]), .B1_f (Ciphertext_s1_f[10]), .Z0_t (SubCellInst_SboxInst_2_L2), .Z0_f (new_AGEMA_signal_1408), .Z1_t (new_AGEMA_signal_1409), .Z1_f (new_AGEMA_signal_1410) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_2_L0), .A0_f (new_AGEMA_signal_3281), .A1_t (new_AGEMA_signal_3282), .A1_f (new_AGEMA_signal_3283), .B0_t (SubCellInst_SboxInst_2_L2), .B0_f (new_AGEMA_signal_1408), .B1_t (new_AGEMA_signal_1409), .B1_f (new_AGEMA_signal_1410), .Z0_t (SubCellInst_SboxInst_2_YY_3), .Z0_f (new_AGEMA_signal_3441), .Z1_t (new_AGEMA_signal_3442), .Z1_f (new_AGEMA_signal_3443) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_2_L0), .A0_f (new_AGEMA_signal_3281), .A1_t (new_AGEMA_signal_3282), .A1_f (new_AGEMA_signal_3283), .B0_t (SubCellInst_SboxInst_2_T3), .B0_f (new_AGEMA_signal_3059), .B1_t (new_AGEMA_signal_3060), .B1_f (new_AGEMA_signal_3061), .Z0_t (ShiftRowsOutput[12]), .Z0_f (new_AGEMA_signal_3444), .Z1_t (new_AGEMA_signal_3445), .Z1_f (new_AGEMA_signal_3446) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_2_XX[2]), .A0_f (new_AGEMA_signal_1399), .A1_t (new_AGEMA_signal_1400), .A1_f (new_AGEMA_signal_1401), .B0_t (SubCellInst_SboxInst_2_T0), .B0_f (new_AGEMA_signal_2719), .B1_t (new_AGEMA_signal_2720), .B1_f (new_AGEMA_signal_2721), .Z0_t (SubCellInst_SboxInst_2_L3), .Z0_f (new_AGEMA_signal_2873), .Z1_t (new_AGEMA_signal_2874), .Z1_f (new_AGEMA_signal_2875) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_2_L3), .A0_f (new_AGEMA_signal_2873), .A1_t (new_AGEMA_signal_2874), .A1_f (new_AGEMA_signal_2875), .B0_t (SubCellInst_SboxInst_2_T2), .B0_f (new_AGEMA_signal_2343), .B1_t (new_AGEMA_signal_2344), .B1_f (new_AGEMA_signal_2345), .Z0_t (SubCellInst_SboxInst_2_YY[1]), .Z0_f (new_AGEMA_signal_3062), .Z1_t (new_AGEMA_signal_3063), .Z1_f (new_AGEMA_signal_3064) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_2_XX[1]), .A0_f (new_AGEMA_signal_1393), .A1_t (new_AGEMA_signal_1394), .A1_f (new_AGEMA_signal_1395), .B0_t (SubCellInst_SboxInst_2_T2), .B0_f (new_AGEMA_signal_2343), .B1_t (new_AGEMA_signal_2344), .B1_f (new_AGEMA_signal_2345), .Z0_t (SubCellInst_SboxInst_2_YY[0]), .Z0_f (new_AGEMA_signal_2725), .Z1_t (new_AGEMA_signal_2726), .Z1_f (new_AGEMA_signal_2727) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_2_YY[1]), .A0_f (new_AGEMA_signal_3062), .A1_t (new_AGEMA_signal_3063), .A1_f (new_AGEMA_signal_3064), .B0_t (SubCellInst_SboxInst_2_YY_3), .B0_f (new_AGEMA_signal_3441), .B1_t (new_AGEMA_signal_3442), .B1_f (new_AGEMA_signal_3443), .Z0_t (ShiftRowsOutput[13]), .Z0_f (new_AGEMA_signal_3642), .Z1_t (new_AGEMA_signal_3643), .Z1_f (new_AGEMA_signal_3644) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[14]), .A0_f (Ciphertext_s0_f[14]), .A1_t (Ciphertext_s1_t[14]), .A1_f (Ciphertext_s1_f[14]), .B0_t (Ciphertext_s0_t[15]), .B0_f (Ciphertext_s0_f[15]), .B1_t (Ciphertext_s1_t[15]), .B1_f (Ciphertext_s1_f[15]), .Z0_t (SubCellInst_SboxInst_3_XX[1]), .Z0_f (new_AGEMA_signal_1417), .Z1_t (new_AGEMA_signal_1418), .Z1_f (new_AGEMA_signal_1419) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[12]), .A0_f (Ciphertext_s0_f[12]), .A1_t (Ciphertext_s1_t[12]), .A1_f (Ciphertext_s1_f[12]), .B0_t (Ciphertext_s0_t[14]), .B0_f (Ciphertext_s0_f[14]), .B1_t (Ciphertext_s1_t[14]), .B1_f (Ciphertext_s1_f[14]), .Z0_t (SubCellInst_SboxInst_3_XX[2]), .Z0_f (new_AGEMA_signal_1423), .Z1_t (new_AGEMA_signal_1424), .Z1_f (new_AGEMA_signal_1425) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR0_U1 ( .A0_t (Ciphertext_s0_t[13]), .A0_f (Ciphertext_s0_f[13]), .A1_t (Ciphertext_s1_t[13]), .A1_f (Ciphertext_s1_f[13]), .B0_t (SubCellInst_SboxInst_3_XX[2]), .B0_f (new_AGEMA_signal_1423), .B1_t (new_AGEMA_signal_1424), .B1_f (new_AGEMA_signal_1425), .Z0_t (SubCellInst_SboxInst_3_Q0), .Z0_f (new_AGEMA_signal_2349), .Z1_t (new_AGEMA_signal_2350), .Z1_f (new_AGEMA_signal_2351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR1_U1 ( .A0_t (Ciphertext_s0_t[13]), .A0_f (Ciphertext_s0_f[13]), .A1_t (Ciphertext_s1_t[13]), .A1_f (Ciphertext_s1_f[13]), .B0_t (SubCellInst_SboxInst_3_XX[1]), .B0_f (new_AGEMA_signal_1417), .B1_t (new_AGEMA_signal_1418), .B1_f (new_AGEMA_signal_1419), .Z0_t (SubCellInst_SboxInst_3_Q1), .Z0_f (new_AGEMA_signal_2352), .Z1_t (new_AGEMA_signal_2353), .Z1_f (new_AGEMA_signal_2354) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_AND1_U1 ( .A0_t (Ciphertext_s0_t[14]), .A0_f (Ciphertext_s0_f[14]), .A1_t (Ciphertext_s1_t[14]), .A1_f (Ciphertext_s1_f[14]), .B0_t (SubCellInst_SboxInst_3_Q1), .B0_f (new_AGEMA_signal_2352), .B1_t (new_AGEMA_signal_2353), .B1_f (new_AGEMA_signal_2354), .Z0_t (SubCellInst_SboxInst_3_T0), .Z0_f (new_AGEMA_signal_2728), .Z1_t (new_AGEMA_signal_2729), .Z1_f (new_AGEMA_signal_2730) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_3_Q0), .A0_f (new_AGEMA_signal_2349), .A1_t (new_AGEMA_signal_2350), .A1_f (new_AGEMA_signal_2351), .B0_t (SubCellInst_SboxInst_3_T0), .B0_f (new_AGEMA_signal_2728), .B1_t (new_AGEMA_signal_2729), .B1_f (new_AGEMA_signal_2730), .Z0_t (SubCellInst_SboxInst_3_Q2), .Z0_f (new_AGEMA_signal_2876), .Z1_t (new_AGEMA_signal_2877), .Z1_f (new_AGEMA_signal_2878) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_AND2_U1 ( .A0_t (Ciphertext_s0_t[13]), .A0_f (Ciphertext_s0_f[13]), .A1_t (Ciphertext_s1_t[13]), .A1_f (Ciphertext_s1_f[13]), .B0_t (SubCellInst_SboxInst_3_Q2), .B0_f (new_AGEMA_signal_2876), .B1_t (new_AGEMA_signal_2877), .B1_f (new_AGEMA_signal_2878), .Z0_t (SubCellInst_SboxInst_3_T1), .Z0_f (new_AGEMA_signal_3065), .Z1_t (new_AGEMA_signal_3066), .Z1_f (new_AGEMA_signal_3067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_XOR3_U1 ( .A0_t (Ciphertext_s0_t[13]), .A0_f (Ciphertext_s0_f[13]), .A1_t (Ciphertext_s1_t[13]), .A1_f (Ciphertext_s1_f[13]), .B0_t (Ciphertext_s0_t[14]), .B0_f (Ciphertext_s0_f[14]), .B1_t (Ciphertext_s1_t[14]), .B1_f (Ciphertext_s1_f[14]), .Z0_t (SubCellInst_SboxInst_3_Q4), .Z0_f (new_AGEMA_signal_1429), .Z1_t (new_AGEMA_signal_1430), .Z1_f (new_AGEMA_signal_1431) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_AND3_U1 ( .A0_t (Ciphertext_s0_t[14]), .A0_f (Ciphertext_s0_f[14]), .A1_t (Ciphertext_s1_t[14]), .A1_f (Ciphertext_s1_f[14]), .B0_t (SubCellInst_SboxInst_3_Q4), .B0_f (new_AGEMA_signal_1429), .B1_t (new_AGEMA_signal_1430), .B1_f (new_AGEMA_signal_1431), .Z0_t (SubCellInst_SboxInst_3_T2), .Z0_f (new_AGEMA_signal_2355), .Z1_t (new_AGEMA_signal_2356), .Z1_f (new_AGEMA_signal_2357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_3_T1), .A0_f (new_AGEMA_signal_3065), .A1_t (new_AGEMA_signal_3066), .A1_f (new_AGEMA_signal_3067), .B0_t (SubCellInst_SboxInst_3_T2), .B0_f (new_AGEMA_signal_2355), .B1_t (new_AGEMA_signal_2356), .B1_f (new_AGEMA_signal_2357), .Z0_t (SubCellInst_SboxInst_3_L0), .Z0_f (new_AGEMA_signal_3284), .Z1_t (new_AGEMA_signal_3285), .Z1_f (new_AGEMA_signal_3286) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_3_XX[2]), .A0_f (new_AGEMA_signal_1423), .A1_t (new_AGEMA_signal_1424), .A1_f (new_AGEMA_signal_1425), .B0_t (Ciphertext_s0_t[14]), .B0_f (Ciphertext_s0_f[14]), .B1_t (Ciphertext_s1_t[14]), .B1_f (Ciphertext_s1_f[14]), .Z0_t (SubCellInst_SboxInst_3_Q6), .Z0_f (new_AGEMA_signal_2358), .Z1_t (new_AGEMA_signal_2359), .Z1_f (new_AGEMA_signal_2360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_3_Q1), .A0_f (new_AGEMA_signal_2352), .A1_t (new_AGEMA_signal_2353), .A1_f (new_AGEMA_signal_2354), .B0_t (SubCellInst_SboxInst_3_Q6), .B0_f (new_AGEMA_signal_2358), .B1_t (new_AGEMA_signal_2359), .B1_f (new_AGEMA_signal_2360), .Z0_t (SubCellInst_SboxInst_3_L1), .Z0_f (new_AGEMA_signal_2731), .Z1_t (new_AGEMA_signal_2732), .Z1_f (new_AGEMA_signal_2733) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_3_L1), .A0_f (new_AGEMA_signal_2731), .A1_t (new_AGEMA_signal_2732), .A1_f (new_AGEMA_signal_2733), .B0_t (SubCellInst_SboxInst_3_T2), .B0_f (new_AGEMA_signal_2355), .B1_t (new_AGEMA_signal_2356), .B1_f (new_AGEMA_signal_2357), .Z0_t (SubCellInst_SboxInst_3_Q7), .Z0_f (new_AGEMA_signal_2879), .Z1_t (new_AGEMA_signal_2880), .Z1_f (new_AGEMA_signal_2881) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_AND4_U1 ( .A0_t (SubCellInst_SboxInst_3_Q6), .A0_f (new_AGEMA_signal_2358), .A1_t (new_AGEMA_signal_2359), .A1_f (new_AGEMA_signal_2360), .B0_t (SubCellInst_SboxInst_3_Q7), .B0_f (new_AGEMA_signal_2879), .B1_t (new_AGEMA_signal_2880), .B1_f (new_AGEMA_signal_2881), .Z0_t (SubCellInst_SboxInst_3_T3), .Z0_f (new_AGEMA_signal_3068), .Z1_t (new_AGEMA_signal_3069), .Z1_f (new_AGEMA_signal_3070) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR8_U1 ( .A0_t (Ciphertext_s0_t[13]), .A0_f (Ciphertext_s0_f[13]), .A1_t (Ciphertext_s1_t[13]), .A1_f (Ciphertext_s1_f[13]), .B0_t (Ciphertext_s0_t[14]), .B0_f (Ciphertext_s0_f[14]), .B1_t (Ciphertext_s1_t[14]), .B1_f (Ciphertext_s1_f[14]), .Z0_t (SubCellInst_SboxInst_3_L2), .Z0_f (new_AGEMA_signal_1432), .Z1_t (new_AGEMA_signal_1433), .Z1_f (new_AGEMA_signal_1434) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_3_L0), .A0_f (new_AGEMA_signal_3284), .A1_t (new_AGEMA_signal_3285), .A1_f (new_AGEMA_signal_3286), .B0_t (SubCellInst_SboxInst_3_L2), .B0_f (new_AGEMA_signal_1432), .B1_t (new_AGEMA_signal_1433), .B1_f (new_AGEMA_signal_1434), .Z0_t (SubCellInst_SboxInst_3_YY_3), .Z0_f (new_AGEMA_signal_3447), .Z1_t (new_AGEMA_signal_3448), .Z1_f (new_AGEMA_signal_3449) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_3_L0), .A0_f (new_AGEMA_signal_3284), .A1_t (new_AGEMA_signal_3285), .A1_f (new_AGEMA_signal_3286), .B0_t (SubCellInst_SboxInst_3_T3), .B0_f (new_AGEMA_signal_3068), .B1_t (new_AGEMA_signal_3069), .B1_f (new_AGEMA_signal_3070), .Z0_t (ShiftRowsOutput[0]), .Z0_f (new_AGEMA_signal_3450), .Z1_t (new_AGEMA_signal_3451), .Z1_f (new_AGEMA_signal_3452) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_3_XX[2]), .A0_f (new_AGEMA_signal_1423), .A1_t (new_AGEMA_signal_1424), .A1_f (new_AGEMA_signal_1425), .B0_t (SubCellInst_SboxInst_3_T0), .B0_f (new_AGEMA_signal_2728), .B1_t (new_AGEMA_signal_2729), .B1_f (new_AGEMA_signal_2730), .Z0_t (SubCellInst_SboxInst_3_L3), .Z0_f (new_AGEMA_signal_2882), .Z1_t (new_AGEMA_signal_2883), .Z1_f (new_AGEMA_signal_2884) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_3_L3), .A0_f (new_AGEMA_signal_2882), .A1_t (new_AGEMA_signal_2883), .A1_f (new_AGEMA_signal_2884), .B0_t (SubCellInst_SboxInst_3_T2), .B0_f (new_AGEMA_signal_2355), .B1_t (new_AGEMA_signal_2356), .B1_f (new_AGEMA_signal_2357), .Z0_t (SubCellInst_SboxInst_3_YY[1]), .Z0_f (new_AGEMA_signal_3071), .Z1_t (new_AGEMA_signal_3072), .Z1_f (new_AGEMA_signal_3073) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_3_XX[1]), .A0_f (new_AGEMA_signal_1417), .A1_t (new_AGEMA_signal_1418), .A1_f (new_AGEMA_signal_1419), .B0_t (SubCellInst_SboxInst_3_T2), .B0_f (new_AGEMA_signal_2355), .B1_t (new_AGEMA_signal_2356), .B1_f (new_AGEMA_signal_2357), .Z0_t (SubCellInst_SboxInst_3_YY[0]), .Z0_f (new_AGEMA_signal_2734), .Z1_t (new_AGEMA_signal_2735), .Z1_f (new_AGEMA_signal_2736) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_3_YY[1]), .A0_f (new_AGEMA_signal_3071), .A1_t (new_AGEMA_signal_3072), .A1_f (new_AGEMA_signal_3073), .B0_t (SubCellInst_SboxInst_3_YY_3), .B0_f (new_AGEMA_signal_3447), .B1_t (new_AGEMA_signal_3448), .B1_f (new_AGEMA_signal_3449), .Z0_t (ShiftRowsOutput[1]), .Z0_f (new_AGEMA_signal_3645), .Z1_t (new_AGEMA_signal_3646), .Z1_f (new_AGEMA_signal_3647) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[18]), .A0_f (Ciphertext_s0_f[18]), .A1_t (Ciphertext_s1_t[18]), .A1_f (Ciphertext_s1_f[18]), .B0_t (Ciphertext_s0_t[19]), .B0_f (Ciphertext_s0_f[19]), .B1_t (Ciphertext_s1_t[19]), .B1_f (Ciphertext_s1_f[19]), .Z0_t (SubCellInst_SboxInst_4_XX[1]), .Z0_f (new_AGEMA_signal_1441), .Z1_t (new_AGEMA_signal_1442), .Z1_f (new_AGEMA_signal_1443) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[16]), .A0_f (Ciphertext_s0_f[16]), .A1_t (Ciphertext_s1_t[16]), .A1_f (Ciphertext_s1_f[16]), .B0_t (Ciphertext_s0_t[18]), .B0_f (Ciphertext_s0_f[18]), .B1_t (Ciphertext_s1_t[18]), .B1_f (Ciphertext_s1_f[18]), .Z0_t (SubCellInst_SboxInst_4_XX[2]), .Z0_f (new_AGEMA_signal_1447), .Z1_t (new_AGEMA_signal_1448), .Z1_f (new_AGEMA_signal_1449) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR0_U1 ( .A0_t (Ciphertext_s0_t[17]), .A0_f (Ciphertext_s0_f[17]), .A1_t (Ciphertext_s1_t[17]), .A1_f (Ciphertext_s1_f[17]), .B0_t (SubCellInst_SboxInst_4_XX[2]), .B0_f (new_AGEMA_signal_1447), .B1_t (new_AGEMA_signal_1448), .B1_f (new_AGEMA_signal_1449), .Z0_t (SubCellInst_SboxInst_4_Q0), .Z0_f (new_AGEMA_signal_2361), .Z1_t (new_AGEMA_signal_2362), .Z1_f (new_AGEMA_signal_2363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR1_U1 ( .A0_t (Ciphertext_s0_t[17]), .A0_f (Ciphertext_s0_f[17]), .A1_t (Ciphertext_s1_t[17]), .A1_f (Ciphertext_s1_f[17]), .B0_t (SubCellInst_SboxInst_4_XX[1]), .B0_f (new_AGEMA_signal_1441), .B1_t (new_AGEMA_signal_1442), .B1_f (new_AGEMA_signal_1443), .Z0_t (SubCellInst_SboxInst_4_Q1), .Z0_f (new_AGEMA_signal_2364), .Z1_t (new_AGEMA_signal_2365), .Z1_f (new_AGEMA_signal_2366) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_AND1_U1 ( .A0_t (Ciphertext_s0_t[18]), .A0_f (Ciphertext_s0_f[18]), .A1_t (Ciphertext_s1_t[18]), .A1_f (Ciphertext_s1_f[18]), .B0_t (SubCellInst_SboxInst_4_Q1), .B0_f (new_AGEMA_signal_2364), .B1_t (new_AGEMA_signal_2365), .B1_f (new_AGEMA_signal_2366), .Z0_t (SubCellInst_SboxInst_4_T0), .Z0_f (new_AGEMA_signal_2737), .Z1_t (new_AGEMA_signal_2738), .Z1_f (new_AGEMA_signal_2739) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_4_Q0), .A0_f (new_AGEMA_signal_2361), .A1_t (new_AGEMA_signal_2362), .A1_f (new_AGEMA_signal_2363), .B0_t (SubCellInst_SboxInst_4_T0), .B0_f (new_AGEMA_signal_2737), .B1_t (new_AGEMA_signal_2738), .B1_f (new_AGEMA_signal_2739), .Z0_t (SubCellInst_SboxInst_4_Q2), .Z0_f (new_AGEMA_signal_2885), .Z1_t (new_AGEMA_signal_2886), .Z1_f (new_AGEMA_signal_2887) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_AND2_U1 ( .A0_t (Ciphertext_s0_t[17]), .A0_f (Ciphertext_s0_f[17]), .A1_t (Ciphertext_s1_t[17]), .A1_f (Ciphertext_s1_f[17]), .B0_t (SubCellInst_SboxInst_4_Q2), .B0_f (new_AGEMA_signal_2885), .B1_t (new_AGEMA_signal_2886), .B1_f (new_AGEMA_signal_2887), .Z0_t (SubCellInst_SboxInst_4_T1), .Z0_f (new_AGEMA_signal_3074), .Z1_t (new_AGEMA_signal_3075), .Z1_f (new_AGEMA_signal_3076) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_XOR3_U1 ( .A0_t (Ciphertext_s0_t[17]), .A0_f (Ciphertext_s0_f[17]), .A1_t (Ciphertext_s1_t[17]), .A1_f (Ciphertext_s1_f[17]), .B0_t (Ciphertext_s0_t[18]), .B0_f (Ciphertext_s0_f[18]), .B1_t (Ciphertext_s1_t[18]), .B1_f (Ciphertext_s1_f[18]), .Z0_t (SubCellInst_SboxInst_4_Q4), .Z0_f (new_AGEMA_signal_1453), .Z1_t (new_AGEMA_signal_1454), .Z1_f (new_AGEMA_signal_1455) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_AND3_U1 ( .A0_t (Ciphertext_s0_t[18]), .A0_f (Ciphertext_s0_f[18]), .A1_t (Ciphertext_s1_t[18]), .A1_f (Ciphertext_s1_f[18]), .B0_t (SubCellInst_SboxInst_4_Q4), .B0_f (new_AGEMA_signal_1453), .B1_t (new_AGEMA_signal_1454), .B1_f (new_AGEMA_signal_1455), .Z0_t (SubCellInst_SboxInst_4_T2), .Z0_f (new_AGEMA_signal_2367), .Z1_t (new_AGEMA_signal_2368), .Z1_f (new_AGEMA_signal_2369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_4_T1), .A0_f (new_AGEMA_signal_3074), .A1_t (new_AGEMA_signal_3075), .A1_f (new_AGEMA_signal_3076), .B0_t (SubCellInst_SboxInst_4_T2), .B0_f (new_AGEMA_signal_2367), .B1_t (new_AGEMA_signal_2368), .B1_f (new_AGEMA_signal_2369), .Z0_t (SubCellInst_SboxInst_4_L0), .Z0_f (new_AGEMA_signal_3287), .Z1_t (new_AGEMA_signal_3288), .Z1_f (new_AGEMA_signal_3289) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_4_XX[2]), .A0_f (new_AGEMA_signal_1447), .A1_t (new_AGEMA_signal_1448), .A1_f (new_AGEMA_signal_1449), .B0_t (Ciphertext_s0_t[18]), .B0_f (Ciphertext_s0_f[18]), .B1_t (Ciphertext_s1_t[18]), .B1_f (Ciphertext_s1_f[18]), .Z0_t (SubCellInst_SboxInst_4_Q6), .Z0_f (new_AGEMA_signal_2370), .Z1_t (new_AGEMA_signal_2371), .Z1_f (new_AGEMA_signal_2372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_4_Q1), .A0_f (new_AGEMA_signal_2364), .A1_t (new_AGEMA_signal_2365), .A1_f (new_AGEMA_signal_2366), .B0_t (SubCellInst_SboxInst_4_Q6), .B0_f (new_AGEMA_signal_2370), .B1_t (new_AGEMA_signal_2371), .B1_f (new_AGEMA_signal_2372), .Z0_t (SubCellInst_SboxInst_4_L1), .Z0_f (new_AGEMA_signal_2740), .Z1_t (new_AGEMA_signal_2741), .Z1_f (new_AGEMA_signal_2742) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_4_L1), .A0_f (new_AGEMA_signal_2740), .A1_t (new_AGEMA_signal_2741), .A1_f (new_AGEMA_signal_2742), .B0_t (SubCellInst_SboxInst_4_T2), .B0_f (new_AGEMA_signal_2367), .B1_t (new_AGEMA_signal_2368), .B1_f (new_AGEMA_signal_2369), .Z0_t (SubCellInst_SboxInst_4_Q7), .Z0_f (new_AGEMA_signal_2888), .Z1_t (new_AGEMA_signal_2889), .Z1_f (new_AGEMA_signal_2890) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_AND4_U1 ( .A0_t (SubCellInst_SboxInst_4_Q6), .A0_f (new_AGEMA_signal_2370), .A1_t (new_AGEMA_signal_2371), .A1_f (new_AGEMA_signal_2372), .B0_t (SubCellInst_SboxInst_4_Q7), .B0_f (new_AGEMA_signal_2888), .B1_t (new_AGEMA_signal_2889), .B1_f (new_AGEMA_signal_2890), .Z0_t (SubCellInst_SboxInst_4_T3), .Z0_f (new_AGEMA_signal_3077), .Z1_t (new_AGEMA_signal_3078), .Z1_f (new_AGEMA_signal_3079) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR8_U1 ( .A0_t (Ciphertext_s0_t[17]), .A0_f (Ciphertext_s0_f[17]), .A1_t (Ciphertext_s1_t[17]), .A1_f (Ciphertext_s1_f[17]), .B0_t (Ciphertext_s0_t[18]), .B0_f (Ciphertext_s0_f[18]), .B1_t (Ciphertext_s1_t[18]), .B1_f (Ciphertext_s1_f[18]), .Z0_t (SubCellInst_SboxInst_4_L2), .Z0_f (new_AGEMA_signal_1456), .Z1_t (new_AGEMA_signal_1457), .Z1_f (new_AGEMA_signal_1458) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_4_L0), .A0_f (new_AGEMA_signal_3287), .A1_t (new_AGEMA_signal_3288), .A1_f (new_AGEMA_signal_3289), .B0_t (SubCellInst_SboxInst_4_L2), .B0_f (new_AGEMA_signal_1456), .B1_t (new_AGEMA_signal_1457), .B1_f (new_AGEMA_signal_1458), .Z0_t (SubCellInst_SboxInst_4_YY_3), .Z0_f (new_AGEMA_signal_3453), .Z1_t (new_AGEMA_signal_3454), .Z1_f (new_AGEMA_signal_3455) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_4_L0), .A0_f (new_AGEMA_signal_3287), .A1_t (new_AGEMA_signal_3288), .A1_f (new_AGEMA_signal_3289), .B0_t (SubCellInst_SboxInst_4_T3), .B0_f (new_AGEMA_signal_3077), .B1_t (new_AGEMA_signal_3078), .B1_f (new_AGEMA_signal_3079), .Z0_t (ShiftRowsOutput[24]), .Z0_f (new_AGEMA_signal_3456), .Z1_t (new_AGEMA_signal_3457), .Z1_f (new_AGEMA_signal_3458) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_4_XX[2]), .A0_f (new_AGEMA_signal_1447), .A1_t (new_AGEMA_signal_1448), .A1_f (new_AGEMA_signal_1449), .B0_t (SubCellInst_SboxInst_4_T0), .B0_f (new_AGEMA_signal_2737), .B1_t (new_AGEMA_signal_2738), .B1_f (new_AGEMA_signal_2739), .Z0_t (SubCellInst_SboxInst_4_L3), .Z0_f (new_AGEMA_signal_2891), .Z1_t (new_AGEMA_signal_2892), .Z1_f (new_AGEMA_signal_2893) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_4_L3), .A0_f (new_AGEMA_signal_2891), .A1_t (new_AGEMA_signal_2892), .A1_f (new_AGEMA_signal_2893), .B0_t (SubCellInst_SboxInst_4_T2), .B0_f (new_AGEMA_signal_2367), .B1_t (new_AGEMA_signal_2368), .B1_f (new_AGEMA_signal_2369), .Z0_t (SubCellInst_SboxInst_4_YY[1]), .Z0_f (new_AGEMA_signal_3080), .Z1_t (new_AGEMA_signal_3081), .Z1_f (new_AGEMA_signal_3082) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_4_XX[1]), .A0_f (new_AGEMA_signal_1441), .A1_t (new_AGEMA_signal_1442), .A1_f (new_AGEMA_signal_1443), .B0_t (SubCellInst_SboxInst_4_T2), .B0_f (new_AGEMA_signal_2367), .B1_t (new_AGEMA_signal_2368), .B1_f (new_AGEMA_signal_2369), .Z0_t (SubCellInst_SboxInst_4_YY[0]), .Z0_f (new_AGEMA_signal_2743), .Z1_t (new_AGEMA_signal_2744), .Z1_f (new_AGEMA_signal_2745) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_4_YY[1]), .A0_f (new_AGEMA_signal_3080), .A1_t (new_AGEMA_signal_3081), .A1_f (new_AGEMA_signal_3082), .B0_t (SubCellInst_SboxInst_4_YY_3), .B0_f (new_AGEMA_signal_3453), .B1_t (new_AGEMA_signal_3454), .B1_f (new_AGEMA_signal_3455), .Z0_t (ShiftRowsOutput[25]), .Z0_f (new_AGEMA_signal_3648), .Z1_t (new_AGEMA_signal_3649), .Z1_f (new_AGEMA_signal_3650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[22]), .A0_f (Ciphertext_s0_f[22]), .A1_t (Ciphertext_s1_t[22]), .A1_f (Ciphertext_s1_f[22]), .B0_t (Ciphertext_s0_t[23]), .B0_f (Ciphertext_s0_f[23]), .B1_t (Ciphertext_s1_t[23]), .B1_f (Ciphertext_s1_f[23]), .Z0_t (SubCellInst_SboxInst_5_XX[1]), .Z0_f (new_AGEMA_signal_1465), .Z1_t (new_AGEMA_signal_1466), .Z1_f (new_AGEMA_signal_1467) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[20]), .A0_f (Ciphertext_s0_f[20]), .A1_t (Ciphertext_s1_t[20]), .A1_f (Ciphertext_s1_f[20]), .B0_t (Ciphertext_s0_t[22]), .B0_f (Ciphertext_s0_f[22]), .B1_t (Ciphertext_s1_t[22]), .B1_f (Ciphertext_s1_f[22]), .Z0_t (SubCellInst_SboxInst_5_XX[2]), .Z0_f (new_AGEMA_signal_1471), .Z1_t (new_AGEMA_signal_1472), .Z1_f (new_AGEMA_signal_1473) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR0_U1 ( .A0_t (Ciphertext_s0_t[21]), .A0_f (Ciphertext_s0_f[21]), .A1_t (Ciphertext_s1_t[21]), .A1_f (Ciphertext_s1_f[21]), .B0_t (SubCellInst_SboxInst_5_XX[2]), .B0_f (new_AGEMA_signal_1471), .B1_t (new_AGEMA_signal_1472), .B1_f (new_AGEMA_signal_1473), .Z0_t (SubCellInst_SboxInst_5_Q0), .Z0_f (new_AGEMA_signal_2373), .Z1_t (new_AGEMA_signal_2374), .Z1_f (new_AGEMA_signal_2375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR1_U1 ( .A0_t (Ciphertext_s0_t[21]), .A0_f (Ciphertext_s0_f[21]), .A1_t (Ciphertext_s1_t[21]), .A1_f (Ciphertext_s1_f[21]), .B0_t (SubCellInst_SboxInst_5_XX[1]), .B0_f (new_AGEMA_signal_1465), .B1_t (new_AGEMA_signal_1466), .B1_f (new_AGEMA_signal_1467), .Z0_t (SubCellInst_SboxInst_5_Q1), .Z0_f (new_AGEMA_signal_2376), .Z1_t (new_AGEMA_signal_2377), .Z1_f (new_AGEMA_signal_2378) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_AND1_U1 ( .A0_t (Ciphertext_s0_t[22]), .A0_f (Ciphertext_s0_f[22]), .A1_t (Ciphertext_s1_t[22]), .A1_f (Ciphertext_s1_f[22]), .B0_t (SubCellInst_SboxInst_5_Q1), .B0_f (new_AGEMA_signal_2376), .B1_t (new_AGEMA_signal_2377), .B1_f (new_AGEMA_signal_2378), .Z0_t (SubCellInst_SboxInst_5_T0), .Z0_f (new_AGEMA_signal_2746), .Z1_t (new_AGEMA_signal_2747), .Z1_f (new_AGEMA_signal_2748) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_5_Q0), .A0_f (new_AGEMA_signal_2373), .A1_t (new_AGEMA_signal_2374), .A1_f (new_AGEMA_signal_2375), .B0_t (SubCellInst_SboxInst_5_T0), .B0_f (new_AGEMA_signal_2746), .B1_t (new_AGEMA_signal_2747), .B1_f (new_AGEMA_signal_2748), .Z0_t (SubCellInst_SboxInst_5_Q2), .Z0_f (new_AGEMA_signal_2894), .Z1_t (new_AGEMA_signal_2895), .Z1_f (new_AGEMA_signal_2896) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_AND2_U1 ( .A0_t (Ciphertext_s0_t[21]), .A0_f (Ciphertext_s0_f[21]), .A1_t (Ciphertext_s1_t[21]), .A1_f (Ciphertext_s1_f[21]), .B0_t (SubCellInst_SboxInst_5_Q2), .B0_f (new_AGEMA_signal_2894), .B1_t (new_AGEMA_signal_2895), .B1_f (new_AGEMA_signal_2896), .Z0_t (SubCellInst_SboxInst_5_T1), .Z0_f (new_AGEMA_signal_3083), .Z1_t (new_AGEMA_signal_3084), .Z1_f (new_AGEMA_signal_3085) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_XOR3_U1 ( .A0_t (Ciphertext_s0_t[21]), .A0_f (Ciphertext_s0_f[21]), .A1_t (Ciphertext_s1_t[21]), .A1_f (Ciphertext_s1_f[21]), .B0_t (Ciphertext_s0_t[22]), .B0_f (Ciphertext_s0_f[22]), .B1_t (Ciphertext_s1_t[22]), .B1_f (Ciphertext_s1_f[22]), .Z0_t (SubCellInst_SboxInst_5_Q4), .Z0_f (new_AGEMA_signal_1477), .Z1_t (new_AGEMA_signal_1478), .Z1_f (new_AGEMA_signal_1479) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_AND3_U1 ( .A0_t (Ciphertext_s0_t[22]), .A0_f (Ciphertext_s0_f[22]), .A1_t (Ciphertext_s1_t[22]), .A1_f (Ciphertext_s1_f[22]), .B0_t (SubCellInst_SboxInst_5_Q4), .B0_f (new_AGEMA_signal_1477), .B1_t (new_AGEMA_signal_1478), .B1_f (new_AGEMA_signal_1479), .Z0_t (SubCellInst_SboxInst_5_T2), .Z0_f (new_AGEMA_signal_2379), .Z1_t (new_AGEMA_signal_2380), .Z1_f (new_AGEMA_signal_2381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_5_T1), .A0_f (new_AGEMA_signal_3083), .A1_t (new_AGEMA_signal_3084), .A1_f (new_AGEMA_signal_3085), .B0_t (SubCellInst_SboxInst_5_T2), .B0_f (new_AGEMA_signal_2379), .B1_t (new_AGEMA_signal_2380), .B1_f (new_AGEMA_signal_2381), .Z0_t (SubCellInst_SboxInst_5_L0), .Z0_f (new_AGEMA_signal_3290), .Z1_t (new_AGEMA_signal_3291), .Z1_f (new_AGEMA_signal_3292) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_5_XX[2]), .A0_f (new_AGEMA_signal_1471), .A1_t (new_AGEMA_signal_1472), .A1_f (new_AGEMA_signal_1473), .B0_t (Ciphertext_s0_t[22]), .B0_f (Ciphertext_s0_f[22]), .B1_t (Ciphertext_s1_t[22]), .B1_f (Ciphertext_s1_f[22]), .Z0_t (SubCellInst_SboxInst_5_Q6), .Z0_f (new_AGEMA_signal_2382), .Z1_t (new_AGEMA_signal_2383), .Z1_f (new_AGEMA_signal_2384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_5_Q1), .A0_f (new_AGEMA_signal_2376), .A1_t (new_AGEMA_signal_2377), .A1_f (new_AGEMA_signal_2378), .B0_t (SubCellInst_SboxInst_5_Q6), .B0_f (new_AGEMA_signal_2382), .B1_t (new_AGEMA_signal_2383), .B1_f (new_AGEMA_signal_2384), .Z0_t (SubCellInst_SboxInst_5_L1), .Z0_f (new_AGEMA_signal_2749), .Z1_t (new_AGEMA_signal_2750), .Z1_f (new_AGEMA_signal_2751) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_5_L1), .A0_f (new_AGEMA_signal_2749), .A1_t (new_AGEMA_signal_2750), .A1_f (new_AGEMA_signal_2751), .B0_t (SubCellInst_SboxInst_5_T2), .B0_f (new_AGEMA_signal_2379), .B1_t (new_AGEMA_signal_2380), .B1_f (new_AGEMA_signal_2381), .Z0_t (SubCellInst_SboxInst_5_Q7), .Z0_f (new_AGEMA_signal_2897), .Z1_t (new_AGEMA_signal_2898), .Z1_f (new_AGEMA_signal_2899) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_AND4_U1 ( .A0_t (SubCellInst_SboxInst_5_Q6), .A0_f (new_AGEMA_signal_2382), .A1_t (new_AGEMA_signal_2383), .A1_f (new_AGEMA_signal_2384), .B0_t (SubCellInst_SboxInst_5_Q7), .B0_f (new_AGEMA_signal_2897), .B1_t (new_AGEMA_signal_2898), .B1_f (new_AGEMA_signal_2899), .Z0_t (SubCellInst_SboxInst_5_T3), .Z0_f (new_AGEMA_signal_3086), .Z1_t (new_AGEMA_signal_3087), .Z1_f (new_AGEMA_signal_3088) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR8_U1 ( .A0_t (Ciphertext_s0_t[21]), .A0_f (Ciphertext_s0_f[21]), .A1_t (Ciphertext_s1_t[21]), .A1_f (Ciphertext_s1_f[21]), .B0_t (Ciphertext_s0_t[22]), .B0_f (Ciphertext_s0_f[22]), .B1_t (Ciphertext_s1_t[22]), .B1_f (Ciphertext_s1_f[22]), .Z0_t (SubCellInst_SboxInst_5_L2), .Z0_f (new_AGEMA_signal_1480), .Z1_t (new_AGEMA_signal_1481), .Z1_f (new_AGEMA_signal_1482) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_5_L0), .A0_f (new_AGEMA_signal_3290), .A1_t (new_AGEMA_signal_3291), .A1_f (new_AGEMA_signal_3292), .B0_t (SubCellInst_SboxInst_5_L2), .B0_f (new_AGEMA_signal_1480), .B1_t (new_AGEMA_signal_1481), .B1_f (new_AGEMA_signal_1482), .Z0_t (SubCellInst_SboxInst_5_YY_3), .Z0_f (new_AGEMA_signal_3459), .Z1_t (new_AGEMA_signal_3460), .Z1_f (new_AGEMA_signal_3461) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_5_L0), .A0_f (new_AGEMA_signal_3290), .A1_t (new_AGEMA_signal_3291), .A1_f (new_AGEMA_signal_3292), .B0_t (SubCellInst_SboxInst_5_T3), .B0_f (new_AGEMA_signal_3086), .B1_t (new_AGEMA_signal_3087), .B1_f (new_AGEMA_signal_3088), .Z0_t (ShiftRowsOutput[28]), .Z0_f (new_AGEMA_signal_3462), .Z1_t (new_AGEMA_signal_3463), .Z1_f (new_AGEMA_signal_3464) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_5_XX[2]), .A0_f (new_AGEMA_signal_1471), .A1_t (new_AGEMA_signal_1472), .A1_f (new_AGEMA_signal_1473), .B0_t (SubCellInst_SboxInst_5_T0), .B0_f (new_AGEMA_signal_2746), .B1_t (new_AGEMA_signal_2747), .B1_f (new_AGEMA_signal_2748), .Z0_t (SubCellInst_SboxInst_5_L3), .Z0_f (new_AGEMA_signal_2900), .Z1_t (new_AGEMA_signal_2901), .Z1_f (new_AGEMA_signal_2902) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_5_L3), .A0_f (new_AGEMA_signal_2900), .A1_t (new_AGEMA_signal_2901), .A1_f (new_AGEMA_signal_2902), .B0_t (SubCellInst_SboxInst_5_T2), .B0_f (new_AGEMA_signal_2379), .B1_t (new_AGEMA_signal_2380), .B1_f (new_AGEMA_signal_2381), .Z0_t (SubCellInst_SboxInst_5_YY[1]), .Z0_f (new_AGEMA_signal_3089), .Z1_t (new_AGEMA_signal_3090), .Z1_f (new_AGEMA_signal_3091) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_5_XX[1]), .A0_f (new_AGEMA_signal_1465), .A1_t (new_AGEMA_signal_1466), .A1_f (new_AGEMA_signal_1467), .B0_t (SubCellInst_SboxInst_5_T2), .B0_f (new_AGEMA_signal_2379), .B1_t (new_AGEMA_signal_2380), .B1_f (new_AGEMA_signal_2381), .Z0_t (SubCellInst_SboxInst_5_YY[0]), .Z0_f (new_AGEMA_signal_2752), .Z1_t (new_AGEMA_signal_2753), .Z1_f (new_AGEMA_signal_2754) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_5_YY[1]), .A0_f (new_AGEMA_signal_3089), .A1_t (new_AGEMA_signal_3090), .A1_f (new_AGEMA_signal_3091), .B0_t (SubCellInst_SboxInst_5_YY_3), .B0_f (new_AGEMA_signal_3459), .B1_t (new_AGEMA_signal_3460), .B1_f (new_AGEMA_signal_3461), .Z0_t (ShiftRowsOutput[29]), .Z0_f (new_AGEMA_signal_3651), .Z1_t (new_AGEMA_signal_3652), .Z1_f (new_AGEMA_signal_3653) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[26]), .A0_f (Ciphertext_s0_f[26]), .A1_t (Ciphertext_s1_t[26]), .A1_f (Ciphertext_s1_f[26]), .B0_t (Ciphertext_s0_t[27]), .B0_f (Ciphertext_s0_f[27]), .B1_t (Ciphertext_s1_t[27]), .B1_f (Ciphertext_s1_f[27]), .Z0_t (SubCellInst_SboxInst_6_XX[1]), .Z0_f (new_AGEMA_signal_1489), .Z1_t (new_AGEMA_signal_1490), .Z1_f (new_AGEMA_signal_1491) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[24]), .A0_f (Ciphertext_s0_f[24]), .A1_t (Ciphertext_s1_t[24]), .A1_f (Ciphertext_s1_f[24]), .B0_t (Ciphertext_s0_t[26]), .B0_f (Ciphertext_s0_f[26]), .B1_t (Ciphertext_s1_t[26]), .B1_f (Ciphertext_s1_f[26]), .Z0_t (SubCellInst_SboxInst_6_XX[2]), .Z0_f (new_AGEMA_signal_1495), .Z1_t (new_AGEMA_signal_1496), .Z1_f (new_AGEMA_signal_1497) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR0_U1 ( .A0_t (Ciphertext_s0_t[25]), .A0_f (Ciphertext_s0_f[25]), .A1_t (Ciphertext_s1_t[25]), .A1_f (Ciphertext_s1_f[25]), .B0_t (SubCellInst_SboxInst_6_XX[2]), .B0_f (new_AGEMA_signal_1495), .B1_t (new_AGEMA_signal_1496), .B1_f (new_AGEMA_signal_1497), .Z0_t (SubCellInst_SboxInst_6_Q0), .Z0_f (new_AGEMA_signal_2385), .Z1_t (new_AGEMA_signal_2386), .Z1_f (new_AGEMA_signal_2387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR1_U1 ( .A0_t (Ciphertext_s0_t[25]), .A0_f (Ciphertext_s0_f[25]), .A1_t (Ciphertext_s1_t[25]), .A1_f (Ciphertext_s1_f[25]), .B0_t (SubCellInst_SboxInst_6_XX[1]), .B0_f (new_AGEMA_signal_1489), .B1_t (new_AGEMA_signal_1490), .B1_f (new_AGEMA_signal_1491), .Z0_t (SubCellInst_SboxInst_6_Q1), .Z0_f (new_AGEMA_signal_2388), .Z1_t (new_AGEMA_signal_2389), .Z1_f (new_AGEMA_signal_2390) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_AND1_U1 ( .A0_t (Ciphertext_s0_t[26]), .A0_f (Ciphertext_s0_f[26]), .A1_t (Ciphertext_s1_t[26]), .A1_f (Ciphertext_s1_f[26]), .B0_t (SubCellInst_SboxInst_6_Q1), .B0_f (new_AGEMA_signal_2388), .B1_t (new_AGEMA_signal_2389), .B1_f (new_AGEMA_signal_2390), .Z0_t (SubCellInst_SboxInst_6_T0), .Z0_f (new_AGEMA_signal_2755), .Z1_t (new_AGEMA_signal_2756), .Z1_f (new_AGEMA_signal_2757) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_6_Q0), .A0_f (new_AGEMA_signal_2385), .A1_t (new_AGEMA_signal_2386), .A1_f (new_AGEMA_signal_2387), .B0_t (SubCellInst_SboxInst_6_T0), .B0_f (new_AGEMA_signal_2755), .B1_t (new_AGEMA_signal_2756), .B1_f (new_AGEMA_signal_2757), .Z0_t (SubCellInst_SboxInst_6_Q2), .Z0_f (new_AGEMA_signal_2903), .Z1_t (new_AGEMA_signal_2904), .Z1_f (new_AGEMA_signal_2905) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_AND2_U1 ( .A0_t (Ciphertext_s0_t[25]), .A0_f (Ciphertext_s0_f[25]), .A1_t (Ciphertext_s1_t[25]), .A1_f (Ciphertext_s1_f[25]), .B0_t (SubCellInst_SboxInst_6_Q2), .B0_f (new_AGEMA_signal_2903), .B1_t (new_AGEMA_signal_2904), .B1_f (new_AGEMA_signal_2905), .Z0_t (SubCellInst_SboxInst_6_T1), .Z0_f (new_AGEMA_signal_3092), .Z1_t (new_AGEMA_signal_3093), .Z1_f (new_AGEMA_signal_3094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_XOR3_U1 ( .A0_t (Ciphertext_s0_t[25]), .A0_f (Ciphertext_s0_f[25]), .A1_t (Ciphertext_s1_t[25]), .A1_f (Ciphertext_s1_f[25]), .B0_t (Ciphertext_s0_t[26]), .B0_f (Ciphertext_s0_f[26]), .B1_t (Ciphertext_s1_t[26]), .B1_f (Ciphertext_s1_f[26]), .Z0_t (SubCellInst_SboxInst_6_Q4), .Z0_f (new_AGEMA_signal_1501), .Z1_t (new_AGEMA_signal_1502), .Z1_f (new_AGEMA_signal_1503) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_AND3_U1 ( .A0_t (Ciphertext_s0_t[26]), .A0_f (Ciphertext_s0_f[26]), .A1_t (Ciphertext_s1_t[26]), .A1_f (Ciphertext_s1_f[26]), .B0_t (SubCellInst_SboxInst_6_Q4), .B0_f (new_AGEMA_signal_1501), .B1_t (new_AGEMA_signal_1502), .B1_f (new_AGEMA_signal_1503), .Z0_t (SubCellInst_SboxInst_6_T2), .Z0_f (new_AGEMA_signal_2391), .Z1_t (new_AGEMA_signal_2392), .Z1_f (new_AGEMA_signal_2393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_6_T1), .A0_f (new_AGEMA_signal_3092), .A1_t (new_AGEMA_signal_3093), .A1_f (new_AGEMA_signal_3094), .B0_t (SubCellInst_SboxInst_6_T2), .B0_f (new_AGEMA_signal_2391), .B1_t (new_AGEMA_signal_2392), .B1_f (new_AGEMA_signal_2393), .Z0_t (SubCellInst_SboxInst_6_L0), .Z0_f (new_AGEMA_signal_3293), .Z1_t (new_AGEMA_signal_3294), .Z1_f (new_AGEMA_signal_3295) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_6_XX[2]), .A0_f (new_AGEMA_signal_1495), .A1_t (new_AGEMA_signal_1496), .A1_f (new_AGEMA_signal_1497), .B0_t (Ciphertext_s0_t[26]), .B0_f (Ciphertext_s0_f[26]), .B1_t (Ciphertext_s1_t[26]), .B1_f (Ciphertext_s1_f[26]), .Z0_t (SubCellInst_SboxInst_6_Q6), .Z0_f (new_AGEMA_signal_2394), .Z1_t (new_AGEMA_signal_2395), .Z1_f (new_AGEMA_signal_2396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_6_Q1), .A0_f (new_AGEMA_signal_2388), .A1_t (new_AGEMA_signal_2389), .A1_f (new_AGEMA_signal_2390), .B0_t (SubCellInst_SboxInst_6_Q6), .B0_f (new_AGEMA_signal_2394), .B1_t (new_AGEMA_signal_2395), .B1_f (new_AGEMA_signal_2396), .Z0_t (SubCellInst_SboxInst_6_L1), .Z0_f (new_AGEMA_signal_2758), .Z1_t (new_AGEMA_signal_2759), .Z1_f (new_AGEMA_signal_2760) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_6_L1), .A0_f (new_AGEMA_signal_2758), .A1_t (new_AGEMA_signal_2759), .A1_f (new_AGEMA_signal_2760), .B0_t (SubCellInst_SboxInst_6_T2), .B0_f (new_AGEMA_signal_2391), .B1_t (new_AGEMA_signal_2392), .B1_f (new_AGEMA_signal_2393), .Z0_t (SubCellInst_SboxInst_6_Q7), .Z0_f (new_AGEMA_signal_2906), .Z1_t (new_AGEMA_signal_2907), .Z1_f (new_AGEMA_signal_2908) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_AND4_U1 ( .A0_t (SubCellInst_SboxInst_6_Q6), .A0_f (new_AGEMA_signal_2394), .A1_t (new_AGEMA_signal_2395), .A1_f (new_AGEMA_signal_2396), .B0_t (SubCellInst_SboxInst_6_Q7), .B0_f (new_AGEMA_signal_2906), .B1_t (new_AGEMA_signal_2907), .B1_f (new_AGEMA_signal_2908), .Z0_t (SubCellInst_SboxInst_6_T3), .Z0_f (new_AGEMA_signal_3095), .Z1_t (new_AGEMA_signal_3096), .Z1_f (new_AGEMA_signal_3097) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR8_U1 ( .A0_t (Ciphertext_s0_t[25]), .A0_f (Ciphertext_s0_f[25]), .A1_t (Ciphertext_s1_t[25]), .A1_f (Ciphertext_s1_f[25]), .B0_t (Ciphertext_s0_t[26]), .B0_f (Ciphertext_s0_f[26]), .B1_t (Ciphertext_s1_t[26]), .B1_f (Ciphertext_s1_f[26]), .Z0_t (SubCellInst_SboxInst_6_L2), .Z0_f (new_AGEMA_signal_1504), .Z1_t (new_AGEMA_signal_1505), .Z1_f (new_AGEMA_signal_1506) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_6_L0), .A0_f (new_AGEMA_signal_3293), .A1_t (new_AGEMA_signal_3294), .A1_f (new_AGEMA_signal_3295), .B0_t (SubCellInst_SboxInst_6_L2), .B0_f (new_AGEMA_signal_1504), .B1_t (new_AGEMA_signal_1505), .B1_f (new_AGEMA_signal_1506), .Z0_t (SubCellInst_SboxInst_6_YY_3), .Z0_f (new_AGEMA_signal_3465), .Z1_t (new_AGEMA_signal_3466), .Z1_f (new_AGEMA_signal_3467) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_6_L0), .A0_f (new_AGEMA_signal_3293), .A1_t (new_AGEMA_signal_3294), .A1_f (new_AGEMA_signal_3295), .B0_t (SubCellInst_SboxInst_6_T3), .B0_f (new_AGEMA_signal_3095), .B1_t (new_AGEMA_signal_3096), .B1_f (new_AGEMA_signal_3097), .Z0_t (ShiftRowsOutput[16]), .Z0_f (new_AGEMA_signal_3468), .Z1_t (new_AGEMA_signal_3469), .Z1_f (new_AGEMA_signal_3470) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_6_XX[2]), .A0_f (new_AGEMA_signal_1495), .A1_t (new_AGEMA_signal_1496), .A1_f (new_AGEMA_signal_1497), .B0_t (SubCellInst_SboxInst_6_T0), .B0_f (new_AGEMA_signal_2755), .B1_t (new_AGEMA_signal_2756), .B1_f (new_AGEMA_signal_2757), .Z0_t (SubCellInst_SboxInst_6_L3), .Z0_f (new_AGEMA_signal_2909), .Z1_t (new_AGEMA_signal_2910), .Z1_f (new_AGEMA_signal_2911) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_6_L3), .A0_f (new_AGEMA_signal_2909), .A1_t (new_AGEMA_signal_2910), .A1_f (new_AGEMA_signal_2911), .B0_t (SubCellInst_SboxInst_6_T2), .B0_f (new_AGEMA_signal_2391), .B1_t (new_AGEMA_signal_2392), .B1_f (new_AGEMA_signal_2393), .Z0_t (SubCellInst_SboxInst_6_YY[1]), .Z0_f (new_AGEMA_signal_3098), .Z1_t (new_AGEMA_signal_3099), .Z1_f (new_AGEMA_signal_3100) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_6_XX[1]), .A0_f (new_AGEMA_signal_1489), .A1_t (new_AGEMA_signal_1490), .A1_f (new_AGEMA_signal_1491), .B0_t (SubCellInst_SboxInst_6_T2), .B0_f (new_AGEMA_signal_2391), .B1_t (new_AGEMA_signal_2392), .B1_f (new_AGEMA_signal_2393), .Z0_t (SubCellInst_SboxInst_6_YY[0]), .Z0_f (new_AGEMA_signal_2761), .Z1_t (new_AGEMA_signal_2762), .Z1_f (new_AGEMA_signal_2763) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_6_YY[1]), .A0_f (new_AGEMA_signal_3098), .A1_t (new_AGEMA_signal_3099), .A1_f (new_AGEMA_signal_3100), .B0_t (SubCellInst_SboxInst_6_YY_3), .B0_f (new_AGEMA_signal_3465), .B1_t (new_AGEMA_signal_3466), .B1_f (new_AGEMA_signal_3467), .Z0_t (ShiftRowsOutput[17]), .Z0_f (new_AGEMA_signal_3654), .Z1_t (new_AGEMA_signal_3655), .Z1_f (new_AGEMA_signal_3656) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[30]), .A0_f (Ciphertext_s0_f[30]), .A1_t (Ciphertext_s1_t[30]), .A1_f (Ciphertext_s1_f[30]), .B0_t (Ciphertext_s0_t[31]), .B0_f (Ciphertext_s0_f[31]), .B1_t (Ciphertext_s1_t[31]), .B1_f (Ciphertext_s1_f[31]), .Z0_t (SubCellInst_SboxInst_7_XX[1]), .Z0_f (new_AGEMA_signal_1513), .Z1_t (new_AGEMA_signal_1514), .Z1_f (new_AGEMA_signal_1515) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[28]), .A0_f (Ciphertext_s0_f[28]), .A1_t (Ciphertext_s1_t[28]), .A1_f (Ciphertext_s1_f[28]), .B0_t (Ciphertext_s0_t[30]), .B0_f (Ciphertext_s0_f[30]), .B1_t (Ciphertext_s1_t[30]), .B1_f (Ciphertext_s1_f[30]), .Z0_t (SubCellInst_SboxInst_7_XX[2]), .Z0_f (new_AGEMA_signal_1519), .Z1_t (new_AGEMA_signal_1520), .Z1_f (new_AGEMA_signal_1521) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR0_U1 ( .A0_t (Ciphertext_s0_t[29]), .A0_f (Ciphertext_s0_f[29]), .A1_t (Ciphertext_s1_t[29]), .A1_f (Ciphertext_s1_f[29]), .B0_t (SubCellInst_SboxInst_7_XX[2]), .B0_f (new_AGEMA_signal_1519), .B1_t (new_AGEMA_signal_1520), .B1_f (new_AGEMA_signal_1521), .Z0_t (SubCellInst_SboxInst_7_Q0), .Z0_f (new_AGEMA_signal_2397), .Z1_t (new_AGEMA_signal_2398), .Z1_f (new_AGEMA_signal_2399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR1_U1 ( .A0_t (Ciphertext_s0_t[29]), .A0_f (Ciphertext_s0_f[29]), .A1_t (Ciphertext_s1_t[29]), .A1_f (Ciphertext_s1_f[29]), .B0_t (SubCellInst_SboxInst_7_XX[1]), .B0_f (new_AGEMA_signal_1513), .B1_t (new_AGEMA_signal_1514), .B1_f (new_AGEMA_signal_1515), .Z0_t (SubCellInst_SboxInst_7_Q1), .Z0_f (new_AGEMA_signal_2400), .Z1_t (new_AGEMA_signal_2401), .Z1_f (new_AGEMA_signal_2402) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_AND1_U1 ( .A0_t (Ciphertext_s0_t[30]), .A0_f (Ciphertext_s0_f[30]), .A1_t (Ciphertext_s1_t[30]), .A1_f (Ciphertext_s1_f[30]), .B0_t (SubCellInst_SboxInst_7_Q1), .B0_f (new_AGEMA_signal_2400), .B1_t (new_AGEMA_signal_2401), .B1_f (new_AGEMA_signal_2402), .Z0_t (SubCellInst_SboxInst_7_T0), .Z0_f (new_AGEMA_signal_2764), .Z1_t (new_AGEMA_signal_2765), .Z1_f (new_AGEMA_signal_2766) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_7_Q0), .A0_f (new_AGEMA_signal_2397), .A1_t (new_AGEMA_signal_2398), .A1_f (new_AGEMA_signal_2399), .B0_t (SubCellInst_SboxInst_7_T0), .B0_f (new_AGEMA_signal_2764), .B1_t (new_AGEMA_signal_2765), .B1_f (new_AGEMA_signal_2766), .Z0_t (SubCellInst_SboxInst_7_Q2), .Z0_f (new_AGEMA_signal_2912), .Z1_t (new_AGEMA_signal_2913), .Z1_f (new_AGEMA_signal_2914) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_AND2_U1 ( .A0_t (Ciphertext_s0_t[29]), .A0_f (Ciphertext_s0_f[29]), .A1_t (Ciphertext_s1_t[29]), .A1_f (Ciphertext_s1_f[29]), .B0_t (SubCellInst_SboxInst_7_Q2), .B0_f (new_AGEMA_signal_2912), .B1_t (new_AGEMA_signal_2913), .B1_f (new_AGEMA_signal_2914), .Z0_t (SubCellInst_SboxInst_7_T1), .Z0_f (new_AGEMA_signal_3101), .Z1_t (new_AGEMA_signal_3102), .Z1_f (new_AGEMA_signal_3103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_XOR3_U1 ( .A0_t (Ciphertext_s0_t[29]), .A0_f (Ciphertext_s0_f[29]), .A1_t (Ciphertext_s1_t[29]), .A1_f (Ciphertext_s1_f[29]), .B0_t (Ciphertext_s0_t[30]), .B0_f (Ciphertext_s0_f[30]), .B1_t (Ciphertext_s1_t[30]), .B1_f (Ciphertext_s1_f[30]), .Z0_t (SubCellInst_SboxInst_7_Q4), .Z0_f (new_AGEMA_signal_1525), .Z1_t (new_AGEMA_signal_1526), .Z1_f (new_AGEMA_signal_1527) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_AND3_U1 ( .A0_t (Ciphertext_s0_t[30]), .A0_f (Ciphertext_s0_f[30]), .A1_t (Ciphertext_s1_t[30]), .A1_f (Ciphertext_s1_f[30]), .B0_t (SubCellInst_SboxInst_7_Q4), .B0_f (new_AGEMA_signal_1525), .B1_t (new_AGEMA_signal_1526), .B1_f (new_AGEMA_signal_1527), .Z0_t (SubCellInst_SboxInst_7_T2), .Z0_f (new_AGEMA_signal_2403), .Z1_t (new_AGEMA_signal_2404), .Z1_f (new_AGEMA_signal_2405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_7_T1), .A0_f (new_AGEMA_signal_3101), .A1_t (new_AGEMA_signal_3102), .A1_f (new_AGEMA_signal_3103), .B0_t (SubCellInst_SboxInst_7_T2), .B0_f (new_AGEMA_signal_2403), .B1_t (new_AGEMA_signal_2404), .B1_f (new_AGEMA_signal_2405), .Z0_t (SubCellInst_SboxInst_7_L0), .Z0_f (new_AGEMA_signal_3296), .Z1_t (new_AGEMA_signal_3297), .Z1_f (new_AGEMA_signal_3298) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_7_XX[2]), .A0_f (new_AGEMA_signal_1519), .A1_t (new_AGEMA_signal_1520), .A1_f (new_AGEMA_signal_1521), .B0_t (Ciphertext_s0_t[30]), .B0_f (Ciphertext_s0_f[30]), .B1_t (Ciphertext_s1_t[30]), .B1_f (Ciphertext_s1_f[30]), .Z0_t (SubCellInst_SboxInst_7_Q6), .Z0_f (new_AGEMA_signal_2406), .Z1_t (new_AGEMA_signal_2407), .Z1_f (new_AGEMA_signal_2408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_7_Q1), .A0_f (new_AGEMA_signal_2400), .A1_t (new_AGEMA_signal_2401), .A1_f (new_AGEMA_signal_2402), .B0_t (SubCellInst_SboxInst_7_Q6), .B0_f (new_AGEMA_signal_2406), .B1_t (new_AGEMA_signal_2407), .B1_f (new_AGEMA_signal_2408), .Z0_t (SubCellInst_SboxInst_7_L1), .Z0_f (new_AGEMA_signal_2767), .Z1_t (new_AGEMA_signal_2768), .Z1_f (new_AGEMA_signal_2769) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_7_L1), .A0_f (new_AGEMA_signal_2767), .A1_t (new_AGEMA_signal_2768), .A1_f (new_AGEMA_signal_2769), .B0_t (SubCellInst_SboxInst_7_T2), .B0_f (new_AGEMA_signal_2403), .B1_t (new_AGEMA_signal_2404), .B1_f (new_AGEMA_signal_2405), .Z0_t (SubCellInst_SboxInst_7_Q7), .Z0_f (new_AGEMA_signal_2915), .Z1_t (new_AGEMA_signal_2916), .Z1_f (new_AGEMA_signal_2917) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_AND4_U1 ( .A0_t (SubCellInst_SboxInst_7_Q6), .A0_f (new_AGEMA_signal_2406), .A1_t (new_AGEMA_signal_2407), .A1_f (new_AGEMA_signal_2408), .B0_t (SubCellInst_SboxInst_7_Q7), .B0_f (new_AGEMA_signal_2915), .B1_t (new_AGEMA_signal_2916), .B1_f (new_AGEMA_signal_2917), .Z0_t (SubCellInst_SboxInst_7_T3), .Z0_f (new_AGEMA_signal_3104), .Z1_t (new_AGEMA_signal_3105), .Z1_f (new_AGEMA_signal_3106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR8_U1 ( .A0_t (Ciphertext_s0_t[29]), .A0_f (Ciphertext_s0_f[29]), .A1_t (Ciphertext_s1_t[29]), .A1_f (Ciphertext_s1_f[29]), .B0_t (Ciphertext_s0_t[30]), .B0_f (Ciphertext_s0_f[30]), .B1_t (Ciphertext_s1_t[30]), .B1_f (Ciphertext_s1_f[30]), .Z0_t (SubCellInst_SboxInst_7_L2), .Z0_f (new_AGEMA_signal_1528), .Z1_t (new_AGEMA_signal_1529), .Z1_f (new_AGEMA_signal_1530) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_7_L0), .A0_f (new_AGEMA_signal_3296), .A1_t (new_AGEMA_signal_3297), .A1_f (new_AGEMA_signal_3298), .B0_t (SubCellInst_SboxInst_7_L2), .B0_f (new_AGEMA_signal_1528), .B1_t (new_AGEMA_signal_1529), .B1_f (new_AGEMA_signal_1530), .Z0_t (SubCellInst_SboxInst_7_YY_3), .Z0_f (new_AGEMA_signal_3471), .Z1_t (new_AGEMA_signal_3472), .Z1_f (new_AGEMA_signal_3473) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_7_L0), .A0_f (new_AGEMA_signal_3296), .A1_t (new_AGEMA_signal_3297), .A1_f (new_AGEMA_signal_3298), .B0_t (SubCellInst_SboxInst_7_T3), .B0_f (new_AGEMA_signal_3104), .B1_t (new_AGEMA_signal_3105), .B1_f (new_AGEMA_signal_3106), .Z0_t (ShiftRowsOutput[20]), .Z0_f (new_AGEMA_signal_3474), .Z1_t (new_AGEMA_signal_3475), .Z1_f (new_AGEMA_signal_3476) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_7_XX[2]), .A0_f (new_AGEMA_signal_1519), .A1_t (new_AGEMA_signal_1520), .A1_f (new_AGEMA_signal_1521), .B0_t (SubCellInst_SboxInst_7_T0), .B0_f (new_AGEMA_signal_2764), .B1_t (new_AGEMA_signal_2765), .B1_f (new_AGEMA_signal_2766), .Z0_t (SubCellInst_SboxInst_7_L3), .Z0_f (new_AGEMA_signal_2918), .Z1_t (new_AGEMA_signal_2919), .Z1_f (new_AGEMA_signal_2920) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_7_L3), .A0_f (new_AGEMA_signal_2918), .A1_t (new_AGEMA_signal_2919), .A1_f (new_AGEMA_signal_2920), .B0_t (SubCellInst_SboxInst_7_T2), .B0_f (new_AGEMA_signal_2403), .B1_t (new_AGEMA_signal_2404), .B1_f (new_AGEMA_signal_2405), .Z0_t (SubCellInst_SboxInst_7_YY[1]), .Z0_f (new_AGEMA_signal_3107), .Z1_t (new_AGEMA_signal_3108), .Z1_f (new_AGEMA_signal_3109) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_7_XX[1]), .A0_f (new_AGEMA_signal_1513), .A1_t (new_AGEMA_signal_1514), .A1_f (new_AGEMA_signal_1515), .B0_t (SubCellInst_SboxInst_7_T2), .B0_f (new_AGEMA_signal_2403), .B1_t (new_AGEMA_signal_2404), .B1_f (new_AGEMA_signal_2405), .Z0_t (SubCellInst_SboxInst_7_YY[0]), .Z0_f (new_AGEMA_signal_2770), .Z1_t (new_AGEMA_signal_2771), .Z1_f (new_AGEMA_signal_2772) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_7_YY[1]), .A0_f (new_AGEMA_signal_3107), .A1_t (new_AGEMA_signal_3108), .A1_f (new_AGEMA_signal_3109), .B0_t (SubCellInst_SboxInst_7_YY_3), .B0_f (new_AGEMA_signal_3471), .B1_t (new_AGEMA_signal_3472), .B1_f (new_AGEMA_signal_3473), .Z0_t (SubCellOutput[29]), .Z0_f (new_AGEMA_signal_3657), .Z1_t (new_AGEMA_signal_3658), .Z1_f (new_AGEMA_signal_3659) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[34]), .A0_f (Ciphertext_s0_f[34]), .A1_t (Ciphertext_s1_t[34]), .A1_f (Ciphertext_s1_f[34]), .B0_t (Ciphertext_s0_t[35]), .B0_f (Ciphertext_s0_f[35]), .B1_t (Ciphertext_s1_t[35]), .B1_f (Ciphertext_s1_f[35]), .Z0_t (SubCellInst_SboxInst_8_XX[1]), .Z0_f (new_AGEMA_signal_1537), .Z1_t (new_AGEMA_signal_1538), .Z1_f (new_AGEMA_signal_1539) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[32]), .A0_f (Ciphertext_s0_f[32]), .A1_t (Ciphertext_s1_t[32]), .A1_f (Ciphertext_s1_f[32]), .B0_t (Ciphertext_s0_t[34]), .B0_f (Ciphertext_s0_f[34]), .B1_t (Ciphertext_s1_t[34]), .B1_f (Ciphertext_s1_f[34]), .Z0_t (SubCellInst_SboxInst_8_XX[2]), .Z0_f (new_AGEMA_signal_1543), .Z1_t (new_AGEMA_signal_1544), .Z1_f (new_AGEMA_signal_1545) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR0_U1 ( .A0_t (Ciphertext_s0_t[33]), .A0_f (Ciphertext_s0_f[33]), .A1_t (Ciphertext_s1_t[33]), .A1_f (Ciphertext_s1_f[33]), .B0_t (SubCellInst_SboxInst_8_XX[2]), .B0_f (new_AGEMA_signal_1543), .B1_t (new_AGEMA_signal_1544), .B1_f (new_AGEMA_signal_1545), .Z0_t (SubCellInst_SboxInst_8_Q0), .Z0_f (new_AGEMA_signal_2409), .Z1_t (new_AGEMA_signal_2410), .Z1_f (new_AGEMA_signal_2411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR1_U1 ( .A0_t (Ciphertext_s0_t[33]), .A0_f (Ciphertext_s0_f[33]), .A1_t (Ciphertext_s1_t[33]), .A1_f (Ciphertext_s1_f[33]), .B0_t (SubCellInst_SboxInst_8_XX[1]), .B0_f (new_AGEMA_signal_1537), .B1_t (new_AGEMA_signal_1538), .B1_f (new_AGEMA_signal_1539), .Z0_t (SubCellInst_SboxInst_8_Q1), .Z0_f (new_AGEMA_signal_2412), .Z1_t (new_AGEMA_signal_2413), .Z1_f (new_AGEMA_signal_2414) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_AND1_U1 ( .A0_t (Ciphertext_s0_t[34]), .A0_f (Ciphertext_s0_f[34]), .A1_t (Ciphertext_s1_t[34]), .A1_f (Ciphertext_s1_f[34]), .B0_t (SubCellInst_SboxInst_8_Q1), .B0_f (new_AGEMA_signal_2412), .B1_t (new_AGEMA_signal_2413), .B1_f (new_AGEMA_signal_2414), .Z0_t (SubCellInst_SboxInst_8_T0), .Z0_f (new_AGEMA_signal_2773), .Z1_t (new_AGEMA_signal_2774), .Z1_f (new_AGEMA_signal_2775) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_8_Q0), .A0_f (new_AGEMA_signal_2409), .A1_t (new_AGEMA_signal_2410), .A1_f (new_AGEMA_signal_2411), .B0_t (SubCellInst_SboxInst_8_T0), .B0_f (new_AGEMA_signal_2773), .B1_t (new_AGEMA_signal_2774), .B1_f (new_AGEMA_signal_2775), .Z0_t (SubCellInst_SboxInst_8_Q2), .Z0_f (new_AGEMA_signal_2921), .Z1_t (new_AGEMA_signal_2922), .Z1_f (new_AGEMA_signal_2923) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_AND2_U1 ( .A0_t (Ciphertext_s0_t[33]), .A0_f (Ciphertext_s0_f[33]), .A1_t (Ciphertext_s1_t[33]), .A1_f (Ciphertext_s1_f[33]), .B0_t (SubCellInst_SboxInst_8_Q2), .B0_f (new_AGEMA_signal_2921), .B1_t (new_AGEMA_signal_2922), .B1_f (new_AGEMA_signal_2923), .Z0_t (SubCellInst_SboxInst_8_T1), .Z0_f (new_AGEMA_signal_3110), .Z1_t (new_AGEMA_signal_3111), .Z1_f (new_AGEMA_signal_3112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_XOR3_U1 ( .A0_t (Ciphertext_s0_t[33]), .A0_f (Ciphertext_s0_f[33]), .A1_t (Ciphertext_s1_t[33]), .A1_f (Ciphertext_s1_f[33]), .B0_t (Ciphertext_s0_t[34]), .B0_f (Ciphertext_s0_f[34]), .B1_t (Ciphertext_s1_t[34]), .B1_f (Ciphertext_s1_f[34]), .Z0_t (SubCellInst_SboxInst_8_Q4), .Z0_f (new_AGEMA_signal_1549), .Z1_t (new_AGEMA_signal_1550), .Z1_f (new_AGEMA_signal_1551) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_AND3_U1 ( .A0_t (Ciphertext_s0_t[34]), .A0_f (Ciphertext_s0_f[34]), .A1_t (Ciphertext_s1_t[34]), .A1_f (Ciphertext_s1_f[34]), .B0_t (SubCellInst_SboxInst_8_Q4), .B0_f (new_AGEMA_signal_1549), .B1_t (new_AGEMA_signal_1550), .B1_f (new_AGEMA_signal_1551), .Z0_t (SubCellInst_SboxInst_8_T2), .Z0_f (new_AGEMA_signal_2415), .Z1_t (new_AGEMA_signal_2416), .Z1_f (new_AGEMA_signal_2417) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_8_T1), .A0_f (new_AGEMA_signal_3110), .A1_t (new_AGEMA_signal_3111), .A1_f (new_AGEMA_signal_3112), .B0_t (SubCellInst_SboxInst_8_T2), .B0_f (new_AGEMA_signal_2415), .B1_t (new_AGEMA_signal_2416), .B1_f (new_AGEMA_signal_2417), .Z0_t (SubCellInst_SboxInst_8_L0), .Z0_f (new_AGEMA_signal_3299), .Z1_t (new_AGEMA_signal_3300), .Z1_f (new_AGEMA_signal_3301) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_8_XX[2]), .A0_f (new_AGEMA_signal_1543), .A1_t (new_AGEMA_signal_1544), .A1_f (new_AGEMA_signal_1545), .B0_t (Ciphertext_s0_t[34]), .B0_f (Ciphertext_s0_f[34]), .B1_t (Ciphertext_s1_t[34]), .B1_f (Ciphertext_s1_f[34]), .Z0_t (SubCellInst_SboxInst_8_Q6), .Z0_f (new_AGEMA_signal_2418), .Z1_t (new_AGEMA_signal_2419), .Z1_f (new_AGEMA_signal_2420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_8_Q1), .A0_f (new_AGEMA_signal_2412), .A1_t (new_AGEMA_signal_2413), .A1_f (new_AGEMA_signal_2414), .B0_t (SubCellInst_SboxInst_8_Q6), .B0_f (new_AGEMA_signal_2418), .B1_t (new_AGEMA_signal_2419), .B1_f (new_AGEMA_signal_2420), .Z0_t (SubCellInst_SboxInst_8_L1), .Z0_f (new_AGEMA_signal_2776), .Z1_t (new_AGEMA_signal_2777), .Z1_f (new_AGEMA_signal_2778) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_8_L1), .A0_f (new_AGEMA_signal_2776), .A1_t (new_AGEMA_signal_2777), .A1_f (new_AGEMA_signal_2778), .B0_t (SubCellInst_SboxInst_8_T2), .B0_f (new_AGEMA_signal_2415), .B1_t (new_AGEMA_signal_2416), .B1_f (new_AGEMA_signal_2417), .Z0_t (SubCellInst_SboxInst_8_Q7), .Z0_f (new_AGEMA_signal_2924), .Z1_t (new_AGEMA_signal_2925), .Z1_f (new_AGEMA_signal_2926) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_AND4_U1 ( .A0_t (SubCellInst_SboxInst_8_Q6), .A0_f (new_AGEMA_signal_2418), .A1_t (new_AGEMA_signal_2419), .A1_f (new_AGEMA_signal_2420), .B0_t (SubCellInst_SboxInst_8_Q7), .B0_f (new_AGEMA_signal_2924), .B1_t (new_AGEMA_signal_2925), .B1_f (new_AGEMA_signal_2926), .Z0_t (SubCellInst_SboxInst_8_T3), .Z0_f (new_AGEMA_signal_3113), .Z1_t (new_AGEMA_signal_3114), .Z1_f (new_AGEMA_signal_3115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR8_U1 ( .A0_t (Ciphertext_s0_t[33]), .A0_f (Ciphertext_s0_f[33]), .A1_t (Ciphertext_s1_t[33]), .A1_f (Ciphertext_s1_f[33]), .B0_t (Ciphertext_s0_t[34]), .B0_f (Ciphertext_s0_f[34]), .B1_t (Ciphertext_s1_t[34]), .B1_f (Ciphertext_s1_f[34]), .Z0_t (SubCellInst_SboxInst_8_L2), .Z0_f (new_AGEMA_signal_1552), .Z1_t (new_AGEMA_signal_1553), .Z1_f (new_AGEMA_signal_1554) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_8_L0), .A0_f (new_AGEMA_signal_3299), .A1_t (new_AGEMA_signal_3300), .A1_f (new_AGEMA_signal_3301), .B0_t (SubCellInst_SboxInst_8_L2), .B0_f (new_AGEMA_signal_1552), .B1_t (new_AGEMA_signal_1553), .B1_f (new_AGEMA_signal_1554), .Z0_t (SubCellInst_SboxInst_8_YY_3), .Z0_f (new_AGEMA_signal_3477), .Z1_t (new_AGEMA_signal_3478), .Z1_f (new_AGEMA_signal_3479) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_8_L0), .A0_f (new_AGEMA_signal_3299), .A1_t (new_AGEMA_signal_3300), .A1_f (new_AGEMA_signal_3301), .B0_t (SubCellInst_SboxInst_8_T3), .B0_f (new_AGEMA_signal_3113), .B1_t (new_AGEMA_signal_3114), .B1_f (new_AGEMA_signal_3115), .Z0_t (AddRoundConstantOutput[32]), .Z0_f (new_AGEMA_signal_3480), .Z1_t (new_AGEMA_signal_3481), .Z1_f (new_AGEMA_signal_3482) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_8_XX[2]), .A0_f (new_AGEMA_signal_1543), .A1_t (new_AGEMA_signal_1544), .A1_f (new_AGEMA_signal_1545), .B0_t (SubCellInst_SboxInst_8_T0), .B0_f (new_AGEMA_signal_2773), .B1_t (new_AGEMA_signal_2774), .B1_f (new_AGEMA_signal_2775), .Z0_t (SubCellInst_SboxInst_8_L3), .Z0_f (new_AGEMA_signal_2927), .Z1_t (new_AGEMA_signal_2928), .Z1_f (new_AGEMA_signal_2929) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_8_L3), .A0_f (new_AGEMA_signal_2927), .A1_t (new_AGEMA_signal_2928), .A1_f (new_AGEMA_signal_2929), .B0_t (SubCellInst_SboxInst_8_T2), .B0_f (new_AGEMA_signal_2415), .B1_t (new_AGEMA_signal_2416), .B1_f (new_AGEMA_signal_2417), .Z0_t (SubCellInst_SboxInst_8_YY[1]), .Z0_f (new_AGEMA_signal_3116), .Z1_t (new_AGEMA_signal_3117), .Z1_f (new_AGEMA_signal_3118) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_8_XX[1]), .A0_f (new_AGEMA_signal_1537), .A1_t (new_AGEMA_signal_1538), .A1_f (new_AGEMA_signal_1539), .B0_t (SubCellInst_SboxInst_8_T2), .B0_f (new_AGEMA_signal_2415), .B1_t (new_AGEMA_signal_2416), .B1_f (new_AGEMA_signal_2417), .Z0_t (SubCellInst_SboxInst_8_YY[0]), .Z0_f (new_AGEMA_signal_2779), .Z1_t (new_AGEMA_signal_2780), .Z1_f (new_AGEMA_signal_2781) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_8_YY[1]), .A0_f (new_AGEMA_signal_3116), .A1_t (new_AGEMA_signal_3117), .A1_f (new_AGEMA_signal_3118), .B0_t (SubCellInst_SboxInst_8_YY_3), .B0_f (new_AGEMA_signal_3477), .B1_t (new_AGEMA_signal_3478), .B1_f (new_AGEMA_signal_3479), .Z0_t (AddRoundConstantOutput[33]), .Z0_f (new_AGEMA_signal_3660), .Z1_t (new_AGEMA_signal_3661), .Z1_f (new_AGEMA_signal_3662) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[38]), .A0_f (Ciphertext_s0_f[38]), .A1_t (Ciphertext_s1_t[38]), .A1_f (Ciphertext_s1_f[38]), .B0_t (Ciphertext_s0_t[39]), .B0_f (Ciphertext_s0_f[39]), .B1_t (Ciphertext_s1_t[39]), .B1_f (Ciphertext_s1_f[39]), .Z0_t (SubCellInst_SboxInst_9_XX[1]), .Z0_f (new_AGEMA_signal_1561), .Z1_t (new_AGEMA_signal_1562), .Z1_f (new_AGEMA_signal_1563) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[36]), .A0_f (Ciphertext_s0_f[36]), .A1_t (Ciphertext_s1_t[36]), .A1_f (Ciphertext_s1_f[36]), .B0_t (Ciphertext_s0_t[38]), .B0_f (Ciphertext_s0_f[38]), .B1_t (Ciphertext_s1_t[38]), .B1_f (Ciphertext_s1_f[38]), .Z0_t (SubCellInst_SboxInst_9_XX[2]), .Z0_f (new_AGEMA_signal_1567), .Z1_t (new_AGEMA_signal_1568), .Z1_f (new_AGEMA_signal_1569) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR0_U1 ( .A0_t (Ciphertext_s0_t[37]), .A0_f (Ciphertext_s0_f[37]), .A1_t (Ciphertext_s1_t[37]), .A1_f (Ciphertext_s1_f[37]), .B0_t (SubCellInst_SboxInst_9_XX[2]), .B0_f (new_AGEMA_signal_1567), .B1_t (new_AGEMA_signal_1568), .B1_f (new_AGEMA_signal_1569), .Z0_t (SubCellInst_SboxInst_9_Q0), .Z0_f (new_AGEMA_signal_2421), .Z1_t (new_AGEMA_signal_2422), .Z1_f (new_AGEMA_signal_2423) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR1_U1 ( .A0_t (Ciphertext_s0_t[37]), .A0_f (Ciphertext_s0_f[37]), .A1_t (Ciphertext_s1_t[37]), .A1_f (Ciphertext_s1_f[37]), .B0_t (SubCellInst_SboxInst_9_XX[1]), .B0_f (new_AGEMA_signal_1561), .B1_t (new_AGEMA_signal_1562), .B1_f (new_AGEMA_signal_1563), .Z0_t (SubCellInst_SboxInst_9_Q1), .Z0_f (new_AGEMA_signal_2424), .Z1_t (new_AGEMA_signal_2425), .Z1_f (new_AGEMA_signal_2426) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_AND1_U1 ( .A0_t (Ciphertext_s0_t[38]), .A0_f (Ciphertext_s0_f[38]), .A1_t (Ciphertext_s1_t[38]), .A1_f (Ciphertext_s1_f[38]), .B0_t (SubCellInst_SboxInst_9_Q1), .B0_f (new_AGEMA_signal_2424), .B1_t (new_AGEMA_signal_2425), .B1_f (new_AGEMA_signal_2426), .Z0_t (SubCellInst_SboxInst_9_T0), .Z0_f (new_AGEMA_signal_2782), .Z1_t (new_AGEMA_signal_2783), .Z1_f (new_AGEMA_signal_2784) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_9_Q0), .A0_f (new_AGEMA_signal_2421), .A1_t (new_AGEMA_signal_2422), .A1_f (new_AGEMA_signal_2423), .B0_t (SubCellInst_SboxInst_9_T0), .B0_f (new_AGEMA_signal_2782), .B1_t (new_AGEMA_signal_2783), .B1_f (new_AGEMA_signal_2784), .Z0_t (SubCellInst_SboxInst_9_Q2), .Z0_f (new_AGEMA_signal_2930), .Z1_t (new_AGEMA_signal_2931), .Z1_f (new_AGEMA_signal_2932) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_AND2_U1 ( .A0_t (Ciphertext_s0_t[37]), .A0_f (Ciphertext_s0_f[37]), .A1_t (Ciphertext_s1_t[37]), .A1_f (Ciphertext_s1_f[37]), .B0_t (SubCellInst_SboxInst_9_Q2), .B0_f (new_AGEMA_signal_2930), .B1_t (new_AGEMA_signal_2931), .B1_f (new_AGEMA_signal_2932), .Z0_t (SubCellInst_SboxInst_9_T1), .Z0_f (new_AGEMA_signal_3119), .Z1_t (new_AGEMA_signal_3120), .Z1_f (new_AGEMA_signal_3121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_XOR3_U1 ( .A0_t (Ciphertext_s0_t[37]), .A0_f (Ciphertext_s0_f[37]), .A1_t (Ciphertext_s1_t[37]), .A1_f (Ciphertext_s1_f[37]), .B0_t (Ciphertext_s0_t[38]), .B0_f (Ciphertext_s0_f[38]), .B1_t (Ciphertext_s1_t[38]), .B1_f (Ciphertext_s1_f[38]), .Z0_t (SubCellInst_SboxInst_9_Q4), .Z0_f (new_AGEMA_signal_1573), .Z1_t (new_AGEMA_signal_1574), .Z1_f (new_AGEMA_signal_1575) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_AND3_U1 ( .A0_t (Ciphertext_s0_t[38]), .A0_f (Ciphertext_s0_f[38]), .A1_t (Ciphertext_s1_t[38]), .A1_f (Ciphertext_s1_f[38]), .B0_t (SubCellInst_SboxInst_9_Q4), .B0_f (new_AGEMA_signal_1573), .B1_t (new_AGEMA_signal_1574), .B1_f (new_AGEMA_signal_1575), .Z0_t (SubCellInst_SboxInst_9_T2), .Z0_f (new_AGEMA_signal_2427), .Z1_t (new_AGEMA_signal_2428), .Z1_f (new_AGEMA_signal_2429) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_9_T1), .A0_f (new_AGEMA_signal_3119), .A1_t (new_AGEMA_signal_3120), .A1_f (new_AGEMA_signal_3121), .B0_t (SubCellInst_SboxInst_9_T2), .B0_f (new_AGEMA_signal_2427), .B1_t (new_AGEMA_signal_2428), .B1_f (new_AGEMA_signal_2429), .Z0_t (SubCellInst_SboxInst_9_L0), .Z0_f (new_AGEMA_signal_3302), .Z1_t (new_AGEMA_signal_3303), .Z1_f (new_AGEMA_signal_3304) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_9_XX[2]), .A0_f (new_AGEMA_signal_1567), .A1_t (new_AGEMA_signal_1568), .A1_f (new_AGEMA_signal_1569), .B0_t (Ciphertext_s0_t[38]), .B0_f (Ciphertext_s0_f[38]), .B1_t (Ciphertext_s1_t[38]), .B1_f (Ciphertext_s1_f[38]), .Z0_t (SubCellInst_SboxInst_9_Q6), .Z0_f (new_AGEMA_signal_2430), .Z1_t (new_AGEMA_signal_2431), .Z1_f (new_AGEMA_signal_2432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_9_Q1), .A0_f (new_AGEMA_signal_2424), .A1_t (new_AGEMA_signal_2425), .A1_f (new_AGEMA_signal_2426), .B0_t (SubCellInst_SboxInst_9_Q6), .B0_f (new_AGEMA_signal_2430), .B1_t (new_AGEMA_signal_2431), .B1_f (new_AGEMA_signal_2432), .Z0_t (SubCellInst_SboxInst_9_L1), .Z0_f (new_AGEMA_signal_2785), .Z1_t (new_AGEMA_signal_2786), .Z1_f (new_AGEMA_signal_2787) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_9_L1), .A0_f (new_AGEMA_signal_2785), .A1_t (new_AGEMA_signal_2786), .A1_f (new_AGEMA_signal_2787), .B0_t (SubCellInst_SboxInst_9_T2), .B0_f (new_AGEMA_signal_2427), .B1_t (new_AGEMA_signal_2428), .B1_f (new_AGEMA_signal_2429), .Z0_t (SubCellInst_SboxInst_9_Q7), .Z0_f (new_AGEMA_signal_2933), .Z1_t (new_AGEMA_signal_2934), .Z1_f (new_AGEMA_signal_2935) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_AND4_U1 ( .A0_t (SubCellInst_SboxInst_9_Q6), .A0_f (new_AGEMA_signal_2430), .A1_t (new_AGEMA_signal_2431), .A1_f (new_AGEMA_signal_2432), .B0_t (SubCellInst_SboxInst_9_Q7), .B0_f (new_AGEMA_signal_2933), .B1_t (new_AGEMA_signal_2934), .B1_f (new_AGEMA_signal_2935), .Z0_t (SubCellInst_SboxInst_9_T3), .Z0_f (new_AGEMA_signal_3122), .Z1_t (new_AGEMA_signal_3123), .Z1_f (new_AGEMA_signal_3124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR8_U1 ( .A0_t (Ciphertext_s0_t[37]), .A0_f (Ciphertext_s0_f[37]), .A1_t (Ciphertext_s1_t[37]), .A1_f (Ciphertext_s1_f[37]), .B0_t (Ciphertext_s0_t[38]), .B0_f (Ciphertext_s0_f[38]), .B1_t (Ciphertext_s1_t[38]), .B1_f (Ciphertext_s1_f[38]), .Z0_t (SubCellInst_SboxInst_9_L2), .Z0_f (new_AGEMA_signal_1576), .Z1_t (new_AGEMA_signal_1577), .Z1_f (new_AGEMA_signal_1578) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_9_L0), .A0_f (new_AGEMA_signal_3302), .A1_t (new_AGEMA_signal_3303), .A1_f (new_AGEMA_signal_3304), .B0_t (SubCellInst_SboxInst_9_L2), .B0_f (new_AGEMA_signal_1576), .B1_t (new_AGEMA_signal_1577), .B1_f (new_AGEMA_signal_1578), .Z0_t (SubCellInst_SboxInst_9_YY_3), .Z0_f (new_AGEMA_signal_3483), .Z1_t (new_AGEMA_signal_3484), .Z1_f (new_AGEMA_signal_3485) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_9_L0), .A0_f (new_AGEMA_signal_3302), .A1_t (new_AGEMA_signal_3303), .A1_f (new_AGEMA_signal_3304), .B0_t (SubCellInst_SboxInst_9_T3), .B0_f (new_AGEMA_signal_3122), .B1_t (new_AGEMA_signal_3123), .B1_f (new_AGEMA_signal_3124), .Z0_t (AddRoundConstantOutput[36]), .Z0_f (new_AGEMA_signal_3486), .Z1_t (new_AGEMA_signal_3487), .Z1_f (new_AGEMA_signal_3488) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_9_XX[2]), .A0_f (new_AGEMA_signal_1567), .A1_t (new_AGEMA_signal_1568), .A1_f (new_AGEMA_signal_1569), .B0_t (SubCellInst_SboxInst_9_T0), .B0_f (new_AGEMA_signal_2782), .B1_t (new_AGEMA_signal_2783), .B1_f (new_AGEMA_signal_2784), .Z0_t (SubCellInst_SboxInst_9_L3), .Z0_f (new_AGEMA_signal_2936), .Z1_t (new_AGEMA_signal_2937), .Z1_f (new_AGEMA_signal_2938) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_9_L3), .A0_f (new_AGEMA_signal_2936), .A1_t (new_AGEMA_signal_2937), .A1_f (new_AGEMA_signal_2938), .B0_t (SubCellInst_SboxInst_9_T2), .B0_f (new_AGEMA_signal_2427), .B1_t (new_AGEMA_signal_2428), .B1_f (new_AGEMA_signal_2429), .Z0_t (SubCellInst_SboxInst_9_YY[1]), .Z0_f (new_AGEMA_signal_3125), .Z1_t (new_AGEMA_signal_3126), .Z1_f (new_AGEMA_signal_3127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_9_XX[1]), .A0_f (new_AGEMA_signal_1561), .A1_t (new_AGEMA_signal_1562), .A1_f (new_AGEMA_signal_1563), .B0_t (SubCellInst_SboxInst_9_T2), .B0_f (new_AGEMA_signal_2427), .B1_t (new_AGEMA_signal_2428), .B1_f (new_AGEMA_signal_2429), .Z0_t (SubCellInst_SboxInst_9_YY[0]), .Z0_f (new_AGEMA_signal_2788), .Z1_t (new_AGEMA_signal_2789), .Z1_f (new_AGEMA_signal_2790) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_9_YY[1]), .A0_f (new_AGEMA_signal_3125), .A1_t (new_AGEMA_signal_3126), .A1_f (new_AGEMA_signal_3127), .B0_t (SubCellInst_SboxInst_9_YY_3), .B0_f (new_AGEMA_signal_3483), .B1_t (new_AGEMA_signal_3484), .B1_f (new_AGEMA_signal_3485), .Z0_t (AddRoundConstantOutput[37]), .Z0_f (new_AGEMA_signal_3663), .Z1_t (new_AGEMA_signal_3664), .Z1_f (new_AGEMA_signal_3665) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[42]), .A0_f (Ciphertext_s0_f[42]), .A1_t (Ciphertext_s1_t[42]), .A1_f (Ciphertext_s1_f[42]), .B0_t (Ciphertext_s0_t[43]), .B0_f (Ciphertext_s0_f[43]), .B1_t (Ciphertext_s1_t[43]), .B1_f (Ciphertext_s1_f[43]), .Z0_t (SubCellInst_SboxInst_10_XX[1]), .Z0_f (new_AGEMA_signal_1585), .Z1_t (new_AGEMA_signal_1586), .Z1_f (new_AGEMA_signal_1587) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[40]), .A0_f (Ciphertext_s0_f[40]), .A1_t (Ciphertext_s1_t[40]), .A1_f (Ciphertext_s1_f[40]), .B0_t (Ciphertext_s0_t[42]), .B0_f (Ciphertext_s0_f[42]), .B1_t (Ciphertext_s1_t[42]), .B1_f (Ciphertext_s1_f[42]), .Z0_t (SubCellInst_SboxInst_10_XX[2]), .Z0_f (new_AGEMA_signal_1591), .Z1_t (new_AGEMA_signal_1592), .Z1_f (new_AGEMA_signal_1593) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR0_U1 ( .A0_t (Ciphertext_s0_t[41]), .A0_f (Ciphertext_s0_f[41]), .A1_t (Ciphertext_s1_t[41]), .A1_f (Ciphertext_s1_f[41]), .B0_t (SubCellInst_SboxInst_10_XX[2]), .B0_f (new_AGEMA_signal_1591), .B1_t (new_AGEMA_signal_1592), .B1_f (new_AGEMA_signal_1593), .Z0_t (SubCellInst_SboxInst_10_Q0), .Z0_f (new_AGEMA_signal_2433), .Z1_t (new_AGEMA_signal_2434), .Z1_f (new_AGEMA_signal_2435) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR1_U1 ( .A0_t (Ciphertext_s0_t[41]), .A0_f (Ciphertext_s0_f[41]), .A1_t (Ciphertext_s1_t[41]), .A1_f (Ciphertext_s1_f[41]), .B0_t (SubCellInst_SboxInst_10_XX[1]), .B0_f (new_AGEMA_signal_1585), .B1_t (new_AGEMA_signal_1586), .B1_f (new_AGEMA_signal_1587), .Z0_t (SubCellInst_SboxInst_10_Q1), .Z0_f (new_AGEMA_signal_2436), .Z1_t (new_AGEMA_signal_2437), .Z1_f (new_AGEMA_signal_2438) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_AND1_U1 ( .A0_t (Ciphertext_s0_t[42]), .A0_f (Ciphertext_s0_f[42]), .A1_t (Ciphertext_s1_t[42]), .A1_f (Ciphertext_s1_f[42]), .B0_t (SubCellInst_SboxInst_10_Q1), .B0_f (new_AGEMA_signal_2436), .B1_t (new_AGEMA_signal_2437), .B1_f (new_AGEMA_signal_2438), .Z0_t (SubCellInst_SboxInst_10_T0), .Z0_f (new_AGEMA_signal_2791), .Z1_t (new_AGEMA_signal_2792), .Z1_f (new_AGEMA_signal_2793) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_10_Q0), .A0_f (new_AGEMA_signal_2433), .A1_t (new_AGEMA_signal_2434), .A1_f (new_AGEMA_signal_2435), .B0_t (SubCellInst_SboxInst_10_T0), .B0_f (new_AGEMA_signal_2791), .B1_t (new_AGEMA_signal_2792), .B1_f (new_AGEMA_signal_2793), .Z0_t (SubCellInst_SboxInst_10_Q2), .Z0_f (new_AGEMA_signal_2939), .Z1_t (new_AGEMA_signal_2940), .Z1_f (new_AGEMA_signal_2941) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_AND2_U1 ( .A0_t (Ciphertext_s0_t[41]), .A0_f (Ciphertext_s0_f[41]), .A1_t (Ciphertext_s1_t[41]), .A1_f (Ciphertext_s1_f[41]), .B0_t (SubCellInst_SboxInst_10_Q2), .B0_f (new_AGEMA_signal_2939), .B1_t (new_AGEMA_signal_2940), .B1_f (new_AGEMA_signal_2941), .Z0_t (SubCellInst_SboxInst_10_T1), .Z0_f (new_AGEMA_signal_3128), .Z1_t (new_AGEMA_signal_3129), .Z1_f (new_AGEMA_signal_3130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_XOR3_U1 ( .A0_t (Ciphertext_s0_t[41]), .A0_f (Ciphertext_s0_f[41]), .A1_t (Ciphertext_s1_t[41]), .A1_f (Ciphertext_s1_f[41]), .B0_t (Ciphertext_s0_t[42]), .B0_f (Ciphertext_s0_f[42]), .B1_t (Ciphertext_s1_t[42]), .B1_f (Ciphertext_s1_f[42]), .Z0_t (SubCellInst_SboxInst_10_Q4), .Z0_f (new_AGEMA_signal_1597), .Z1_t (new_AGEMA_signal_1598), .Z1_f (new_AGEMA_signal_1599) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_AND3_U1 ( .A0_t (Ciphertext_s0_t[42]), .A0_f (Ciphertext_s0_f[42]), .A1_t (Ciphertext_s1_t[42]), .A1_f (Ciphertext_s1_f[42]), .B0_t (SubCellInst_SboxInst_10_Q4), .B0_f (new_AGEMA_signal_1597), .B1_t (new_AGEMA_signal_1598), .B1_f (new_AGEMA_signal_1599), .Z0_t (SubCellInst_SboxInst_10_T2), .Z0_f (new_AGEMA_signal_2439), .Z1_t (new_AGEMA_signal_2440), .Z1_f (new_AGEMA_signal_2441) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_10_T1), .A0_f (new_AGEMA_signal_3128), .A1_t (new_AGEMA_signal_3129), .A1_f (new_AGEMA_signal_3130), .B0_t (SubCellInst_SboxInst_10_T2), .B0_f (new_AGEMA_signal_2439), .B1_t (new_AGEMA_signal_2440), .B1_f (new_AGEMA_signal_2441), .Z0_t (SubCellInst_SboxInst_10_L0), .Z0_f (new_AGEMA_signal_3305), .Z1_t (new_AGEMA_signal_3306), .Z1_f (new_AGEMA_signal_3307) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_10_XX[2]), .A0_f (new_AGEMA_signal_1591), .A1_t (new_AGEMA_signal_1592), .A1_f (new_AGEMA_signal_1593), .B0_t (Ciphertext_s0_t[42]), .B0_f (Ciphertext_s0_f[42]), .B1_t (Ciphertext_s1_t[42]), .B1_f (Ciphertext_s1_f[42]), .Z0_t (SubCellInst_SboxInst_10_Q6), .Z0_f (new_AGEMA_signal_2442), .Z1_t (new_AGEMA_signal_2443), .Z1_f (new_AGEMA_signal_2444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_10_Q1), .A0_f (new_AGEMA_signal_2436), .A1_t (new_AGEMA_signal_2437), .A1_f (new_AGEMA_signal_2438), .B0_t (SubCellInst_SboxInst_10_Q6), .B0_f (new_AGEMA_signal_2442), .B1_t (new_AGEMA_signal_2443), .B1_f (new_AGEMA_signal_2444), .Z0_t (SubCellInst_SboxInst_10_L1), .Z0_f (new_AGEMA_signal_2794), .Z1_t (new_AGEMA_signal_2795), .Z1_f (new_AGEMA_signal_2796) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_10_L1), .A0_f (new_AGEMA_signal_2794), .A1_t (new_AGEMA_signal_2795), .A1_f (new_AGEMA_signal_2796), .B0_t (SubCellInst_SboxInst_10_T2), .B0_f (new_AGEMA_signal_2439), .B1_t (new_AGEMA_signal_2440), .B1_f (new_AGEMA_signal_2441), .Z0_t (SubCellInst_SboxInst_10_Q7), .Z0_f (new_AGEMA_signal_2942), .Z1_t (new_AGEMA_signal_2943), .Z1_f (new_AGEMA_signal_2944) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_AND4_U1 ( .A0_t (SubCellInst_SboxInst_10_Q6), .A0_f (new_AGEMA_signal_2442), .A1_t (new_AGEMA_signal_2443), .A1_f (new_AGEMA_signal_2444), .B0_t (SubCellInst_SboxInst_10_Q7), .B0_f (new_AGEMA_signal_2942), .B1_t (new_AGEMA_signal_2943), .B1_f (new_AGEMA_signal_2944), .Z0_t (SubCellInst_SboxInst_10_T3), .Z0_f (new_AGEMA_signal_3131), .Z1_t (new_AGEMA_signal_3132), .Z1_f (new_AGEMA_signal_3133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR8_U1 ( .A0_t (Ciphertext_s0_t[41]), .A0_f (Ciphertext_s0_f[41]), .A1_t (Ciphertext_s1_t[41]), .A1_f (Ciphertext_s1_f[41]), .B0_t (Ciphertext_s0_t[42]), .B0_f (Ciphertext_s0_f[42]), .B1_t (Ciphertext_s1_t[42]), .B1_f (Ciphertext_s1_f[42]), .Z0_t (SubCellInst_SboxInst_10_L2), .Z0_f (new_AGEMA_signal_1600), .Z1_t (new_AGEMA_signal_1601), .Z1_f (new_AGEMA_signal_1602) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_10_L0), .A0_f (new_AGEMA_signal_3305), .A1_t (new_AGEMA_signal_3306), .A1_f (new_AGEMA_signal_3307), .B0_t (SubCellInst_SboxInst_10_L2), .B0_f (new_AGEMA_signal_1600), .B1_t (new_AGEMA_signal_1601), .B1_f (new_AGEMA_signal_1602), .Z0_t (SubCellInst_SboxInst_10_YY_3), .Z0_f (new_AGEMA_signal_3489), .Z1_t (new_AGEMA_signal_3490), .Z1_f (new_AGEMA_signal_3491) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_10_L0), .A0_f (new_AGEMA_signal_3305), .A1_t (new_AGEMA_signal_3306), .A1_f (new_AGEMA_signal_3307), .B0_t (SubCellInst_SboxInst_10_T3), .B0_f (new_AGEMA_signal_3131), .B1_t (new_AGEMA_signal_3132), .B1_f (new_AGEMA_signal_3133), .Z0_t (AddRoundConstantOutput[40]), .Z0_f (new_AGEMA_signal_3492), .Z1_t (new_AGEMA_signal_3493), .Z1_f (new_AGEMA_signal_3494) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_10_XX[2]), .A0_f (new_AGEMA_signal_1591), .A1_t (new_AGEMA_signal_1592), .A1_f (new_AGEMA_signal_1593), .B0_t (SubCellInst_SboxInst_10_T0), .B0_f (new_AGEMA_signal_2791), .B1_t (new_AGEMA_signal_2792), .B1_f (new_AGEMA_signal_2793), .Z0_t (SubCellInst_SboxInst_10_L3), .Z0_f (new_AGEMA_signal_2945), .Z1_t (new_AGEMA_signal_2946), .Z1_f (new_AGEMA_signal_2947) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_10_L3), .A0_f (new_AGEMA_signal_2945), .A1_t (new_AGEMA_signal_2946), .A1_f (new_AGEMA_signal_2947), .B0_t (SubCellInst_SboxInst_10_T2), .B0_f (new_AGEMA_signal_2439), .B1_t (new_AGEMA_signal_2440), .B1_f (new_AGEMA_signal_2441), .Z0_t (SubCellInst_SboxInst_10_YY[1]), .Z0_f (new_AGEMA_signal_3134), .Z1_t (new_AGEMA_signal_3135), .Z1_f (new_AGEMA_signal_3136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_10_XX[1]), .A0_f (new_AGEMA_signal_1585), .A1_t (new_AGEMA_signal_1586), .A1_f (new_AGEMA_signal_1587), .B0_t (SubCellInst_SboxInst_10_T2), .B0_f (new_AGEMA_signal_2439), .B1_t (new_AGEMA_signal_2440), .B1_f (new_AGEMA_signal_2441), .Z0_t (SubCellInst_SboxInst_10_YY[0]), .Z0_f (new_AGEMA_signal_2797), .Z1_t (new_AGEMA_signal_2798), .Z1_f (new_AGEMA_signal_2799) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_10_YY[1]), .A0_f (new_AGEMA_signal_3134), .A1_t (new_AGEMA_signal_3135), .A1_f (new_AGEMA_signal_3136), .B0_t (SubCellInst_SboxInst_10_YY_3), .B0_f (new_AGEMA_signal_3489), .B1_t (new_AGEMA_signal_3490), .B1_f (new_AGEMA_signal_3491), .Z0_t (AddRoundConstantOutput[41]), .Z0_f (new_AGEMA_signal_3666), .Z1_t (new_AGEMA_signal_3667), .Z1_f (new_AGEMA_signal_3668) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[46]), .A0_f (Ciphertext_s0_f[46]), .A1_t (Ciphertext_s1_t[46]), .A1_f (Ciphertext_s1_f[46]), .B0_t (Ciphertext_s0_t[47]), .B0_f (Ciphertext_s0_f[47]), .B1_t (Ciphertext_s1_t[47]), .B1_f (Ciphertext_s1_f[47]), .Z0_t (SubCellInst_SboxInst_11_XX[1]), .Z0_f (new_AGEMA_signal_1609), .Z1_t (new_AGEMA_signal_1610), .Z1_f (new_AGEMA_signal_1611) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[44]), .A0_f (Ciphertext_s0_f[44]), .A1_t (Ciphertext_s1_t[44]), .A1_f (Ciphertext_s1_f[44]), .B0_t (Ciphertext_s0_t[46]), .B0_f (Ciphertext_s0_f[46]), .B1_t (Ciphertext_s1_t[46]), .B1_f (Ciphertext_s1_f[46]), .Z0_t (SubCellInst_SboxInst_11_XX[2]), .Z0_f (new_AGEMA_signal_1615), .Z1_t (new_AGEMA_signal_1616), .Z1_f (new_AGEMA_signal_1617) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR0_U1 ( .A0_t (Ciphertext_s0_t[45]), .A0_f (Ciphertext_s0_f[45]), .A1_t (Ciphertext_s1_t[45]), .A1_f (Ciphertext_s1_f[45]), .B0_t (SubCellInst_SboxInst_11_XX[2]), .B0_f (new_AGEMA_signal_1615), .B1_t (new_AGEMA_signal_1616), .B1_f (new_AGEMA_signal_1617), .Z0_t (SubCellInst_SboxInst_11_Q0), .Z0_f (new_AGEMA_signal_2445), .Z1_t (new_AGEMA_signal_2446), .Z1_f (new_AGEMA_signal_2447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR1_U1 ( .A0_t (Ciphertext_s0_t[45]), .A0_f (Ciphertext_s0_f[45]), .A1_t (Ciphertext_s1_t[45]), .A1_f (Ciphertext_s1_f[45]), .B0_t (SubCellInst_SboxInst_11_XX[1]), .B0_f (new_AGEMA_signal_1609), .B1_t (new_AGEMA_signal_1610), .B1_f (new_AGEMA_signal_1611), .Z0_t (SubCellInst_SboxInst_11_Q1), .Z0_f (new_AGEMA_signal_2448), .Z1_t (new_AGEMA_signal_2449), .Z1_f (new_AGEMA_signal_2450) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_AND1_U1 ( .A0_t (Ciphertext_s0_t[46]), .A0_f (Ciphertext_s0_f[46]), .A1_t (Ciphertext_s1_t[46]), .A1_f (Ciphertext_s1_f[46]), .B0_t (SubCellInst_SboxInst_11_Q1), .B0_f (new_AGEMA_signal_2448), .B1_t (new_AGEMA_signal_2449), .B1_f (new_AGEMA_signal_2450), .Z0_t (SubCellInst_SboxInst_11_T0), .Z0_f (new_AGEMA_signal_2800), .Z1_t (new_AGEMA_signal_2801), .Z1_f (new_AGEMA_signal_2802) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_11_Q0), .A0_f (new_AGEMA_signal_2445), .A1_t (new_AGEMA_signal_2446), .A1_f (new_AGEMA_signal_2447), .B0_t (SubCellInst_SboxInst_11_T0), .B0_f (new_AGEMA_signal_2800), .B1_t (new_AGEMA_signal_2801), .B1_f (new_AGEMA_signal_2802), .Z0_t (SubCellInst_SboxInst_11_Q2), .Z0_f (new_AGEMA_signal_2948), .Z1_t (new_AGEMA_signal_2949), .Z1_f (new_AGEMA_signal_2950) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_AND2_U1 ( .A0_t (Ciphertext_s0_t[45]), .A0_f (Ciphertext_s0_f[45]), .A1_t (Ciphertext_s1_t[45]), .A1_f (Ciphertext_s1_f[45]), .B0_t (SubCellInst_SboxInst_11_Q2), .B0_f (new_AGEMA_signal_2948), .B1_t (new_AGEMA_signal_2949), .B1_f (new_AGEMA_signal_2950), .Z0_t (SubCellInst_SboxInst_11_T1), .Z0_f (new_AGEMA_signal_3137), .Z1_t (new_AGEMA_signal_3138), .Z1_f (new_AGEMA_signal_3139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_XOR3_U1 ( .A0_t (Ciphertext_s0_t[45]), .A0_f (Ciphertext_s0_f[45]), .A1_t (Ciphertext_s1_t[45]), .A1_f (Ciphertext_s1_f[45]), .B0_t (Ciphertext_s0_t[46]), .B0_f (Ciphertext_s0_f[46]), .B1_t (Ciphertext_s1_t[46]), .B1_f (Ciphertext_s1_f[46]), .Z0_t (SubCellInst_SboxInst_11_Q4), .Z0_f (new_AGEMA_signal_1621), .Z1_t (new_AGEMA_signal_1622), .Z1_f (new_AGEMA_signal_1623) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_AND3_U1 ( .A0_t (Ciphertext_s0_t[46]), .A0_f (Ciphertext_s0_f[46]), .A1_t (Ciphertext_s1_t[46]), .A1_f (Ciphertext_s1_f[46]), .B0_t (SubCellInst_SboxInst_11_Q4), .B0_f (new_AGEMA_signal_1621), .B1_t (new_AGEMA_signal_1622), .B1_f (new_AGEMA_signal_1623), .Z0_t (SubCellInst_SboxInst_11_T2), .Z0_f (new_AGEMA_signal_2451), .Z1_t (new_AGEMA_signal_2452), .Z1_f (new_AGEMA_signal_2453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_11_T1), .A0_f (new_AGEMA_signal_3137), .A1_t (new_AGEMA_signal_3138), .A1_f (new_AGEMA_signal_3139), .B0_t (SubCellInst_SboxInst_11_T2), .B0_f (new_AGEMA_signal_2451), .B1_t (new_AGEMA_signal_2452), .B1_f (new_AGEMA_signal_2453), .Z0_t (SubCellInst_SboxInst_11_L0), .Z0_f (new_AGEMA_signal_3308), .Z1_t (new_AGEMA_signal_3309), .Z1_f (new_AGEMA_signal_3310) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_11_XX[2]), .A0_f (new_AGEMA_signal_1615), .A1_t (new_AGEMA_signal_1616), .A1_f (new_AGEMA_signal_1617), .B0_t (Ciphertext_s0_t[46]), .B0_f (Ciphertext_s0_f[46]), .B1_t (Ciphertext_s1_t[46]), .B1_f (Ciphertext_s1_f[46]), .Z0_t (SubCellInst_SboxInst_11_Q6), .Z0_f (new_AGEMA_signal_2454), .Z1_t (new_AGEMA_signal_2455), .Z1_f (new_AGEMA_signal_2456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_11_Q1), .A0_f (new_AGEMA_signal_2448), .A1_t (new_AGEMA_signal_2449), .A1_f (new_AGEMA_signal_2450), .B0_t (SubCellInst_SboxInst_11_Q6), .B0_f (new_AGEMA_signal_2454), .B1_t (new_AGEMA_signal_2455), .B1_f (new_AGEMA_signal_2456), .Z0_t (SubCellInst_SboxInst_11_L1), .Z0_f (new_AGEMA_signal_2803), .Z1_t (new_AGEMA_signal_2804), .Z1_f (new_AGEMA_signal_2805) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_11_L1), .A0_f (new_AGEMA_signal_2803), .A1_t (new_AGEMA_signal_2804), .A1_f (new_AGEMA_signal_2805), .B0_t (SubCellInst_SboxInst_11_T2), .B0_f (new_AGEMA_signal_2451), .B1_t (new_AGEMA_signal_2452), .B1_f (new_AGEMA_signal_2453), .Z0_t (SubCellInst_SboxInst_11_Q7), .Z0_f (new_AGEMA_signal_2951), .Z1_t (new_AGEMA_signal_2952), .Z1_f (new_AGEMA_signal_2953) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_AND4_U1 ( .A0_t (SubCellInst_SboxInst_11_Q6), .A0_f (new_AGEMA_signal_2454), .A1_t (new_AGEMA_signal_2455), .A1_f (new_AGEMA_signal_2456), .B0_t (SubCellInst_SboxInst_11_Q7), .B0_f (new_AGEMA_signal_2951), .B1_t (new_AGEMA_signal_2952), .B1_f (new_AGEMA_signal_2953), .Z0_t (SubCellInst_SboxInst_11_T3), .Z0_f (new_AGEMA_signal_3140), .Z1_t (new_AGEMA_signal_3141), .Z1_f (new_AGEMA_signal_3142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR8_U1 ( .A0_t (Ciphertext_s0_t[45]), .A0_f (Ciphertext_s0_f[45]), .A1_t (Ciphertext_s1_t[45]), .A1_f (Ciphertext_s1_f[45]), .B0_t (Ciphertext_s0_t[46]), .B0_f (Ciphertext_s0_f[46]), .B1_t (Ciphertext_s1_t[46]), .B1_f (Ciphertext_s1_f[46]), .Z0_t (SubCellInst_SboxInst_11_L2), .Z0_f (new_AGEMA_signal_1624), .Z1_t (new_AGEMA_signal_1625), .Z1_f (new_AGEMA_signal_1626) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_11_L0), .A0_f (new_AGEMA_signal_3308), .A1_t (new_AGEMA_signal_3309), .A1_f (new_AGEMA_signal_3310), .B0_t (SubCellInst_SboxInst_11_L2), .B0_f (new_AGEMA_signal_1624), .B1_t (new_AGEMA_signal_1625), .B1_f (new_AGEMA_signal_1626), .Z0_t (SubCellInst_SboxInst_11_YY_3), .Z0_f (new_AGEMA_signal_3495), .Z1_t (new_AGEMA_signal_3496), .Z1_f (new_AGEMA_signal_3497) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_11_L0), .A0_f (new_AGEMA_signal_3308), .A1_t (new_AGEMA_signal_3309), .A1_f (new_AGEMA_signal_3310), .B0_t (SubCellInst_SboxInst_11_T3), .B0_f (new_AGEMA_signal_3140), .B1_t (new_AGEMA_signal_3141), .B1_f (new_AGEMA_signal_3142), .Z0_t (SubCellOutput[44]), .Z0_f (new_AGEMA_signal_3498), .Z1_t (new_AGEMA_signal_3499), .Z1_f (new_AGEMA_signal_3500) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_11_XX[2]), .A0_f (new_AGEMA_signal_1615), .A1_t (new_AGEMA_signal_1616), .A1_f (new_AGEMA_signal_1617), .B0_t (SubCellInst_SboxInst_11_T0), .B0_f (new_AGEMA_signal_2800), .B1_t (new_AGEMA_signal_2801), .B1_f (new_AGEMA_signal_2802), .Z0_t (SubCellInst_SboxInst_11_L3), .Z0_f (new_AGEMA_signal_2954), .Z1_t (new_AGEMA_signal_2955), .Z1_f (new_AGEMA_signal_2956) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_11_L3), .A0_f (new_AGEMA_signal_2954), .A1_t (new_AGEMA_signal_2955), .A1_f (new_AGEMA_signal_2956), .B0_t (SubCellInst_SboxInst_11_T2), .B0_f (new_AGEMA_signal_2451), .B1_t (new_AGEMA_signal_2452), .B1_f (new_AGEMA_signal_2453), .Z0_t (SubCellInst_SboxInst_11_YY[1]), .Z0_f (new_AGEMA_signal_3143), .Z1_t (new_AGEMA_signal_3144), .Z1_f (new_AGEMA_signal_3145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_11_XX[1]), .A0_f (new_AGEMA_signal_1609), .A1_t (new_AGEMA_signal_1610), .A1_f (new_AGEMA_signal_1611), .B0_t (SubCellInst_SboxInst_11_T2), .B0_f (new_AGEMA_signal_2451), .B1_t (new_AGEMA_signal_2452), .B1_f (new_AGEMA_signal_2453), .Z0_t (SubCellInst_SboxInst_11_YY[0]), .Z0_f (new_AGEMA_signal_2806), .Z1_t (new_AGEMA_signal_2807), .Z1_f (new_AGEMA_signal_2808) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_11_YY[1]), .A0_f (new_AGEMA_signal_3143), .A1_t (new_AGEMA_signal_3144), .A1_f (new_AGEMA_signal_3145), .B0_t (SubCellInst_SboxInst_11_YY_3), .B0_f (new_AGEMA_signal_3495), .B1_t (new_AGEMA_signal_3496), .B1_f (new_AGEMA_signal_3497), .Z0_t (SubCellOutput[45]), .Z0_f (new_AGEMA_signal_3669), .Z1_t (new_AGEMA_signal_3670), .Z1_f (new_AGEMA_signal_3671) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[50]), .A0_f (Ciphertext_s0_f[50]), .A1_t (Ciphertext_s1_t[50]), .A1_f (Ciphertext_s1_f[50]), .B0_t (Ciphertext_s0_t[51]), .B0_f (Ciphertext_s0_f[51]), .B1_t (Ciphertext_s1_t[51]), .B1_f (Ciphertext_s1_f[51]), .Z0_t (SubCellInst_SboxInst_12_XX[1]), .Z0_f (new_AGEMA_signal_1633), .Z1_t (new_AGEMA_signal_1634), .Z1_f (new_AGEMA_signal_1635) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[48]), .A0_f (Ciphertext_s0_f[48]), .A1_t (Ciphertext_s1_t[48]), .A1_f (Ciphertext_s1_f[48]), .B0_t (Ciphertext_s0_t[50]), .B0_f (Ciphertext_s0_f[50]), .B1_t (Ciphertext_s1_t[50]), .B1_f (Ciphertext_s1_f[50]), .Z0_t (SubCellInst_SboxInst_12_XX[2]), .Z0_f (new_AGEMA_signal_1639), .Z1_t (new_AGEMA_signal_1640), .Z1_f (new_AGEMA_signal_1641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR0_U1 ( .A0_t (Ciphertext_s0_t[49]), .A0_f (Ciphertext_s0_f[49]), .A1_t (Ciphertext_s1_t[49]), .A1_f (Ciphertext_s1_f[49]), .B0_t (SubCellInst_SboxInst_12_XX[2]), .B0_f (new_AGEMA_signal_1639), .B1_t (new_AGEMA_signal_1640), .B1_f (new_AGEMA_signal_1641), .Z0_t (SubCellInst_SboxInst_12_Q0), .Z0_f (new_AGEMA_signal_2457), .Z1_t (new_AGEMA_signal_2458), .Z1_f (new_AGEMA_signal_2459) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR1_U1 ( .A0_t (Ciphertext_s0_t[49]), .A0_f (Ciphertext_s0_f[49]), .A1_t (Ciphertext_s1_t[49]), .A1_f (Ciphertext_s1_f[49]), .B0_t (SubCellInst_SboxInst_12_XX[1]), .B0_f (new_AGEMA_signal_1633), .B1_t (new_AGEMA_signal_1634), .B1_f (new_AGEMA_signal_1635), .Z0_t (SubCellInst_SboxInst_12_Q1), .Z0_f (new_AGEMA_signal_2460), .Z1_t (new_AGEMA_signal_2461), .Z1_f (new_AGEMA_signal_2462) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_AND1_U1 ( .A0_t (Ciphertext_s0_t[50]), .A0_f (Ciphertext_s0_f[50]), .A1_t (Ciphertext_s1_t[50]), .A1_f (Ciphertext_s1_f[50]), .B0_t (SubCellInst_SboxInst_12_Q1), .B0_f (new_AGEMA_signal_2460), .B1_t (new_AGEMA_signal_2461), .B1_f (new_AGEMA_signal_2462), .Z0_t (SubCellInst_SboxInst_12_T0), .Z0_f (new_AGEMA_signal_2809), .Z1_t (new_AGEMA_signal_2810), .Z1_f (new_AGEMA_signal_2811) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_12_Q0), .A0_f (new_AGEMA_signal_2457), .A1_t (new_AGEMA_signal_2458), .A1_f (new_AGEMA_signal_2459), .B0_t (SubCellInst_SboxInst_12_T0), .B0_f (new_AGEMA_signal_2809), .B1_t (new_AGEMA_signal_2810), .B1_f (new_AGEMA_signal_2811), .Z0_t (SubCellInst_SboxInst_12_Q2), .Z0_f (new_AGEMA_signal_2957), .Z1_t (new_AGEMA_signal_2958), .Z1_f (new_AGEMA_signal_2959) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_AND2_U1 ( .A0_t (Ciphertext_s0_t[49]), .A0_f (Ciphertext_s0_f[49]), .A1_t (Ciphertext_s1_t[49]), .A1_f (Ciphertext_s1_f[49]), .B0_t (SubCellInst_SboxInst_12_Q2), .B0_f (new_AGEMA_signal_2957), .B1_t (new_AGEMA_signal_2958), .B1_f (new_AGEMA_signal_2959), .Z0_t (SubCellInst_SboxInst_12_T1), .Z0_f (new_AGEMA_signal_3146), .Z1_t (new_AGEMA_signal_3147), .Z1_f (new_AGEMA_signal_3148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_XOR3_U1 ( .A0_t (Ciphertext_s0_t[49]), .A0_f (Ciphertext_s0_f[49]), .A1_t (Ciphertext_s1_t[49]), .A1_f (Ciphertext_s1_f[49]), .B0_t (Ciphertext_s0_t[50]), .B0_f (Ciphertext_s0_f[50]), .B1_t (Ciphertext_s1_t[50]), .B1_f (Ciphertext_s1_f[50]), .Z0_t (SubCellInst_SboxInst_12_Q4), .Z0_f (new_AGEMA_signal_1645), .Z1_t (new_AGEMA_signal_1646), .Z1_f (new_AGEMA_signal_1647) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_AND3_U1 ( .A0_t (Ciphertext_s0_t[50]), .A0_f (Ciphertext_s0_f[50]), .A1_t (Ciphertext_s1_t[50]), .A1_f (Ciphertext_s1_f[50]), .B0_t (SubCellInst_SboxInst_12_Q4), .B0_f (new_AGEMA_signal_1645), .B1_t (new_AGEMA_signal_1646), .B1_f (new_AGEMA_signal_1647), .Z0_t (SubCellInst_SboxInst_12_T2), .Z0_f (new_AGEMA_signal_2463), .Z1_t (new_AGEMA_signal_2464), .Z1_f (new_AGEMA_signal_2465) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_12_T1), .A0_f (new_AGEMA_signal_3146), .A1_t (new_AGEMA_signal_3147), .A1_f (new_AGEMA_signal_3148), .B0_t (SubCellInst_SboxInst_12_T2), .B0_f (new_AGEMA_signal_2463), .B1_t (new_AGEMA_signal_2464), .B1_f (new_AGEMA_signal_2465), .Z0_t (SubCellInst_SboxInst_12_L0), .Z0_f (new_AGEMA_signal_3311), .Z1_t (new_AGEMA_signal_3312), .Z1_f (new_AGEMA_signal_3313) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_12_XX[2]), .A0_f (new_AGEMA_signal_1639), .A1_t (new_AGEMA_signal_1640), .A1_f (new_AGEMA_signal_1641), .B0_t (Ciphertext_s0_t[50]), .B0_f (Ciphertext_s0_f[50]), .B1_t (Ciphertext_s1_t[50]), .B1_f (Ciphertext_s1_f[50]), .Z0_t (SubCellInst_SboxInst_12_Q6), .Z0_f (new_AGEMA_signal_2466), .Z1_t (new_AGEMA_signal_2467), .Z1_f (new_AGEMA_signal_2468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_12_Q1), .A0_f (new_AGEMA_signal_2460), .A1_t (new_AGEMA_signal_2461), .A1_f (new_AGEMA_signal_2462), .B0_t (SubCellInst_SboxInst_12_Q6), .B0_f (new_AGEMA_signal_2466), .B1_t (new_AGEMA_signal_2467), .B1_f (new_AGEMA_signal_2468), .Z0_t (SubCellInst_SboxInst_12_L1), .Z0_f (new_AGEMA_signal_2812), .Z1_t (new_AGEMA_signal_2813), .Z1_f (new_AGEMA_signal_2814) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_12_L1), .A0_f (new_AGEMA_signal_2812), .A1_t (new_AGEMA_signal_2813), .A1_f (new_AGEMA_signal_2814), .B0_t (SubCellInst_SboxInst_12_T2), .B0_f (new_AGEMA_signal_2463), .B1_t (new_AGEMA_signal_2464), .B1_f (new_AGEMA_signal_2465), .Z0_t (SubCellInst_SboxInst_12_Q7), .Z0_f (new_AGEMA_signal_2960), .Z1_t (new_AGEMA_signal_2961), .Z1_f (new_AGEMA_signal_2962) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_AND4_U1 ( .A0_t (SubCellInst_SboxInst_12_Q6), .A0_f (new_AGEMA_signal_2466), .A1_t (new_AGEMA_signal_2467), .A1_f (new_AGEMA_signal_2468), .B0_t (SubCellInst_SboxInst_12_Q7), .B0_f (new_AGEMA_signal_2960), .B1_t (new_AGEMA_signal_2961), .B1_f (new_AGEMA_signal_2962), .Z0_t (SubCellInst_SboxInst_12_T3), .Z0_f (new_AGEMA_signal_3149), .Z1_t (new_AGEMA_signal_3150), .Z1_f (new_AGEMA_signal_3151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR8_U1 ( .A0_t (Ciphertext_s0_t[49]), .A0_f (Ciphertext_s0_f[49]), .A1_t (Ciphertext_s1_t[49]), .A1_f (Ciphertext_s1_f[49]), .B0_t (Ciphertext_s0_t[50]), .B0_f (Ciphertext_s0_f[50]), .B1_t (Ciphertext_s1_t[50]), .B1_f (Ciphertext_s1_f[50]), .Z0_t (SubCellInst_SboxInst_12_L2), .Z0_f (new_AGEMA_signal_1648), .Z1_t (new_AGEMA_signal_1649), .Z1_f (new_AGEMA_signal_1650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_12_L0), .A0_f (new_AGEMA_signal_3311), .A1_t (new_AGEMA_signal_3312), .A1_f (new_AGEMA_signal_3313), .B0_t (SubCellInst_SboxInst_12_L2), .B0_f (new_AGEMA_signal_1648), .B1_t (new_AGEMA_signal_1649), .B1_f (new_AGEMA_signal_1650), .Z0_t (SubCellInst_SboxInst_12_YY_3), .Z0_f (new_AGEMA_signal_3501), .Z1_t (new_AGEMA_signal_3502), .Z1_f (new_AGEMA_signal_3503) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_12_L0), .A0_f (new_AGEMA_signal_3311), .A1_t (new_AGEMA_signal_3312), .A1_f (new_AGEMA_signal_3313), .B0_t (SubCellInst_SboxInst_12_T3), .B0_f (new_AGEMA_signal_3149), .B1_t (new_AGEMA_signal_3150), .B1_f (new_AGEMA_signal_3151), .Z0_t (AddRoundConstantOutput[48]), .Z0_f (new_AGEMA_signal_3504), .Z1_t (new_AGEMA_signal_3505), .Z1_f (new_AGEMA_signal_3506) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_12_XX[2]), .A0_f (new_AGEMA_signal_1639), .A1_t (new_AGEMA_signal_1640), .A1_f (new_AGEMA_signal_1641), .B0_t (SubCellInst_SboxInst_12_T0), .B0_f (new_AGEMA_signal_2809), .B1_t (new_AGEMA_signal_2810), .B1_f (new_AGEMA_signal_2811), .Z0_t (SubCellInst_SboxInst_12_L3), .Z0_f (new_AGEMA_signal_2963), .Z1_t (new_AGEMA_signal_2964), .Z1_f (new_AGEMA_signal_2965) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_12_L3), .A0_f (new_AGEMA_signal_2963), .A1_t (new_AGEMA_signal_2964), .A1_f (new_AGEMA_signal_2965), .B0_t (SubCellInst_SboxInst_12_T2), .B0_f (new_AGEMA_signal_2463), .B1_t (new_AGEMA_signal_2464), .B1_f (new_AGEMA_signal_2465), .Z0_t (SubCellInst_SboxInst_12_YY[1]), .Z0_f (new_AGEMA_signal_3152), .Z1_t (new_AGEMA_signal_3153), .Z1_f (new_AGEMA_signal_3154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_12_XX[1]), .A0_f (new_AGEMA_signal_1633), .A1_t (new_AGEMA_signal_1634), .A1_f (new_AGEMA_signal_1635), .B0_t (SubCellInst_SboxInst_12_T2), .B0_f (new_AGEMA_signal_2463), .B1_t (new_AGEMA_signal_2464), .B1_f (new_AGEMA_signal_2465), .Z0_t (SubCellInst_SboxInst_12_YY[0]), .Z0_f (new_AGEMA_signal_2815), .Z1_t (new_AGEMA_signal_2816), .Z1_f (new_AGEMA_signal_2817) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_12_YY[1]), .A0_f (new_AGEMA_signal_3152), .A1_t (new_AGEMA_signal_3153), .A1_f (new_AGEMA_signal_3154), .B0_t (SubCellInst_SboxInst_12_YY_3), .B0_f (new_AGEMA_signal_3501), .B1_t (new_AGEMA_signal_3502), .B1_f (new_AGEMA_signal_3503), .Z0_t (AddRoundConstantOutput[49]), .Z0_f (new_AGEMA_signal_3672), .Z1_t (new_AGEMA_signal_3673), .Z1_f (new_AGEMA_signal_3674) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[54]), .A0_f (Ciphertext_s0_f[54]), .A1_t (Ciphertext_s1_t[54]), .A1_f (Ciphertext_s1_f[54]), .B0_t (Ciphertext_s0_t[55]), .B0_f (Ciphertext_s0_f[55]), .B1_t (Ciphertext_s1_t[55]), .B1_f (Ciphertext_s1_f[55]), .Z0_t (SubCellInst_SboxInst_13_XX[1]), .Z0_f (new_AGEMA_signal_1657), .Z1_t (new_AGEMA_signal_1658), .Z1_f (new_AGEMA_signal_1659) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[52]), .A0_f (Ciphertext_s0_f[52]), .A1_t (Ciphertext_s1_t[52]), .A1_f (Ciphertext_s1_f[52]), .B0_t (Ciphertext_s0_t[54]), .B0_f (Ciphertext_s0_f[54]), .B1_t (Ciphertext_s1_t[54]), .B1_f (Ciphertext_s1_f[54]), .Z0_t (SubCellInst_SboxInst_13_XX[2]), .Z0_f (new_AGEMA_signal_1663), .Z1_t (new_AGEMA_signal_1664), .Z1_f (new_AGEMA_signal_1665) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR0_U1 ( .A0_t (Ciphertext_s0_t[53]), .A0_f (Ciphertext_s0_f[53]), .A1_t (Ciphertext_s1_t[53]), .A1_f (Ciphertext_s1_f[53]), .B0_t (SubCellInst_SboxInst_13_XX[2]), .B0_f (new_AGEMA_signal_1663), .B1_t (new_AGEMA_signal_1664), .B1_f (new_AGEMA_signal_1665), .Z0_t (SubCellInst_SboxInst_13_Q0), .Z0_f (new_AGEMA_signal_2469), .Z1_t (new_AGEMA_signal_2470), .Z1_f (new_AGEMA_signal_2471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR1_U1 ( .A0_t (Ciphertext_s0_t[53]), .A0_f (Ciphertext_s0_f[53]), .A1_t (Ciphertext_s1_t[53]), .A1_f (Ciphertext_s1_f[53]), .B0_t (SubCellInst_SboxInst_13_XX[1]), .B0_f (new_AGEMA_signal_1657), .B1_t (new_AGEMA_signal_1658), .B1_f (new_AGEMA_signal_1659), .Z0_t (SubCellInst_SboxInst_13_Q1), .Z0_f (new_AGEMA_signal_2472), .Z1_t (new_AGEMA_signal_2473), .Z1_f (new_AGEMA_signal_2474) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_AND1_U1 ( .A0_t (Ciphertext_s0_t[54]), .A0_f (Ciphertext_s0_f[54]), .A1_t (Ciphertext_s1_t[54]), .A1_f (Ciphertext_s1_f[54]), .B0_t (SubCellInst_SboxInst_13_Q1), .B0_f (new_AGEMA_signal_2472), .B1_t (new_AGEMA_signal_2473), .B1_f (new_AGEMA_signal_2474), .Z0_t (SubCellInst_SboxInst_13_T0), .Z0_f (new_AGEMA_signal_2818), .Z1_t (new_AGEMA_signal_2819), .Z1_f (new_AGEMA_signal_2820) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_13_Q0), .A0_f (new_AGEMA_signal_2469), .A1_t (new_AGEMA_signal_2470), .A1_f (new_AGEMA_signal_2471), .B0_t (SubCellInst_SboxInst_13_T0), .B0_f (new_AGEMA_signal_2818), .B1_t (new_AGEMA_signal_2819), .B1_f (new_AGEMA_signal_2820), .Z0_t (SubCellInst_SboxInst_13_Q2), .Z0_f (new_AGEMA_signal_2966), .Z1_t (new_AGEMA_signal_2967), .Z1_f (new_AGEMA_signal_2968) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_AND2_U1 ( .A0_t (Ciphertext_s0_t[53]), .A0_f (Ciphertext_s0_f[53]), .A1_t (Ciphertext_s1_t[53]), .A1_f (Ciphertext_s1_f[53]), .B0_t (SubCellInst_SboxInst_13_Q2), .B0_f (new_AGEMA_signal_2966), .B1_t (new_AGEMA_signal_2967), .B1_f (new_AGEMA_signal_2968), .Z0_t (SubCellInst_SboxInst_13_T1), .Z0_f (new_AGEMA_signal_3155), .Z1_t (new_AGEMA_signal_3156), .Z1_f (new_AGEMA_signal_3157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_XOR3_U1 ( .A0_t (Ciphertext_s0_t[53]), .A0_f (Ciphertext_s0_f[53]), .A1_t (Ciphertext_s1_t[53]), .A1_f (Ciphertext_s1_f[53]), .B0_t (Ciphertext_s0_t[54]), .B0_f (Ciphertext_s0_f[54]), .B1_t (Ciphertext_s1_t[54]), .B1_f (Ciphertext_s1_f[54]), .Z0_t (SubCellInst_SboxInst_13_Q4), .Z0_f (new_AGEMA_signal_1669), .Z1_t (new_AGEMA_signal_1670), .Z1_f (new_AGEMA_signal_1671) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_AND3_U1 ( .A0_t (Ciphertext_s0_t[54]), .A0_f (Ciphertext_s0_f[54]), .A1_t (Ciphertext_s1_t[54]), .A1_f (Ciphertext_s1_f[54]), .B0_t (SubCellInst_SboxInst_13_Q4), .B0_f (new_AGEMA_signal_1669), .B1_t (new_AGEMA_signal_1670), .B1_f (new_AGEMA_signal_1671), .Z0_t (SubCellInst_SboxInst_13_T2), .Z0_f (new_AGEMA_signal_2475), .Z1_t (new_AGEMA_signal_2476), .Z1_f (new_AGEMA_signal_2477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_13_T1), .A0_f (new_AGEMA_signal_3155), .A1_t (new_AGEMA_signal_3156), .A1_f (new_AGEMA_signal_3157), .B0_t (SubCellInst_SboxInst_13_T2), .B0_f (new_AGEMA_signal_2475), .B1_t (new_AGEMA_signal_2476), .B1_f (new_AGEMA_signal_2477), .Z0_t (SubCellInst_SboxInst_13_L0), .Z0_f (new_AGEMA_signal_3314), .Z1_t (new_AGEMA_signal_3315), .Z1_f (new_AGEMA_signal_3316) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_13_XX[2]), .A0_f (new_AGEMA_signal_1663), .A1_t (new_AGEMA_signal_1664), .A1_f (new_AGEMA_signal_1665), .B0_t (Ciphertext_s0_t[54]), .B0_f (Ciphertext_s0_f[54]), .B1_t (Ciphertext_s1_t[54]), .B1_f (Ciphertext_s1_f[54]), .Z0_t (SubCellInst_SboxInst_13_Q6), .Z0_f (new_AGEMA_signal_2478), .Z1_t (new_AGEMA_signal_2479), .Z1_f (new_AGEMA_signal_2480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_13_Q1), .A0_f (new_AGEMA_signal_2472), .A1_t (new_AGEMA_signal_2473), .A1_f (new_AGEMA_signal_2474), .B0_t (SubCellInst_SboxInst_13_Q6), .B0_f (new_AGEMA_signal_2478), .B1_t (new_AGEMA_signal_2479), .B1_f (new_AGEMA_signal_2480), .Z0_t (SubCellInst_SboxInst_13_L1), .Z0_f (new_AGEMA_signal_2821), .Z1_t (new_AGEMA_signal_2822), .Z1_f (new_AGEMA_signal_2823) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_13_L1), .A0_f (new_AGEMA_signal_2821), .A1_t (new_AGEMA_signal_2822), .A1_f (new_AGEMA_signal_2823), .B0_t (SubCellInst_SboxInst_13_T2), .B0_f (new_AGEMA_signal_2475), .B1_t (new_AGEMA_signal_2476), .B1_f (new_AGEMA_signal_2477), .Z0_t (SubCellInst_SboxInst_13_Q7), .Z0_f (new_AGEMA_signal_2969), .Z1_t (new_AGEMA_signal_2970), .Z1_f (new_AGEMA_signal_2971) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_AND4_U1 ( .A0_t (SubCellInst_SboxInst_13_Q6), .A0_f (new_AGEMA_signal_2478), .A1_t (new_AGEMA_signal_2479), .A1_f (new_AGEMA_signal_2480), .B0_t (SubCellInst_SboxInst_13_Q7), .B0_f (new_AGEMA_signal_2969), .B1_t (new_AGEMA_signal_2970), .B1_f (new_AGEMA_signal_2971), .Z0_t (SubCellInst_SboxInst_13_T3), .Z0_f (new_AGEMA_signal_3158), .Z1_t (new_AGEMA_signal_3159), .Z1_f (new_AGEMA_signal_3160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR8_U1 ( .A0_t (Ciphertext_s0_t[53]), .A0_f (Ciphertext_s0_f[53]), .A1_t (Ciphertext_s1_t[53]), .A1_f (Ciphertext_s1_f[53]), .B0_t (Ciphertext_s0_t[54]), .B0_f (Ciphertext_s0_f[54]), .B1_t (Ciphertext_s1_t[54]), .B1_f (Ciphertext_s1_f[54]), .Z0_t (SubCellInst_SboxInst_13_L2), .Z0_f (new_AGEMA_signal_1672), .Z1_t (new_AGEMA_signal_1673), .Z1_f (new_AGEMA_signal_1674) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_13_L0), .A0_f (new_AGEMA_signal_3314), .A1_t (new_AGEMA_signal_3315), .A1_f (new_AGEMA_signal_3316), .B0_t (SubCellInst_SboxInst_13_L2), .B0_f (new_AGEMA_signal_1672), .B1_t (new_AGEMA_signal_1673), .B1_f (new_AGEMA_signal_1674), .Z0_t (SubCellInst_SboxInst_13_YY_3), .Z0_f (new_AGEMA_signal_3507), .Z1_t (new_AGEMA_signal_3508), .Z1_f (new_AGEMA_signal_3509) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_13_L0), .A0_f (new_AGEMA_signal_3314), .A1_t (new_AGEMA_signal_3315), .A1_f (new_AGEMA_signal_3316), .B0_t (SubCellInst_SboxInst_13_T3), .B0_f (new_AGEMA_signal_3158), .B1_t (new_AGEMA_signal_3159), .B1_f (new_AGEMA_signal_3160), .Z0_t (AddRoundConstantOutput[52]), .Z0_f (new_AGEMA_signal_3510), .Z1_t (new_AGEMA_signal_3511), .Z1_f (new_AGEMA_signal_3512) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_13_XX[2]), .A0_f (new_AGEMA_signal_1663), .A1_t (new_AGEMA_signal_1664), .A1_f (new_AGEMA_signal_1665), .B0_t (SubCellInst_SboxInst_13_T0), .B0_f (new_AGEMA_signal_2818), .B1_t (new_AGEMA_signal_2819), .B1_f (new_AGEMA_signal_2820), .Z0_t (SubCellInst_SboxInst_13_L3), .Z0_f (new_AGEMA_signal_2972), .Z1_t (new_AGEMA_signal_2973), .Z1_f (new_AGEMA_signal_2974) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_13_L3), .A0_f (new_AGEMA_signal_2972), .A1_t (new_AGEMA_signal_2973), .A1_f (new_AGEMA_signal_2974), .B0_t (SubCellInst_SboxInst_13_T2), .B0_f (new_AGEMA_signal_2475), .B1_t (new_AGEMA_signal_2476), .B1_f (new_AGEMA_signal_2477), .Z0_t (SubCellInst_SboxInst_13_YY[1]), .Z0_f (new_AGEMA_signal_3161), .Z1_t (new_AGEMA_signal_3162), .Z1_f (new_AGEMA_signal_3163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_13_XX[1]), .A0_f (new_AGEMA_signal_1657), .A1_t (new_AGEMA_signal_1658), .A1_f (new_AGEMA_signal_1659), .B0_t (SubCellInst_SboxInst_13_T2), .B0_f (new_AGEMA_signal_2475), .B1_t (new_AGEMA_signal_2476), .B1_f (new_AGEMA_signal_2477), .Z0_t (SubCellInst_SboxInst_13_YY[0]), .Z0_f (new_AGEMA_signal_2824), .Z1_t (new_AGEMA_signal_2825), .Z1_f (new_AGEMA_signal_2826) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_13_YY[1]), .A0_f (new_AGEMA_signal_3161), .A1_t (new_AGEMA_signal_3162), .A1_f (new_AGEMA_signal_3163), .B0_t (SubCellInst_SboxInst_13_YY_3), .B0_f (new_AGEMA_signal_3507), .B1_t (new_AGEMA_signal_3508), .B1_f (new_AGEMA_signal_3509), .Z0_t (AddRoundConstantOutput[53]), .Z0_f (new_AGEMA_signal_3675), .Z1_t (new_AGEMA_signal_3676), .Z1_f (new_AGEMA_signal_3677) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[58]), .A0_f (Ciphertext_s0_f[58]), .A1_t (Ciphertext_s1_t[58]), .A1_f (Ciphertext_s1_f[58]), .B0_t (Ciphertext_s0_t[59]), .B0_f (Ciphertext_s0_f[59]), .B1_t (Ciphertext_s1_t[59]), .B1_f (Ciphertext_s1_f[59]), .Z0_t (SubCellInst_SboxInst_14_XX[1]), .Z0_f (new_AGEMA_signal_1681), .Z1_t (new_AGEMA_signal_1682), .Z1_f (new_AGEMA_signal_1683) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[56]), .A0_f (Ciphertext_s0_f[56]), .A1_t (Ciphertext_s1_t[56]), .A1_f (Ciphertext_s1_f[56]), .B0_t (Ciphertext_s0_t[58]), .B0_f (Ciphertext_s0_f[58]), .B1_t (Ciphertext_s1_t[58]), .B1_f (Ciphertext_s1_f[58]), .Z0_t (SubCellInst_SboxInst_14_XX[2]), .Z0_f (new_AGEMA_signal_1687), .Z1_t (new_AGEMA_signal_1688), .Z1_f (new_AGEMA_signal_1689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR0_U1 ( .A0_t (Ciphertext_s0_t[57]), .A0_f (Ciphertext_s0_f[57]), .A1_t (Ciphertext_s1_t[57]), .A1_f (Ciphertext_s1_f[57]), .B0_t (SubCellInst_SboxInst_14_XX[2]), .B0_f (new_AGEMA_signal_1687), .B1_t (new_AGEMA_signal_1688), .B1_f (new_AGEMA_signal_1689), .Z0_t (SubCellInst_SboxInst_14_Q0), .Z0_f (new_AGEMA_signal_2481), .Z1_t (new_AGEMA_signal_2482), .Z1_f (new_AGEMA_signal_2483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR1_U1 ( .A0_t (Ciphertext_s0_t[57]), .A0_f (Ciphertext_s0_f[57]), .A1_t (Ciphertext_s1_t[57]), .A1_f (Ciphertext_s1_f[57]), .B0_t (SubCellInst_SboxInst_14_XX[1]), .B0_f (new_AGEMA_signal_1681), .B1_t (new_AGEMA_signal_1682), .B1_f (new_AGEMA_signal_1683), .Z0_t (SubCellInst_SboxInst_14_Q1), .Z0_f (new_AGEMA_signal_2484), .Z1_t (new_AGEMA_signal_2485), .Z1_f (new_AGEMA_signal_2486) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_AND1_U1 ( .A0_t (Ciphertext_s0_t[58]), .A0_f (Ciphertext_s0_f[58]), .A1_t (Ciphertext_s1_t[58]), .A1_f (Ciphertext_s1_f[58]), .B0_t (SubCellInst_SboxInst_14_Q1), .B0_f (new_AGEMA_signal_2484), .B1_t (new_AGEMA_signal_2485), .B1_f (new_AGEMA_signal_2486), .Z0_t (SubCellInst_SboxInst_14_T0), .Z0_f (new_AGEMA_signal_2827), .Z1_t (new_AGEMA_signal_2828), .Z1_f (new_AGEMA_signal_2829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_14_Q0), .A0_f (new_AGEMA_signal_2481), .A1_t (new_AGEMA_signal_2482), .A1_f (new_AGEMA_signal_2483), .B0_t (SubCellInst_SboxInst_14_T0), .B0_f (new_AGEMA_signal_2827), .B1_t (new_AGEMA_signal_2828), .B1_f (new_AGEMA_signal_2829), .Z0_t (SubCellInst_SboxInst_14_Q2), .Z0_f (new_AGEMA_signal_2975), .Z1_t (new_AGEMA_signal_2976), .Z1_f (new_AGEMA_signal_2977) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_AND2_U1 ( .A0_t (Ciphertext_s0_t[57]), .A0_f (Ciphertext_s0_f[57]), .A1_t (Ciphertext_s1_t[57]), .A1_f (Ciphertext_s1_f[57]), .B0_t (SubCellInst_SboxInst_14_Q2), .B0_f (new_AGEMA_signal_2975), .B1_t (new_AGEMA_signal_2976), .B1_f (new_AGEMA_signal_2977), .Z0_t (SubCellInst_SboxInst_14_T1), .Z0_f (new_AGEMA_signal_3164), .Z1_t (new_AGEMA_signal_3165), .Z1_f (new_AGEMA_signal_3166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_XOR3_U1 ( .A0_t (Ciphertext_s0_t[57]), .A0_f (Ciphertext_s0_f[57]), .A1_t (Ciphertext_s1_t[57]), .A1_f (Ciphertext_s1_f[57]), .B0_t (Ciphertext_s0_t[58]), .B0_f (Ciphertext_s0_f[58]), .B1_t (Ciphertext_s1_t[58]), .B1_f (Ciphertext_s1_f[58]), .Z0_t (SubCellInst_SboxInst_14_Q4), .Z0_f (new_AGEMA_signal_1693), .Z1_t (new_AGEMA_signal_1694), .Z1_f (new_AGEMA_signal_1695) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_AND3_U1 ( .A0_t (Ciphertext_s0_t[58]), .A0_f (Ciphertext_s0_f[58]), .A1_t (Ciphertext_s1_t[58]), .A1_f (Ciphertext_s1_f[58]), .B0_t (SubCellInst_SboxInst_14_Q4), .B0_f (new_AGEMA_signal_1693), .B1_t (new_AGEMA_signal_1694), .B1_f (new_AGEMA_signal_1695), .Z0_t (SubCellInst_SboxInst_14_T2), .Z0_f (new_AGEMA_signal_2487), .Z1_t (new_AGEMA_signal_2488), .Z1_f (new_AGEMA_signal_2489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_14_T1), .A0_f (new_AGEMA_signal_3164), .A1_t (new_AGEMA_signal_3165), .A1_f (new_AGEMA_signal_3166), .B0_t (SubCellInst_SboxInst_14_T2), .B0_f (new_AGEMA_signal_2487), .B1_t (new_AGEMA_signal_2488), .B1_f (new_AGEMA_signal_2489), .Z0_t (SubCellInst_SboxInst_14_L0), .Z0_f (new_AGEMA_signal_3317), .Z1_t (new_AGEMA_signal_3318), .Z1_f (new_AGEMA_signal_3319) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_14_XX[2]), .A0_f (new_AGEMA_signal_1687), .A1_t (new_AGEMA_signal_1688), .A1_f (new_AGEMA_signal_1689), .B0_t (Ciphertext_s0_t[58]), .B0_f (Ciphertext_s0_f[58]), .B1_t (Ciphertext_s1_t[58]), .B1_f (Ciphertext_s1_f[58]), .Z0_t (SubCellInst_SboxInst_14_Q6), .Z0_f (new_AGEMA_signal_2490), .Z1_t (new_AGEMA_signal_2491), .Z1_f (new_AGEMA_signal_2492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_14_Q1), .A0_f (new_AGEMA_signal_2484), .A1_t (new_AGEMA_signal_2485), .A1_f (new_AGEMA_signal_2486), .B0_t (SubCellInst_SboxInst_14_Q6), .B0_f (new_AGEMA_signal_2490), .B1_t (new_AGEMA_signal_2491), .B1_f (new_AGEMA_signal_2492), .Z0_t (SubCellInst_SboxInst_14_L1), .Z0_f (new_AGEMA_signal_2830), .Z1_t (new_AGEMA_signal_2831), .Z1_f (new_AGEMA_signal_2832) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_14_L1), .A0_f (new_AGEMA_signal_2830), .A1_t (new_AGEMA_signal_2831), .A1_f (new_AGEMA_signal_2832), .B0_t (SubCellInst_SboxInst_14_T2), .B0_f (new_AGEMA_signal_2487), .B1_t (new_AGEMA_signal_2488), .B1_f (new_AGEMA_signal_2489), .Z0_t (SubCellInst_SboxInst_14_Q7), .Z0_f (new_AGEMA_signal_2978), .Z1_t (new_AGEMA_signal_2979), .Z1_f (new_AGEMA_signal_2980) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_AND4_U1 ( .A0_t (SubCellInst_SboxInst_14_Q6), .A0_f (new_AGEMA_signal_2490), .A1_t (new_AGEMA_signal_2491), .A1_f (new_AGEMA_signal_2492), .B0_t (SubCellInst_SboxInst_14_Q7), .B0_f (new_AGEMA_signal_2978), .B1_t (new_AGEMA_signal_2979), .B1_f (new_AGEMA_signal_2980), .Z0_t (SubCellInst_SboxInst_14_T3), .Z0_f (new_AGEMA_signal_3167), .Z1_t (new_AGEMA_signal_3168), .Z1_f (new_AGEMA_signal_3169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR8_U1 ( .A0_t (Ciphertext_s0_t[57]), .A0_f (Ciphertext_s0_f[57]), .A1_t (Ciphertext_s1_t[57]), .A1_f (Ciphertext_s1_f[57]), .B0_t (Ciphertext_s0_t[58]), .B0_f (Ciphertext_s0_f[58]), .B1_t (Ciphertext_s1_t[58]), .B1_f (Ciphertext_s1_f[58]), .Z0_t (SubCellInst_SboxInst_14_L2), .Z0_f (new_AGEMA_signal_1696), .Z1_t (new_AGEMA_signal_1697), .Z1_f (new_AGEMA_signal_1698) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_14_L0), .A0_f (new_AGEMA_signal_3317), .A1_t (new_AGEMA_signal_3318), .A1_f (new_AGEMA_signal_3319), .B0_t (SubCellInst_SboxInst_14_L2), .B0_f (new_AGEMA_signal_1696), .B1_t (new_AGEMA_signal_1697), .B1_f (new_AGEMA_signal_1698), .Z0_t (SubCellInst_SboxInst_14_YY_3), .Z0_f (new_AGEMA_signal_3513), .Z1_t (new_AGEMA_signal_3514), .Z1_f (new_AGEMA_signal_3515) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_14_L0), .A0_f (new_AGEMA_signal_3317), .A1_t (new_AGEMA_signal_3318), .A1_f (new_AGEMA_signal_3319), .B0_t (SubCellInst_SboxInst_14_T3), .B0_f (new_AGEMA_signal_3167), .B1_t (new_AGEMA_signal_3168), .B1_f (new_AGEMA_signal_3169), .Z0_t (AddRoundConstantOutput[56]), .Z0_f (new_AGEMA_signal_3516), .Z1_t (new_AGEMA_signal_3517), .Z1_f (new_AGEMA_signal_3518) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_14_XX[2]), .A0_f (new_AGEMA_signal_1687), .A1_t (new_AGEMA_signal_1688), .A1_f (new_AGEMA_signal_1689), .B0_t (SubCellInst_SboxInst_14_T0), .B0_f (new_AGEMA_signal_2827), .B1_t (new_AGEMA_signal_2828), .B1_f (new_AGEMA_signal_2829), .Z0_t (SubCellInst_SboxInst_14_L3), .Z0_f (new_AGEMA_signal_2981), .Z1_t (new_AGEMA_signal_2982), .Z1_f (new_AGEMA_signal_2983) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_14_L3), .A0_f (new_AGEMA_signal_2981), .A1_t (new_AGEMA_signal_2982), .A1_f (new_AGEMA_signal_2983), .B0_t (SubCellInst_SboxInst_14_T2), .B0_f (new_AGEMA_signal_2487), .B1_t (new_AGEMA_signal_2488), .B1_f (new_AGEMA_signal_2489), .Z0_t (SubCellInst_SboxInst_14_YY[1]), .Z0_f (new_AGEMA_signal_3170), .Z1_t (new_AGEMA_signal_3171), .Z1_f (new_AGEMA_signal_3172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_14_XX[1]), .A0_f (new_AGEMA_signal_1681), .A1_t (new_AGEMA_signal_1682), .A1_f (new_AGEMA_signal_1683), .B0_t (SubCellInst_SboxInst_14_T2), .B0_f (new_AGEMA_signal_2487), .B1_t (new_AGEMA_signal_2488), .B1_f (new_AGEMA_signal_2489), .Z0_t (SubCellInst_SboxInst_14_YY[0]), .Z0_f (new_AGEMA_signal_2833), .Z1_t (new_AGEMA_signal_2834), .Z1_f (new_AGEMA_signal_2835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_14_YY[1]), .A0_f (new_AGEMA_signal_3170), .A1_t (new_AGEMA_signal_3171), .A1_f (new_AGEMA_signal_3172), .B0_t (SubCellInst_SboxInst_14_YY_3), .B0_f (new_AGEMA_signal_3513), .B1_t (new_AGEMA_signal_3514), .B1_f (new_AGEMA_signal_3515), .Z0_t (AddRoundConstantOutput[57]), .Z0_f (new_AGEMA_signal_3678), .Z1_t (new_AGEMA_signal_3679), .Z1_f (new_AGEMA_signal_3680) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR_i1_U1 ( .A0_t (Ciphertext_s0_t[62]), .A0_f (Ciphertext_s0_f[62]), .A1_t (Ciphertext_s1_t[62]), .A1_f (Ciphertext_s1_f[62]), .B0_t (Ciphertext_s0_t[63]), .B0_f (Ciphertext_s0_f[63]), .B1_t (Ciphertext_s1_t[63]), .B1_f (Ciphertext_s1_f[63]), .Z0_t (SubCellInst_SboxInst_15_XX[1]), .Z0_f (new_AGEMA_signal_1705), .Z1_t (new_AGEMA_signal_1706), .Z1_f (new_AGEMA_signal_1707) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR_i2_U1 ( .A0_t (Ciphertext_s0_t[60]), .A0_f (Ciphertext_s0_f[60]), .A1_t (Ciphertext_s1_t[60]), .A1_f (Ciphertext_s1_f[60]), .B0_t (Ciphertext_s0_t[62]), .B0_f (Ciphertext_s0_f[62]), .B1_t (Ciphertext_s1_t[62]), .B1_f (Ciphertext_s1_f[62]), .Z0_t (SubCellInst_SboxInst_15_XX[2]), .Z0_f (new_AGEMA_signal_1711), .Z1_t (new_AGEMA_signal_1712), .Z1_f (new_AGEMA_signal_1713) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR0_U1 ( .A0_t (Ciphertext_s0_t[61]), .A0_f (Ciphertext_s0_f[61]), .A1_t (Ciphertext_s1_t[61]), .A1_f (Ciphertext_s1_f[61]), .B0_t (SubCellInst_SboxInst_15_XX[2]), .B0_f (new_AGEMA_signal_1711), .B1_t (new_AGEMA_signal_1712), .B1_f (new_AGEMA_signal_1713), .Z0_t (SubCellInst_SboxInst_15_Q0), .Z0_f (new_AGEMA_signal_2493), .Z1_t (new_AGEMA_signal_2494), .Z1_f (new_AGEMA_signal_2495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR1_U1 ( .A0_t (Ciphertext_s0_t[61]), .A0_f (Ciphertext_s0_f[61]), .A1_t (Ciphertext_s1_t[61]), .A1_f (Ciphertext_s1_f[61]), .B0_t (SubCellInst_SboxInst_15_XX[1]), .B0_f (new_AGEMA_signal_1705), .B1_t (new_AGEMA_signal_1706), .B1_f (new_AGEMA_signal_1707), .Z0_t (SubCellInst_SboxInst_15_Q1), .Z0_f (new_AGEMA_signal_2496), .Z1_t (new_AGEMA_signal_2497), .Z1_f (new_AGEMA_signal_2498) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_AND1_U1 ( .A0_t (Ciphertext_s0_t[62]), .A0_f (Ciphertext_s0_f[62]), .A1_t (Ciphertext_s1_t[62]), .A1_f (Ciphertext_s1_f[62]), .B0_t (SubCellInst_SboxInst_15_Q1), .B0_f (new_AGEMA_signal_2496), .B1_t (new_AGEMA_signal_2497), .B1_f (new_AGEMA_signal_2498), .Z0_t (SubCellInst_SboxInst_15_T0), .Z0_f (new_AGEMA_signal_2836), .Z1_t (new_AGEMA_signal_2837), .Z1_f (new_AGEMA_signal_2838) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_15_Q0), .A0_f (new_AGEMA_signal_2493), .A1_t (new_AGEMA_signal_2494), .A1_f (new_AGEMA_signal_2495), .B0_t (SubCellInst_SboxInst_15_T0), .B0_f (new_AGEMA_signal_2836), .B1_t (new_AGEMA_signal_2837), .B1_f (new_AGEMA_signal_2838), .Z0_t (SubCellInst_SboxInst_15_Q2), .Z0_f (new_AGEMA_signal_2984), .Z1_t (new_AGEMA_signal_2985), .Z1_f (new_AGEMA_signal_2986) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_AND2_U1 ( .A0_t (Ciphertext_s0_t[61]), .A0_f (Ciphertext_s0_f[61]), .A1_t (Ciphertext_s1_t[61]), .A1_f (Ciphertext_s1_f[61]), .B0_t (SubCellInst_SboxInst_15_Q2), .B0_f (new_AGEMA_signal_2984), .B1_t (new_AGEMA_signal_2985), .B1_f (new_AGEMA_signal_2986), .Z0_t (SubCellInst_SboxInst_15_T1), .Z0_f (new_AGEMA_signal_3173), .Z1_t (new_AGEMA_signal_3174), .Z1_f (new_AGEMA_signal_3175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_XOR3_U1 ( .A0_t (Ciphertext_s0_t[61]), .A0_f (Ciphertext_s0_f[61]), .A1_t (Ciphertext_s1_t[61]), .A1_f (Ciphertext_s1_f[61]), .B0_t (Ciphertext_s0_t[62]), .B0_f (Ciphertext_s0_f[62]), .B1_t (Ciphertext_s1_t[62]), .B1_f (Ciphertext_s1_f[62]), .Z0_t (SubCellInst_SboxInst_15_Q4), .Z0_f (new_AGEMA_signal_1717), .Z1_t (new_AGEMA_signal_1718), .Z1_f (new_AGEMA_signal_1719) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_AND3_U1 ( .A0_t (Ciphertext_s0_t[62]), .A0_f (Ciphertext_s0_f[62]), .A1_t (Ciphertext_s1_t[62]), .A1_f (Ciphertext_s1_f[62]), .B0_t (SubCellInst_SboxInst_15_Q4), .B0_f (new_AGEMA_signal_1717), .B1_t (new_AGEMA_signal_1718), .B1_f (new_AGEMA_signal_1719), .Z0_t (SubCellInst_SboxInst_15_T2), .Z0_f (new_AGEMA_signal_2499), .Z1_t (new_AGEMA_signal_2500), .Z1_f (new_AGEMA_signal_2501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_15_T1), .A0_f (new_AGEMA_signal_3173), .A1_t (new_AGEMA_signal_3174), .A1_f (new_AGEMA_signal_3175), .B0_t (SubCellInst_SboxInst_15_T2), .B0_f (new_AGEMA_signal_2499), .B1_t (new_AGEMA_signal_2500), .B1_f (new_AGEMA_signal_2501), .Z0_t (SubCellInst_SboxInst_15_L0), .Z0_f (new_AGEMA_signal_3320), .Z1_t (new_AGEMA_signal_3321), .Z1_f (new_AGEMA_signal_3322) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_15_XX[2]), .A0_f (new_AGEMA_signal_1711), .A1_t (new_AGEMA_signal_1712), .A1_f (new_AGEMA_signal_1713), .B0_t (Ciphertext_s0_t[62]), .B0_f (Ciphertext_s0_f[62]), .B1_t (Ciphertext_s1_t[62]), .B1_f (Ciphertext_s1_f[62]), .Z0_t (SubCellInst_SboxInst_15_Q6), .Z0_f (new_AGEMA_signal_2502), .Z1_t (new_AGEMA_signal_2503), .Z1_f (new_AGEMA_signal_2504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_15_Q1), .A0_f (new_AGEMA_signal_2496), .A1_t (new_AGEMA_signal_2497), .A1_f (new_AGEMA_signal_2498), .B0_t (SubCellInst_SboxInst_15_Q6), .B0_f (new_AGEMA_signal_2502), .B1_t (new_AGEMA_signal_2503), .B1_f (new_AGEMA_signal_2504), .Z0_t (SubCellInst_SboxInst_15_L1), .Z0_f (new_AGEMA_signal_2839), .Z1_t (new_AGEMA_signal_2840), .Z1_f (new_AGEMA_signal_2841) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_15_L1), .A0_f (new_AGEMA_signal_2839), .A1_t (new_AGEMA_signal_2840), .A1_f (new_AGEMA_signal_2841), .B0_t (SubCellInst_SboxInst_15_T2), .B0_f (new_AGEMA_signal_2499), .B1_t (new_AGEMA_signal_2500), .B1_f (new_AGEMA_signal_2501), .Z0_t (SubCellInst_SboxInst_15_Q7), .Z0_f (new_AGEMA_signal_2987), .Z1_t (new_AGEMA_signal_2988), .Z1_f (new_AGEMA_signal_2989) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_AND4_U1 ( .A0_t (SubCellInst_SboxInst_15_Q6), .A0_f (new_AGEMA_signal_2502), .A1_t (new_AGEMA_signal_2503), .A1_f (new_AGEMA_signal_2504), .B0_t (SubCellInst_SboxInst_15_Q7), .B0_f (new_AGEMA_signal_2987), .B1_t (new_AGEMA_signal_2988), .B1_f (new_AGEMA_signal_2989), .Z0_t (SubCellInst_SboxInst_15_T3), .Z0_f (new_AGEMA_signal_3176), .Z1_t (new_AGEMA_signal_3177), .Z1_f (new_AGEMA_signal_3178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR8_U1 ( .A0_t (Ciphertext_s0_t[61]), .A0_f (Ciphertext_s0_f[61]), .A1_t (Ciphertext_s1_t[61]), .A1_f (Ciphertext_s1_f[61]), .B0_t (Ciphertext_s0_t[62]), .B0_f (Ciphertext_s0_f[62]), .B1_t (Ciphertext_s1_t[62]), .B1_f (Ciphertext_s1_f[62]), .Z0_t (SubCellInst_SboxInst_15_L2), .Z0_f (new_AGEMA_signal_1720), .Z1_t (new_AGEMA_signal_1721), .Z1_f (new_AGEMA_signal_1722) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_15_L0), .A0_f (new_AGEMA_signal_3320), .A1_t (new_AGEMA_signal_3321), .A1_f (new_AGEMA_signal_3322), .B0_t (SubCellInst_SboxInst_15_L2), .B0_f (new_AGEMA_signal_1720), .B1_t (new_AGEMA_signal_1721), .B1_f (new_AGEMA_signal_1722), .Z0_t (SubCellInst_SboxInst_15_YY_3), .Z0_f (new_AGEMA_signal_3519), .Z1_t (new_AGEMA_signal_3520), .Z1_f (new_AGEMA_signal_3521) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_15_L0), .A0_f (new_AGEMA_signal_3320), .A1_t (new_AGEMA_signal_3321), .A1_f (new_AGEMA_signal_3322), .B0_t (SubCellInst_SboxInst_15_T3), .B0_f (new_AGEMA_signal_3176), .B1_t (new_AGEMA_signal_3177), .B1_f (new_AGEMA_signal_3178), .Z0_t (SubCellOutput[60]), .Z0_f (new_AGEMA_signal_3522), .Z1_t (new_AGEMA_signal_3523), .Z1_f (new_AGEMA_signal_3524) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_15_XX[2]), .A0_f (new_AGEMA_signal_1711), .A1_t (new_AGEMA_signal_1712), .A1_f (new_AGEMA_signal_1713), .B0_t (SubCellInst_SboxInst_15_T0), .B0_f (new_AGEMA_signal_2836), .B1_t (new_AGEMA_signal_2837), .B1_f (new_AGEMA_signal_2838), .Z0_t (SubCellInst_SboxInst_15_L3), .Z0_f (new_AGEMA_signal_2990), .Z1_t (new_AGEMA_signal_2991), .Z1_f (new_AGEMA_signal_2992) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_15_L3), .A0_f (new_AGEMA_signal_2990), .A1_t (new_AGEMA_signal_2991), .A1_f (new_AGEMA_signal_2992), .B0_t (SubCellInst_SboxInst_15_T2), .B0_f (new_AGEMA_signal_2499), .B1_t (new_AGEMA_signal_2500), .B1_f (new_AGEMA_signal_2501), .Z0_t (SubCellInst_SboxInst_15_YY[1]), .Z0_f (new_AGEMA_signal_3179), .Z1_t (new_AGEMA_signal_3180), .Z1_f (new_AGEMA_signal_3181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_15_XX[1]), .A0_f (new_AGEMA_signal_1705), .A1_t (new_AGEMA_signal_1706), .A1_f (new_AGEMA_signal_1707), .B0_t (SubCellInst_SboxInst_15_T2), .B0_f (new_AGEMA_signal_2499), .B1_t (new_AGEMA_signal_2500), .B1_f (new_AGEMA_signal_2501), .Z0_t (SubCellInst_SboxInst_15_YY[0]), .Z0_f (new_AGEMA_signal_2842), .Z1_t (new_AGEMA_signal_2843), .Z1_f (new_AGEMA_signal_2844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_15_YY[1]), .A0_f (new_AGEMA_signal_3179), .A1_t (new_AGEMA_signal_3180), .A1_f (new_AGEMA_signal_3181), .B0_t (SubCellInst_SboxInst_15_YY_3), .B0_f (new_AGEMA_signal_3519), .B1_t (new_AGEMA_signal_3520), .B1_f (new_AGEMA_signal_3521), .Z0_t (SubCellOutput[61]), .Z0_f (new_AGEMA_signal_3681), .Z1_t (new_AGEMA_signal_3682), .Z1_f (new_AGEMA_signal_3683) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_0_0_U1 ( .A0_t (SubCellOutput[60]), .A0_f (new_AGEMA_signal_3522), .A1_t (new_AGEMA_signal_3523), .A1_f (new_AGEMA_signal_3524), .B0_t (1'b0), .B0_f (1'b1), .B1_t (FSMUpdate[1]), .B1_f (new_AGEMA_signal_2300), .Z0_t (AddRoundConstantOutput[60]), .Z0_f (new_AGEMA_signal_3684), .Z1_t (new_AGEMA_signal_3685), .Z1_f (new_AGEMA_signal_3686) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_0_1_U1 ( .A0_t (SubCellOutput[61]), .A0_f (new_AGEMA_signal_3681), .A1_t (new_AGEMA_signal_3682), .A1_f (new_AGEMA_signal_3683), .B0_t (1'b0), .B0_f (1'b1), .B1_t (FSM[1]), .B1_f (new_AGEMA_signal_2301), .Z0_t (AddRoundConstantOutput[61]), .Z0_f (new_AGEMA_signal_3792), .Z1_t (new_AGEMA_signal_3793), .Z1_f (new_AGEMA_signal_3794) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_0_2_U1 ( .A0_t (SubCellInst_SboxInst_15_YY[0]), .A0_f (new_AGEMA_signal_2842), .A1_t (new_AGEMA_signal_2843), .A1_f (new_AGEMA_signal_2844), .B0_t (1'b0), .B0_f (1'b1), .B1_t (FSMUpdate[3]), .B1_f (new_AGEMA_signal_2302), .Z0_t (AddRoundConstantOutput[62]), .Z0_f (new_AGEMA_signal_2993), .Z1_t (new_AGEMA_signal_2994), .Z1_f (new_AGEMA_signal_2995) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_0_3_U1 ( .A0_t (SubCellInst_SboxInst_15_YY[1]), .A0_f (new_AGEMA_signal_3179), .A1_t (new_AGEMA_signal_3180), .A1_f (new_AGEMA_signal_3181), .B0_t (1'b0), .B0_f (1'b1), .B1_t (FSMUpdate[4]), .B1_f (new_AGEMA_signal_2303), .Z0_t (AddRoundConstantOutput[63]), .Z0_f (new_AGEMA_signal_3323), .Z1_t (new_AGEMA_signal_3324), .Z1_f (new_AGEMA_signal_3325) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_1_0_U1 ( .A0_t (SubCellOutput[44]), .A0_f (new_AGEMA_signal_3498), .A1_t (new_AGEMA_signal_3499), .A1_f (new_AGEMA_signal_3500), .B0_t (1'b0), .B0_f (1'b1), .B1_t (FSM[4]), .B1_f (new_AGEMA_signal_2304), .Z0_t (AddRoundConstantOutput[44]), .Z0_f (new_AGEMA_signal_3687), .Z1_t (new_AGEMA_signal_3688), .Z1_f (new_AGEMA_signal_3689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_1_1_U1 ( .A0_t (SubCellOutput[45]), .A0_f (new_AGEMA_signal_3669), .A1_t (new_AGEMA_signal_3670), .A1_f (new_AGEMA_signal_3671), .B0_t (1'b0), .B0_f (1'b1), .B1_t (FSM[5]), .B1_f (new_AGEMA_signal_2309), .Z0_t (AddRoundConstantOutput[45]), .Z0_f (new_AGEMA_signal_3795), .Z1_t (new_AGEMA_signal_3796), .Z1_f (new_AGEMA_signal_3797) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_0_0_U1 ( .A0_t (AddRoundConstantOutput[32]), .A0_f (new_AGEMA_signal_3480), .A1_t (new_AGEMA_signal_3481), .A1_f (new_AGEMA_signal_3482), .B0_t (TweakeyGeneration_key_Feedback[0]), .B0_f (new_AGEMA_signal_1723), .B1_t (new_AGEMA_signal_1724), .B1_f (new_AGEMA_signal_1725), .Z0_t (ShiftRowsOutput[44]), .Z0_f (new_AGEMA_signal_3690), .Z1_t (new_AGEMA_signal_3691), .Z1_f (new_AGEMA_signal_3692) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_0_1_U1 ( .A0_t (AddRoundConstantOutput[33]), .A0_f (new_AGEMA_signal_3660), .A1_t (new_AGEMA_signal_3661), .A1_f (new_AGEMA_signal_3662), .B0_t (TweakeyGeneration_key_Feedback[1]), .B0_f (new_AGEMA_signal_1732), .B1_t (new_AGEMA_signal_1733), .B1_f (new_AGEMA_signal_1734), .Z0_t (ShiftRowsOutput[45]), .Z0_f (new_AGEMA_signal_3798), .Z1_t (new_AGEMA_signal_3799), .Z1_f (new_AGEMA_signal_3800) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_0_2_U1 ( .A0_t (SubCellInst_SboxInst_8_YY[0]), .A0_f (new_AGEMA_signal_2779), .A1_t (new_AGEMA_signal_2780), .A1_f (new_AGEMA_signal_2781), .B0_t (TweakeyGeneration_key_Feedback[2]), .B0_f (new_AGEMA_signal_1741), .B1_t (new_AGEMA_signal_1742), .B1_f (new_AGEMA_signal_1743), .Z0_t (ShiftRowsOutput[46]), .Z0_f (new_AGEMA_signal_2996), .Z1_t (new_AGEMA_signal_2997), .Z1_f (new_AGEMA_signal_2998) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_0_3_U1 ( .A0_t (SubCellInst_SboxInst_8_YY[1]), .A0_f (new_AGEMA_signal_3116), .A1_t (new_AGEMA_signal_3117), .A1_f (new_AGEMA_signal_3118), .B0_t (TweakeyGeneration_key_Feedback[3]), .B0_f (new_AGEMA_signal_1750), .B1_t (new_AGEMA_signal_1751), .B1_f (new_AGEMA_signal_1752), .Z0_t (ShiftRowsOutput[47]), .Z0_f (new_AGEMA_signal_3326), .Z1_t (new_AGEMA_signal_3327), .Z1_f (new_AGEMA_signal_3328) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_1_0_U1 ( .A0_t (AddRoundConstantOutput[36]), .A0_f (new_AGEMA_signal_3486), .A1_t (new_AGEMA_signal_3487), .A1_f (new_AGEMA_signal_3488), .B0_t (TweakeyGeneration_key_Feedback[4]), .B0_f (new_AGEMA_signal_1759), .B1_t (new_AGEMA_signal_1760), .B1_f (new_AGEMA_signal_1761), .Z0_t (ShiftRowsOutput[32]), .Z0_f (new_AGEMA_signal_3693), .Z1_t (new_AGEMA_signal_3694), .Z1_f (new_AGEMA_signal_3695) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_1_1_U1 ( .A0_t (AddRoundConstantOutput[37]), .A0_f (new_AGEMA_signal_3663), .A1_t (new_AGEMA_signal_3664), .A1_f (new_AGEMA_signal_3665), .B0_t (TweakeyGeneration_key_Feedback[5]), .B0_f (new_AGEMA_signal_1768), .B1_t (new_AGEMA_signal_1769), .B1_f (new_AGEMA_signal_1770), .Z0_t (ShiftRowsOutput[33]), .Z0_f (new_AGEMA_signal_3801), .Z1_t (new_AGEMA_signal_3802), .Z1_f (new_AGEMA_signal_3803) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_1_2_U1 ( .A0_t (SubCellInst_SboxInst_9_YY[0]), .A0_f (new_AGEMA_signal_2788), .A1_t (new_AGEMA_signal_2789), .A1_f (new_AGEMA_signal_2790), .B0_t (TweakeyGeneration_key_Feedback[6]), .B0_f (new_AGEMA_signal_1777), .B1_t (new_AGEMA_signal_1778), .B1_f (new_AGEMA_signal_1779), .Z0_t (ShiftRowsOutput[34]), .Z0_f (new_AGEMA_signal_2999), .Z1_t (new_AGEMA_signal_3000), .Z1_f (new_AGEMA_signal_3001) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_1_3_U1 ( .A0_t (SubCellInst_SboxInst_9_YY[1]), .A0_f (new_AGEMA_signal_3125), .A1_t (new_AGEMA_signal_3126), .A1_f (new_AGEMA_signal_3127), .B0_t (TweakeyGeneration_key_Feedback[7]), .B0_f (new_AGEMA_signal_1786), .B1_t (new_AGEMA_signal_1787), .B1_f (new_AGEMA_signal_1788), .Z0_t (ShiftRowsOutput[35]), .Z0_f (new_AGEMA_signal_3329), .Z1_t (new_AGEMA_signal_3330), .Z1_f (new_AGEMA_signal_3331) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_2_0_U1 ( .A0_t (AddRoundConstantOutput[40]), .A0_f (new_AGEMA_signal_3492), .A1_t (new_AGEMA_signal_3493), .A1_f (new_AGEMA_signal_3494), .B0_t (TweakeyGeneration_key_Feedback[8]), .B0_f (new_AGEMA_signal_1795), .B1_t (new_AGEMA_signal_1796), .B1_f (new_AGEMA_signal_1797), .Z0_t (ShiftRowsOutput[36]), .Z0_f (new_AGEMA_signal_3696), .Z1_t (new_AGEMA_signal_3697), .Z1_f (new_AGEMA_signal_3698) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_2_1_U1 ( .A0_t (AddRoundConstantOutput[41]), .A0_f (new_AGEMA_signal_3666), .A1_t (new_AGEMA_signal_3667), .A1_f (new_AGEMA_signal_3668), .B0_t (TweakeyGeneration_key_Feedback[9]), .B0_f (new_AGEMA_signal_1804), .B1_t (new_AGEMA_signal_1805), .B1_f (new_AGEMA_signal_1806), .Z0_t (ShiftRowsOutput[37]), .Z0_f (new_AGEMA_signal_3804), .Z1_t (new_AGEMA_signal_3805), .Z1_f (new_AGEMA_signal_3806) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_2_2_U1 ( .A0_t (SubCellInst_SboxInst_10_YY[0]), .A0_f (new_AGEMA_signal_2797), .A1_t (new_AGEMA_signal_2798), .A1_f (new_AGEMA_signal_2799), .B0_t (TweakeyGeneration_key_Feedback[10]), .B0_f (new_AGEMA_signal_1813), .B1_t (new_AGEMA_signal_1814), .B1_f (new_AGEMA_signal_1815), .Z0_t (ShiftRowsOutput[38]), .Z0_f (new_AGEMA_signal_3002), .Z1_t (new_AGEMA_signal_3003), .Z1_f (new_AGEMA_signal_3004) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_2_3_U1 ( .A0_t (SubCellInst_SboxInst_10_YY[1]), .A0_f (new_AGEMA_signal_3134), .A1_t (new_AGEMA_signal_3135), .A1_f (new_AGEMA_signal_3136), .B0_t (TweakeyGeneration_key_Feedback[11]), .B0_f (new_AGEMA_signal_1822), .B1_t (new_AGEMA_signal_1823), .B1_f (new_AGEMA_signal_1824), .Z0_t (ShiftRowsOutput[39]), .Z0_f (new_AGEMA_signal_3332), .Z1_t (new_AGEMA_signal_3333), .Z1_f (new_AGEMA_signal_3334) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_3_0_U1 ( .A0_t (AddRoundConstantOutput[44]), .A0_f (new_AGEMA_signal_3687), .A1_t (new_AGEMA_signal_3688), .A1_f (new_AGEMA_signal_3689), .B0_t (TweakeyGeneration_key_Feedback[12]), .B0_f (new_AGEMA_signal_1831), .B1_t (new_AGEMA_signal_1832), .B1_f (new_AGEMA_signal_1833), .Z0_t (ShiftRowsOutput[40]), .Z0_f (new_AGEMA_signal_3807), .Z1_t (new_AGEMA_signal_3808), .Z1_f (new_AGEMA_signal_3809) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_3_1_U1 ( .A0_t (AddRoundConstantOutput[45]), .A0_f (new_AGEMA_signal_3795), .A1_t (new_AGEMA_signal_3796), .A1_f (new_AGEMA_signal_3797), .B0_t (TweakeyGeneration_key_Feedback[13]), .B0_f (new_AGEMA_signal_1840), .B1_t (new_AGEMA_signal_1841), .B1_f (new_AGEMA_signal_1842), .Z0_t (ShiftRowsOutput[41]), .Z0_f (new_AGEMA_signal_3939), .Z1_t (new_AGEMA_signal_3940), .Z1_f (new_AGEMA_signal_3941) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_3_2_U1 ( .A0_t (SubCellInst_SboxInst_11_YY[0]), .A0_f (new_AGEMA_signal_2806), .A1_t (new_AGEMA_signal_2807), .A1_f (new_AGEMA_signal_2808), .B0_t (TweakeyGeneration_key_Feedback[14]), .B0_f (new_AGEMA_signal_1849), .B1_t (new_AGEMA_signal_1850), .B1_f (new_AGEMA_signal_1851), .Z0_t (ShiftRowsOutput[42]), .Z0_f (new_AGEMA_signal_3005), .Z1_t (new_AGEMA_signal_3006), .Z1_f (new_AGEMA_signal_3007) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_3_3_U1 ( .A0_t (SubCellInst_SboxInst_11_YY[1]), .A0_f (new_AGEMA_signal_3143), .A1_t (new_AGEMA_signal_3144), .A1_f (new_AGEMA_signal_3145), .B0_t (TweakeyGeneration_key_Feedback[15]), .B0_f (new_AGEMA_signal_1858), .B1_t (new_AGEMA_signal_1859), .B1_f (new_AGEMA_signal_1860), .Z0_t (ShiftRowsOutput[43]), .Z0_f (new_AGEMA_signal_3335), .Z1_t (new_AGEMA_signal_3336), .Z1_f (new_AGEMA_signal_3337) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_4_0_U1 ( .A0_t (AddRoundConstantOutput[48]), .A0_f (new_AGEMA_signal_3504), .A1_t (new_AGEMA_signal_3505), .A1_f (new_AGEMA_signal_3506), .B0_t (TweakeyGeneration_key_Feedback[16]), .B0_f (new_AGEMA_signal_1867), .B1_t (new_AGEMA_signal_1868), .B1_f (new_AGEMA_signal_1869), .Z0_t (MCOutput[32]), .Z0_f (new_AGEMA_signal_3699), .Z1_t (new_AGEMA_signal_3700), .Z1_f (new_AGEMA_signal_3701) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_4_1_U1 ( .A0_t (AddRoundConstantOutput[49]), .A0_f (new_AGEMA_signal_3672), .A1_t (new_AGEMA_signal_3673), .A1_f (new_AGEMA_signal_3674), .B0_t (TweakeyGeneration_key_Feedback[17]), .B0_f (new_AGEMA_signal_1876), .B1_t (new_AGEMA_signal_1877), .B1_f (new_AGEMA_signal_1878), .Z0_t (MCOutput[33]), .Z0_f (new_AGEMA_signal_3810), .Z1_t (new_AGEMA_signal_3811), .Z1_f (new_AGEMA_signal_3812) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_4_2_U1 ( .A0_t (SubCellInst_SboxInst_12_YY[0]), .A0_f (new_AGEMA_signal_2815), .A1_t (new_AGEMA_signal_2816), .A1_f (new_AGEMA_signal_2817), .B0_t (TweakeyGeneration_key_Feedback[18]), .B0_f (new_AGEMA_signal_1885), .B1_t (new_AGEMA_signal_1886), .B1_f (new_AGEMA_signal_1887), .Z0_t (MCOutput[34]), .Z0_f (new_AGEMA_signal_3008), .Z1_t (new_AGEMA_signal_3009), .Z1_f (new_AGEMA_signal_3010) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_4_3_U1 ( .A0_t (SubCellInst_SboxInst_12_YY[1]), .A0_f (new_AGEMA_signal_3152), .A1_t (new_AGEMA_signal_3153), .A1_f (new_AGEMA_signal_3154), .B0_t (TweakeyGeneration_key_Feedback[19]), .B0_f (new_AGEMA_signal_1894), .B1_t (new_AGEMA_signal_1895), .B1_f (new_AGEMA_signal_1896), .Z0_t (MCOutput[35]), .Z0_f (new_AGEMA_signal_3338), .Z1_t (new_AGEMA_signal_3339), .Z1_f (new_AGEMA_signal_3340) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_5_0_U1 ( .A0_t (AddRoundConstantOutput[52]), .A0_f (new_AGEMA_signal_3510), .A1_t (new_AGEMA_signal_3511), .A1_f (new_AGEMA_signal_3512), .B0_t (TweakeyGeneration_key_Feedback[20]), .B0_f (new_AGEMA_signal_1903), .B1_t (new_AGEMA_signal_1904), .B1_f (new_AGEMA_signal_1905), .Z0_t (MCOutput[36]), .Z0_f (new_AGEMA_signal_3702), .Z1_t (new_AGEMA_signal_3703), .Z1_f (new_AGEMA_signal_3704) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_5_1_U1 ( .A0_t (AddRoundConstantOutput[53]), .A0_f (new_AGEMA_signal_3675), .A1_t (new_AGEMA_signal_3676), .A1_f (new_AGEMA_signal_3677), .B0_t (TweakeyGeneration_key_Feedback[21]), .B0_f (new_AGEMA_signal_1912), .B1_t (new_AGEMA_signal_1913), .B1_f (new_AGEMA_signal_1914), .Z0_t (MCOutput[37]), .Z0_f (new_AGEMA_signal_3813), .Z1_t (new_AGEMA_signal_3814), .Z1_f (new_AGEMA_signal_3815) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_5_2_U1 ( .A0_t (SubCellInst_SboxInst_13_YY[0]), .A0_f (new_AGEMA_signal_2824), .A1_t (new_AGEMA_signal_2825), .A1_f (new_AGEMA_signal_2826), .B0_t (TweakeyGeneration_key_Feedback[22]), .B0_f (new_AGEMA_signal_1921), .B1_t (new_AGEMA_signal_1922), .B1_f (new_AGEMA_signal_1923), .Z0_t (MCOutput[38]), .Z0_f (new_AGEMA_signal_3011), .Z1_t (new_AGEMA_signal_3012), .Z1_f (new_AGEMA_signal_3013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_5_3_U1 ( .A0_t (SubCellInst_SboxInst_13_YY[1]), .A0_f (new_AGEMA_signal_3161), .A1_t (new_AGEMA_signal_3162), .A1_f (new_AGEMA_signal_3163), .B0_t (TweakeyGeneration_key_Feedback[23]), .B0_f (new_AGEMA_signal_1930), .B1_t (new_AGEMA_signal_1931), .B1_f (new_AGEMA_signal_1932), .Z0_t (MCOutput[39]), .Z0_f (new_AGEMA_signal_3341), .Z1_t (new_AGEMA_signal_3342), .Z1_f (new_AGEMA_signal_3343) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_6_0_U1 ( .A0_t (AddRoundConstantOutput[56]), .A0_f (new_AGEMA_signal_3516), .A1_t (new_AGEMA_signal_3517), .A1_f (new_AGEMA_signal_3518), .B0_t (TweakeyGeneration_key_Feedback[24]), .B0_f (new_AGEMA_signal_1939), .B1_t (new_AGEMA_signal_1940), .B1_f (new_AGEMA_signal_1941), .Z0_t (MCOutput[40]), .Z0_f (new_AGEMA_signal_3705), .Z1_t (new_AGEMA_signal_3706), .Z1_f (new_AGEMA_signal_3707) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_6_1_U1 ( .A0_t (AddRoundConstantOutput[57]), .A0_f (new_AGEMA_signal_3678), .A1_t (new_AGEMA_signal_3679), .A1_f (new_AGEMA_signal_3680), .B0_t (TweakeyGeneration_key_Feedback[25]), .B0_f (new_AGEMA_signal_1948), .B1_t (new_AGEMA_signal_1949), .B1_f (new_AGEMA_signal_1950), .Z0_t (MCOutput[41]), .Z0_f (new_AGEMA_signal_3816), .Z1_t (new_AGEMA_signal_3817), .Z1_f (new_AGEMA_signal_3818) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_6_2_U1 ( .A0_t (SubCellInst_SboxInst_14_YY[0]), .A0_f (new_AGEMA_signal_2833), .A1_t (new_AGEMA_signal_2834), .A1_f (new_AGEMA_signal_2835), .B0_t (TweakeyGeneration_key_Feedback[26]), .B0_f (new_AGEMA_signal_1957), .B1_t (new_AGEMA_signal_1958), .B1_f (new_AGEMA_signal_1959), .Z0_t (MCOutput[42]), .Z0_f (new_AGEMA_signal_3014), .Z1_t (new_AGEMA_signal_3015), .Z1_f (new_AGEMA_signal_3016) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_6_3_U1 ( .A0_t (SubCellInst_SboxInst_14_YY[1]), .A0_f (new_AGEMA_signal_3170), .A1_t (new_AGEMA_signal_3171), .A1_f (new_AGEMA_signal_3172), .B0_t (TweakeyGeneration_key_Feedback[27]), .B0_f (new_AGEMA_signal_1966), .B1_t (new_AGEMA_signal_1967), .B1_f (new_AGEMA_signal_1968), .Z0_t (MCOutput[43]), .Z0_f (new_AGEMA_signal_3344), .Z1_t (new_AGEMA_signal_3345), .Z1_f (new_AGEMA_signal_3346) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_7_0_U1 ( .A0_t (AddRoundConstantOutput[60]), .A0_f (new_AGEMA_signal_3684), .A1_t (new_AGEMA_signal_3685), .A1_f (new_AGEMA_signal_3686), .B0_t (TweakeyGeneration_key_Feedback[28]), .B0_f (new_AGEMA_signal_1975), .B1_t (new_AGEMA_signal_1976), .B1_f (new_AGEMA_signal_1977), .Z0_t (MCOutput[44]), .Z0_f (new_AGEMA_signal_3819), .Z1_t (new_AGEMA_signal_3820), .Z1_f (new_AGEMA_signal_3821) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_7_1_U1 ( .A0_t (AddRoundConstantOutput[61]), .A0_f (new_AGEMA_signal_3792), .A1_t (new_AGEMA_signal_3793), .A1_f (new_AGEMA_signal_3794), .B0_t (TweakeyGeneration_key_Feedback[29]), .B0_f (new_AGEMA_signal_1984), .B1_t (new_AGEMA_signal_1985), .B1_f (new_AGEMA_signal_1986), .Z0_t (MCOutput[45]), .Z0_f (new_AGEMA_signal_3942), .Z1_t (new_AGEMA_signal_3943), .Z1_f (new_AGEMA_signal_3944) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_7_2_U1 ( .A0_t (AddRoundConstantOutput[62]), .A0_f (new_AGEMA_signal_2993), .A1_t (new_AGEMA_signal_2994), .A1_f (new_AGEMA_signal_2995), .B0_t (TweakeyGeneration_key_Feedback[30]), .B0_f (new_AGEMA_signal_1993), .B1_t (new_AGEMA_signal_1994), .B1_f (new_AGEMA_signal_1995), .Z0_t (MCOutput[46]), .Z0_f (new_AGEMA_signal_3182), .Z1_t (new_AGEMA_signal_3183), .Z1_f (new_AGEMA_signal_3184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_7_3_U1 ( .A0_t (AddRoundConstantOutput[63]), .A0_f (new_AGEMA_signal_3323), .A1_t (new_AGEMA_signal_3324), .A1_f (new_AGEMA_signal_3325), .B0_t (TweakeyGeneration_key_Feedback[31]), .B0_f (new_AGEMA_signal_2002), .B1_t (new_AGEMA_signal_2003), .B1_f (new_AGEMA_signal_2004), .Z0_t (MCOutput[47]), .Z0_f (new_AGEMA_signal_3525), .Z1_t (new_AGEMA_signal_3526), .Z1_f (new_AGEMA_signal_3527) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_0_U2 ( .A0_t (MCInst_MCR0_XORInst_0_0_n1), .A0_f (new_AGEMA_signal_3822), .A1_t (new_AGEMA_signal_3823), .A1_f (new_AGEMA_signal_3824), .B0_t (ShiftRowsOutput[0]), .B0_f (new_AGEMA_signal_3450), .B1_t (new_AGEMA_signal_3451), .B1_f (new_AGEMA_signal_3452), .Z0_t (MCOutput[48]), .Z0_f (new_AGEMA_signal_3945), .Z1_t (new_AGEMA_signal_3946), .Z1_f (new_AGEMA_signal_3947) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_0_U1 ( .A0_t (MCOutput[32]), .A0_f (new_AGEMA_signal_3699), .A1_t (new_AGEMA_signal_3700), .A1_f (new_AGEMA_signal_3701), .B0_t (ShiftRowsOutput[16]), .B0_f (new_AGEMA_signal_3468), .B1_t (new_AGEMA_signal_3469), .B1_f (new_AGEMA_signal_3470), .Z0_t (MCInst_MCR0_XORInst_0_0_n1), .Z0_f (new_AGEMA_signal_3822), .Z1_t (new_AGEMA_signal_3823), .Z1_f (new_AGEMA_signal_3824) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_1_U2 ( .A0_t (MCInst_MCR0_XORInst_0_1_n1), .A0_f (new_AGEMA_signal_3948), .A1_t (new_AGEMA_signal_3949), .A1_f (new_AGEMA_signal_3950), .B0_t (ShiftRowsOutput[1]), .B0_f (new_AGEMA_signal_3645), .B1_t (new_AGEMA_signal_3646), .B1_f (new_AGEMA_signal_3647), .Z0_t (MCOutput[49]), .Z0_f (new_AGEMA_signal_4095), .Z1_t (new_AGEMA_signal_4096), .Z1_f (new_AGEMA_signal_4097) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_1_U1 ( .A0_t (MCOutput[33]), .A0_f (new_AGEMA_signal_3810), .A1_t (new_AGEMA_signal_3811), .A1_f (new_AGEMA_signal_3812), .B0_t (ShiftRowsOutput[17]), .B0_f (new_AGEMA_signal_3654), .B1_t (new_AGEMA_signal_3655), .B1_f (new_AGEMA_signal_3656), .Z0_t (MCInst_MCR0_XORInst_0_1_n1), .Z0_f (new_AGEMA_signal_3948), .Z1_t (new_AGEMA_signal_3949), .Z1_f (new_AGEMA_signal_3950) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_2_U2 ( .A0_t (MCInst_MCR0_XORInst_0_2_n1), .A0_f (new_AGEMA_signal_3185), .A1_t (new_AGEMA_signal_3186), .A1_f (new_AGEMA_signal_3187), .B0_t (SubCellInst_SboxInst_3_YY[0]), .B0_f (new_AGEMA_signal_2734), .B1_t (new_AGEMA_signal_2735), .B1_f (new_AGEMA_signal_2736), .Z0_t (MCOutput[50]), .Z0_f (new_AGEMA_signal_3347), .Z1_t (new_AGEMA_signal_3348), .Z1_f (new_AGEMA_signal_3349) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_2_U1 ( .A0_t (MCOutput[34]), .A0_f (new_AGEMA_signal_3008), .A1_t (new_AGEMA_signal_3009), .A1_f (new_AGEMA_signal_3010), .B0_t (SubCellInst_SboxInst_6_YY[0]), .B0_f (new_AGEMA_signal_2761), .B1_t (new_AGEMA_signal_2762), .B1_f (new_AGEMA_signal_2763), .Z0_t (MCInst_MCR0_XORInst_0_2_n1), .Z0_f (new_AGEMA_signal_3185), .Z1_t (new_AGEMA_signal_3186), .Z1_f (new_AGEMA_signal_3187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_3_U2 ( .A0_t (MCInst_MCR0_XORInst_0_3_n1), .A0_f (new_AGEMA_signal_3528), .A1_t (new_AGEMA_signal_3529), .A1_f (new_AGEMA_signal_3530), .B0_t (SubCellInst_SboxInst_3_YY[1]), .B0_f (new_AGEMA_signal_3071), .B1_t (new_AGEMA_signal_3072), .B1_f (new_AGEMA_signal_3073), .Z0_t (MCOutput[51]), .Z0_f (new_AGEMA_signal_3708), .Z1_t (new_AGEMA_signal_3709), .Z1_f (new_AGEMA_signal_3710) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_3_U1 ( .A0_t (MCOutput[35]), .A0_f (new_AGEMA_signal_3338), .A1_t (new_AGEMA_signal_3339), .A1_f (new_AGEMA_signal_3340), .B0_t (SubCellInst_SboxInst_6_YY[1]), .B0_f (new_AGEMA_signal_3098), .B1_t (new_AGEMA_signal_3099), .B1_f (new_AGEMA_signal_3100), .Z0_t (MCInst_MCR0_XORInst_0_3_n1), .Z0_f (new_AGEMA_signal_3528), .Z1_t (new_AGEMA_signal_3529), .Z1_f (new_AGEMA_signal_3530) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_0_U2 ( .A0_t (MCInst_MCR0_XORInst_1_0_n1), .A0_f (new_AGEMA_signal_3825), .A1_t (new_AGEMA_signal_3826), .A1_f (new_AGEMA_signal_3827), .B0_t (ShiftRowsOutput[4]), .B0_f (new_AGEMA_signal_3432), .B1_t (new_AGEMA_signal_3433), .B1_f (new_AGEMA_signal_3434), .Z0_t (MCOutput[52]), .Z0_f (new_AGEMA_signal_3951), .Z1_t (new_AGEMA_signal_3952), .Z1_f (new_AGEMA_signal_3953) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_0_U1 ( .A0_t (MCOutput[36]), .A0_f (new_AGEMA_signal_3702), .A1_t (new_AGEMA_signal_3703), .A1_f (new_AGEMA_signal_3704), .B0_t (ShiftRowsOutput[20]), .B0_f (new_AGEMA_signal_3474), .B1_t (new_AGEMA_signal_3475), .B1_f (new_AGEMA_signal_3476), .Z0_t (MCInst_MCR0_XORInst_1_0_n1), .Z0_f (new_AGEMA_signal_3825), .Z1_t (new_AGEMA_signal_3826), .Z1_f (new_AGEMA_signal_3827) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_1_U2 ( .A0_t (MCInst_MCR0_XORInst_1_1_n1), .A0_f (new_AGEMA_signal_3954), .A1_t (new_AGEMA_signal_3955), .A1_f (new_AGEMA_signal_3956), .B0_t (ShiftRowsOutput[5]), .B0_f (new_AGEMA_signal_3636), .B1_t (new_AGEMA_signal_3637), .B1_f (new_AGEMA_signal_3638), .Z0_t (MCOutput[53]), .Z0_f (new_AGEMA_signal_4098), .Z1_t (new_AGEMA_signal_4099), .Z1_f (new_AGEMA_signal_4100) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_1_U1 ( .A0_t (MCOutput[37]), .A0_f (new_AGEMA_signal_3813), .A1_t (new_AGEMA_signal_3814), .A1_f (new_AGEMA_signal_3815), .B0_t (SubCellOutput[29]), .B0_f (new_AGEMA_signal_3657), .B1_t (new_AGEMA_signal_3658), .B1_f (new_AGEMA_signal_3659), .Z0_t (MCInst_MCR0_XORInst_1_1_n1), .Z0_f (new_AGEMA_signal_3954), .Z1_t (new_AGEMA_signal_3955), .Z1_f (new_AGEMA_signal_3956) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_2_U2 ( .A0_t (MCInst_MCR0_XORInst_1_2_n1), .A0_f (new_AGEMA_signal_3188), .A1_t (new_AGEMA_signal_3189), .A1_f (new_AGEMA_signal_3190), .B0_t (SubCellInst_SboxInst_0_YY[0]), .B0_f (new_AGEMA_signal_2707), .B1_t (new_AGEMA_signal_2708), .B1_f (new_AGEMA_signal_2709), .Z0_t (MCOutput[54]), .Z0_f (new_AGEMA_signal_3350), .Z1_t (new_AGEMA_signal_3351), .Z1_f (new_AGEMA_signal_3352) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_2_U1 ( .A0_t (MCOutput[38]), .A0_f (new_AGEMA_signal_3011), .A1_t (new_AGEMA_signal_3012), .A1_f (new_AGEMA_signal_3013), .B0_t (SubCellInst_SboxInst_7_YY[0]), .B0_f (new_AGEMA_signal_2770), .B1_t (new_AGEMA_signal_2771), .B1_f (new_AGEMA_signal_2772), .Z0_t (MCInst_MCR0_XORInst_1_2_n1), .Z0_f (new_AGEMA_signal_3188), .Z1_t (new_AGEMA_signal_3189), .Z1_f (new_AGEMA_signal_3190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_3_U2 ( .A0_t (MCInst_MCR0_XORInst_1_3_n1), .A0_f (new_AGEMA_signal_3531), .A1_t (new_AGEMA_signal_3532), .A1_f (new_AGEMA_signal_3533), .B0_t (SubCellInst_SboxInst_0_YY[1]), .B0_f (new_AGEMA_signal_3044), .B1_t (new_AGEMA_signal_3045), .B1_f (new_AGEMA_signal_3046), .Z0_t (MCOutput[55]), .Z0_f (new_AGEMA_signal_3711), .Z1_t (new_AGEMA_signal_3712), .Z1_f (new_AGEMA_signal_3713) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_3_U1 ( .A0_t (MCOutput[39]), .A0_f (new_AGEMA_signal_3341), .A1_t (new_AGEMA_signal_3342), .A1_f (new_AGEMA_signal_3343), .B0_t (SubCellInst_SboxInst_7_YY[1]), .B0_f (new_AGEMA_signal_3107), .B1_t (new_AGEMA_signal_3108), .B1_f (new_AGEMA_signal_3109), .Z0_t (MCInst_MCR0_XORInst_1_3_n1), .Z0_f (new_AGEMA_signal_3531), .Z1_t (new_AGEMA_signal_3532), .Z1_f (new_AGEMA_signal_3533) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_0_U2 ( .A0_t (MCInst_MCR0_XORInst_2_0_n1), .A0_f (new_AGEMA_signal_3828), .A1_t (new_AGEMA_signal_3829), .A1_f (new_AGEMA_signal_3830), .B0_t (ShiftRowsOutput[8]), .B0_f (new_AGEMA_signal_3438), .B1_t (new_AGEMA_signal_3439), .B1_f (new_AGEMA_signal_3440), .Z0_t (MCOutput[56]), .Z0_f (new_AGEMA_signal_3957), .Z1_t (new_AGEMA_signal_3958), .Z1_f (new_AGEMA_signal_3959) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_0_U1 ( .A0_t (MCOutput[40]), .A0_f (new_AGEMA_signal_3705), .A1_t (new_AGEMA_signal_3706), .A1_f (new_AGEMA_signal_3707), .B0_t (ShiftRowsOutput[24]), .B0_f (new_AGEMA_signal_3456), .B1_t (new_AGEMA_signal_3457), .B1_f (new_AGEMA_signal_3458), .Z0_t (MCInst_MCR0_XORInst_2_0_n1), .Z0_f (new_AGEMA_signal_3828), .Z1_t (new_AGEMA_signal_3829), .Z1_f (new_AGEMA_signal_3830) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_1_U2 ( .A0_t (MCInst_MCR0_XORInst_2_1_n1), .A0_f (new_AGEMA_signal_3960), .A1_t (new_AGEMA_signal_3961), .A1_f (new_AGEMA_signal_3962), .B0_t (ShiftRowsOutput[9]), .B0_f (new_AGEMA_signal_3639), .B1_t (new_AGEMA_signal_3640), .B1_f (new_AGEMA_signal_3641), .Z0_t (MCOutput[57]), .Z0_f (new_AGEMA_signal_4101), .Z1_t (new_AGEMA_signal_4102), .Z1_f (new_AGEMA_signal_4103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_1_U1 ( .A0_t (MCOutput[41]), .A0_f (new_AGEMA_signal_3816), .A1_t (new_AGEMA_signal_3817), .A1_f (new_AGEMA_signal_3818), .B0_t (ShiftRowsOutput[25]), .B0_f (new_AGEMA_signal_3648), .B1_t (new_AGEMA_signal_3649), .B1_f (new_AGEMA_signal_3650), .Z0_t (MCInst_MCR0_XORInst_2_1_n1), .Z0_f (new_AGEMA_signal_3960), .Z1_t (new_AGEMA_signal_3961), .Z1_f (new_AGEMA_signal_3962) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_2_U2 ( .A0_t (MCInst_MCR0_XORInst_2_2_n1), .A0_f (new_AGEMA_signal_3191), .A1_t (new_AGEMA_signal_3192), .A1_f (new_AGEMA_signal_3193), .B0_t (SubCellInst_SboxInst_1_YY[0]), .B0_f (new_AGEMA_signal_2716), .B1_t (new_AGEMA_signal_2717), .B1_f (new_AGEMA_signal_2718), .Z0_t (MCOutput[58]), .Z0_f (new_AGEMA_signal_3353), .Z1_t (new_AGEMA_signal_3354), .Z1_f (new_AGEMA_signal_3355) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_2_U1 ( .A0_t (MCOutput[42]), .A0_f (new_AGEMA_signal_3014), .A1_t (new_AGEMA_signal_3015), .A1_f (new_AGEMA_signal_3016), .B0_t (SubCellInst_SboxInst_4_YY[0]), .B0_f (new_AGEMA_signal_2743), .B1_t (new_AGEMA_signal_2744), .B1_f (new_AGEMA_signal_2745), .Z0_t (MCInst_MCR0_XORInst_2_2_n1), .Z0_f (new_AGEMA_signal_3191), .Z1_t (new_AGEMA_signal_3192), .Z1_f (new_AGEMA_signal_3193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_3_U2 ( .A0_t (MCInst_MCR0_XORInst_2_3_n1), .A0_f (new_AGEMA_signal_3534), .A1_t (new_AGEMA_signal_3535), .A1_f (new_AGEMA_signal_3536), .B0_t (SubCellInst_SboxInst_1_YY[1]), .B0_f (new_AGEMA_signal_3053), .B1_t (new_AGEMA_signal_3054), .B1_f (new_AGEMA_signal_3055), .Z0_t (MCOutput[59]), .Z0_f (new_AGEMA_signal_3714), .Z1_t (new_AGEMA_signal_3715), .Z1_f (new_AGEMA_signal_3716) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_3_U1 ( .A0_t (MCOutput[43]), .A0_f (new_AGEMA_signal_3344), .A1_t (new_AGEMA_signal_3345), .A1_f (new_AGEMA_signal_3346), .B0_t (SubCellInst_SboxInst_4_YY[1]), .B0_f (new_AGEMA_signal_3080), .B1_t (new_AGEMA_signal_3081), .B1_f (new_AGEMA_signal_3082), .Z0_t (MCInst_MCR0_XORInst_2_3_n1), .Z0_f (new_AGEMA_signal_3534), .Z1_t (new_AGEMA_signal_3535), .Z1_f (new_AGEMA_signal_3536) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_0_U2 ( .A0_t (MCInst_MCR0_XORInst_3_0_n1), .A0_f (new_AGEMA_signal_3963), .A1_t (new_AGEMA_signal_3964), .A1_f (new_AGEMA_signal_3965), .B0_t (ShiftRowsOutput[12]), .B0_f (new_AGEMA_signal_3444), .B1_t (new_AGEMA_signal_3445), .B1_f (new_AGEMA_signal_3446), .Z0_t (MCOutput[60]), .Z0_f (new_AGEMA_signal_4104), .Z1_t (new_AGEMA_signal_4105), .Z1_f (new_AGEMA_signal_4106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_0_U1 ( .A0_t (MCOutput[44]), .A0_f (new_AGEMA_signal_3819), .A1_t (new_AGEMA_signal_3820), .A1_f (new_AGEMA_signal_3821), .B0_t (ShiftRowsOutput[28]), .B0_f (new_AGEMA_signal_3462), .B1_t (new_AGEMA_signal_3463), .B1_f (new_AGEMA_signal_3464), .Z0_t (MCInst_MCR0_XORInst_3_0_n1), .Z0_f (new_AGEMA_signal_3963), .Z1_t (new_AGEMA_signal_3964), .Z1_f (new_AGEMA_signal_3965) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_1_U2 ( .A0_t (MCInst_MCR0_XORInst_3_1_n1), .A0_f (new_AGEMA_signal_4107), .A1_t (new_AGEMA_signal_4108), .A1_f (new_AGEMA_signal_4109), .B0_t (ShiftRowsOutput[13]), .B0_f (new_AGEMA_signal_3642), .B1_t (new_AGEMA_signal_3643), .B1_f (new_AGEMA_signal_3644), .Z0_t (MCOutput[61]), .Z0_f (new_AGEMA_signal_4188), .Z1_t (new_AGEMA_signal_4189), .Z1_f (new_AGEMA_signal_4190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_1_U1 ( .A0_t (MCOutput[45]), .A0_f (new_AGEMA_signal_3942), .A1_t (new_AGEMA_signal_3943), .A1_f (new_AGEMA_signal_3944), .B0_t (ShiftRowsOutput[29]), .B0_f (new_AGEMA_signal_3651), .B1_t (new_AGEMA_signal_3652), .B1_f (new_AGEMA_signal_3653), .Z0_t (MCInst_MCR0_XORInst_3_1_n1), .Z0_f (new_AGEMA_signal_4107), .Z1_t (new_AGEMA_signal_4108), .Z1_f (new_AGEMA_signal_4109) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_2_U2 ( .A0_t (MCInst_MCR0_XORInst_3_2_n1), .A0_f (new_AGEMA_signal_3356), .A1_t (new_AGEMA_signal_3357), .A1_f (new_AGEMA_signal_3358), .B0_t (SubCellInst_SboxInst_2_YY[0]), .B0_f (new_AGEMA_signal_2725), .B1_t (new_AGEMA_signal_2726), .B1_f (new_AGEMA_signal_2727), .Z0_t (MCOutput[62]), .Z0_f (new_AGEMA_signal_3537), .Z1_t (new_AGEMA_signal_3538), .Z1_f (new_AGEMA_signal_3539) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_2_U1 ( .A0_t (MCOutput[46]), .A0_f (new_AGEMA_signal_3182), .A1_t (new_AGEMA_signal_3183), .A1_f (new_AGEMA_signal_3184), .B0_t (SubCellInst_SboxInst_5_YY[0]), .B0_f (new_AGEMA_signal_2752), .B1_t (new_AGEMA_signal_2753), .B1_f (new_AGEMA_signal_2754), .Z0_t (MCInst_MCR0_XORInst_3_2_n1), .Z0_f (new_AGEMA_signal_3356), .Z1_t (new_AGEMA_signal_3357), .Z1_f (new_AGEMA_signal_3358) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_3_U2 ( .A0_t (MCInst_MCR0_XORInst_3_3_n1), .A0_f (new_AGEMA_signal_3717), .A1_t (new_AGEMA_signal_3718), .A1_f (new_AGEMA_signal_3719), .B0_t (SubCellInst_SboxInst_2_YY[1]), .B0_f (new_AGEMA_signal_3062), .B1_t (new_AGEMA_signal_3063), .B1_f (new_AGEMA_signal_3064), .Z0_t (MCOutput[63]), .Z0_f (new_AGEMA_signal_3831), .Z1_t (new_AGEMA_signal_3832), .Z1_f (new_AGEMA_signal_3833) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_3_U1 ( .A0_t (MCOutput[47]), .A0_f (new_AGEMA_signal_3525), .A1_t (new_AGEMA_signal_3526), .A1_f (new_AGEMA_signal_3527), .B0_t (SubCellInst_SboxInst_5_YY[1]), .B0_f (new_AGEMA_signal_3089), .B1_t (new_AGEMA_signal_3090), .B1_f (new_AGEMA_signal_3091), .Z0_t (MCInst_MCR0_XORInst_3_3_n1), .Z0_f (new_AGEMA_signal_3717), .Z1_t (new_AGEMA_signal_3718), .Z1_f (new_AGEMA_signal_3719) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_0_0_U1 ( .A0_t (ShiftRowsOutput[32]), .A0_f (new_AGEMA_signal_3693), .A1_t (new_AGEMA_signal_3694), .A1_f (new_AGEMA_signal_3695), .B0_t (ShiftRowsOutput[16]), .B0_f (new_AGEMA_signal_3468), .B1_t (new_AGEMA_signal_3469), .B1_f (new_AGEMA_signal_3470), .Z0_t (MCOutput[16]), .Z0_f (new_AGEMA_signal_3834), .Z1_t (new_AGEMA_signal_3835), .Z1_f (new_AGEMA_signal_3836) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_0_1_U1 ( .A0_t (ShiftRowsOutput[33]), .A0_f (new_AGEMA_signal_3801), .A1_t (new_AGEMA_signal_3802), .A1_f (new_AGEMA_signal_3803), .B0_t (ShiftRowsOutput[17]), .B0_f (new_AGEMA_signal_3654), .B1_t (new_AGEMA_signal_3655), .B1_f (new_AGEMA_signal_3656), .Z0_t (MCOutput[17]), .Z0_f (new_AGEMA_signal_3966), .Z1_t (new_AGEMA_signal_3967), .Z1_f (new_AGEMA_signal_3968) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_0_2_U1 ( .A0_t (ShiftRowsOutput[34]), .A0_f (new_AGEMA_signal_2999), .A1_t (new_AGEMA_signal_3000), .A1_f (new_AGEMA_signal_3001), .B0_t (SubCellInst_SboxInst_6_YY[0]), .B0_f (new_AGEMA_signal_2761), .B1_t (new_AGEMA_signal_2762), .B1_f (new_AGEMA_signal_2763), .Z0_t (MCOutput[18]), .Z0_f (new_AGEMA_signal_3194), .Z1_t (new_AGEMA_signal_3195), .Z1_f (new_AGEMA_signal_3196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_0_3_U1 ( .A0_t (ShiftRowsOutput[35]), .A0_f (new_AGEMA_signal_3329), .A1_t (new_AGEMA_signal_3330), .A1_f (new_AGEMA_signal_3331), .B0_t (SubCellInst_SboxInst_6_YY[1]), .B0_f (new_AGEMA_signal_3098), .B1_t (new_AGEMA_signal_3099), .B1_f (new_AGEMA_signal_3100), .Z0_t (MCOutput[19]), .Z0_f (new_AGEMA_signal_3540), .Z1_t (new_AGEMA_signal_3541), .Z1_f (new_AGEMA_signal_3542) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_1_0_U1 ( .A0_t (ShiftRowsOutput[36]), .A0_f (new_AGEMA_signal_3696), .A1_t (new_AGEMA_signal_3697), .A1_f (new_AGEMA_signal_3698), .B0_t (ShiftRowsOutput[20]), .B0_f (new_AGEMA_signal_3474), .B1_t (new_AGEMA_signal_3475), .B1_f (new_AGEMA_signal_3476), .Z0_t (MCOutput[20]), .Z0_f (new_AGEMA_signal_3837), .Z1_t (new_AGEMA_signal_3838), .Z1_f (new_AGEMA_signal_3839) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_1_1_U1 ( .A0_t (ShiftRowsOutput[37]), .A0_f (new_AGEMA_signal_3804), .A1_t (new_AGEMA_signal_3805), .A1_f (new_AGEMA_signal_3806), .B0_t (SubCellOutput[29]), .B0_f (new_AGEMA_signal_3657), .B1_t (new_AGEMA_signal_3658), .B1_f (new_AGEMA_signal_3659), .Z0_t (MCOutput[21]), .Z0_f (new_AGEMA_signal_3969), .Z1_t (new_AGEMA_signal_3970), .Z1_f (new_AGEMA_signal_3971) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_1_2_U1 ( .A0_t (ShiftRowsOutput[38]), .A0_f (new_AGEMA_signal_3002), .A1_t (new_AGEMA_signal_3003), .A1_f (new_AGEMA_signal_3004), .B0_t (SubCellInst_SboxInst_7_YY[0]), .B0_f (new_AGEMA_signal_2770), .B1_t (new_AGEMA_signal_2771), .B1_f (new_AGEMA_signal_2772), .Z0_t (MCOutput[22]), .Z0_f (new_AGEMA_signal_3197), .Z1_t (new_AGEMA_signal_3198), .Z1_f (new_AGEMA_signal_3199) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_1_3_U1 ( .A0_t (ShiftRowsOutput[39]), .A0_f (new_AGEMA_signal_3332), .A1_t (new_AGEMA_signal_3333), .A1_f (new_AGEMA_signal_3334), .B0_t (SubCellInst_SboxInst_7_YY[1]), .B0_f (new_AGEMA_signal_3107), .B1_t (new_AGEMA_signal_3108), .B1_f (new_AGEMA_signal_3109), .Z0_t (MCOutput[23]), .Z0_f (new_AGEMA_signal_3543), .Z1_t (new_AGEMA_signal_3544), .Z1_f (new_AGEMA_signal_3545) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_2_0_U1 ( .A0_t (ShiftRowsOutput[40]), .A0_f (new_AGEMA_signal_3807), .A1_t (new_AGEMA_signal_3808), .A1_f (new_AGEMA_signal_3809), .B0_t (ShiftRowsOutput[24]), .B0_f (new_AGEMA_signal_3456), .B1_t (new_AGEMA_signal_3457), .B1_f (new_AGEMA_signal_3458), .Z0_t (MCOutput[24]), .Z0_f (new_AGEMA_signal_3972), .Z1_t (new_AGEMA_signal_3973), .Z1_f (new_AGEMA_signal_3974) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_2_1_U1 ( .A0_t (ShiftRowsOutput[41]), .A0_f (new_AGEMA_signal_3939), .A1_t (new_AGEMA_signal_3940), .A1_f (new_AGEMA_signal_3941), .B0_t (ShiftRowsOutput[25]), .B0_f (new_AGEMA_signal_3648), .B1_t (new_AGEMA_signal_3649), .B1_f (new_AGEMA_signal_3650), .Z0_t (MCOutput[25]), .Z0_f (new_AGEMA_signal_4110), .Z1_t (new_AGEMA_signal_4111), .Z1_f (new_AGEMA_signal_4112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_2_2_U1 ( .A0_t (ShiftRowsOutput[42]), .A0_f (new_AGEMA_signal_3005), .A1_t (new_AGEMA_signal_3006), .A1_f (new_AGEMA_signal_3007), .B0_t (SubCellInst_SboxInst_4_YY[0]), .B0_f (new_AGEMA_signal_2743), .B1_t (new_AGEMA_signal_2744), .B1_f (new_AGEMA_signal_2745), .Z0_t (MCOutput[26]), .Z0_f (new_AGEMA_signal_3200), .Z1_t (new_AGEMA_signal_3201), .Z1_f (new_AGEMA_signal_3202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_2_3_U1 ( .A0_t (ShiftRowsOutput[43]), .A0_f (new_AGEMA_signal_3335), .A1_t (new_AGEMA_signal_3336), .A1_f (new_AGEMA_signal_3337), .B0_t (SubCellInst_SboxInst_4_YY[1]), .B0_f (new_AGEMA_signal_3080), .B1_t (new_AGEMA_signal_3081), .B1_f (new_AGEMA_signal_3082), .Z0_t (MCOutput[27]), .Z0_f (new_AGEMA_signal_3546), .Z1_t (new_AGEMA_signal_3547), .Z1_f (new_AGEMA_signal_3548) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_3_0_U1 ( .A0_t (ShiftRowsOutput[44]), .A0_f (new_AGEMA_signal_3690), .A1_t (new_AGEMA_signal_3691), .A1_f (new_AGEMA_signal_3692), .B0_t (ShiftRowsOutput[28]), .B0_f (new_AGEMA_signal_3462), .B1_t (new_AGEMA_signal_3463), .B1_f (new_AGEMA_signal_3464), .Z0_t (MCOutput[28]), .Z0_f (new_AGEMA_signal_3840), .Z1_t (new_AGEMA_signal_3841), .Z1_f (new_AGEMA_signal_3842) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_3_1_U1 ( .A0_t (ShiftRowsOutput[45]), .A0_f (new_AGEMA_signal_3798), .A1_t (new_AGEMA_signal_3799), .A1_f (new_AGEMA_signal_3800), .B0_t (ShiftRowsOutput[29]), .B0_f (new_AGEMA_signal_3651), .B1_t (new_AGEMA_signal_3652), .B1_f (new_AGEMA_signal_3653), .Z0_t (MCOutput[29]), .Z0_f (new_AGEMA_signal_3975), .Z1_t (new_AGEMA_signal_3976), .Z1_f (new_AGEMA_signal_3977) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_3_2_U1 ( .A0_t (ShiftRowsOutput[46]), .A0_f (new_AGEMA_signal_2996), .A1_t (new_AGEMA_signal_2997), .A1_f (new_AGEMA_signal_2998), .B0_t (SubCellInst_SboxInst_5_YY[0]), .B0_f (new_AGEMA_signal_2752), .B1_t (new_AGEMA_signal_2753), .B1_f (new_AGEMA_signal_2754), .Z0_t (MCOutput[30]), .Z0_f (new_AGEMA_signal_3203), .Z1_t (new_AGEMA_signal_3204), .Z1_f (new_AGEMA_signal_3205) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_3_3_U1 ( .A0_t (ShiftRowsOutput[47]), .A0_f (new_AGEMA_signal_3326), .A1_t (new_AGEMA_signal_3327), .A1_f (new_AGEMA_signal_3328), .B0_t (SubCellInst_SboxInst_5_YY[1]), .B0_f (new_AGEMA_signal_3089), .B1_t (new_AGEMA_signal_3090), .B1_f (new_AGEMA_signal_3091), .Z0_t (MCOutput[31]), .Z0_f (new_AGEMA_signal_3549), .Z1_t (new_AGEMA_signal_3550), .Z1_f (new_AGEMA_signal_3551) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_0_0_U1 ( .A0_t (MCOutput[32]), .A0_f (new_AGEMA_signal_3699), .A1_t (new_AGEMA_signal_3700), .A1_f (new_AGEMA_signal_3701), .B0_t (ShiftRowsOutput[16]), .B0_f (new_AGEMA_signal_3468), .B1_t (new_AGEMA_signal_3469), .B1_f (new_AGEMA_signal_3470), .Z0_t (MCOutput[0]), .Z0_f (new_AGEMA_signal_3843), .Z1_t (new_AGEMA_signal_3844), .Z1_f (new_AGEMA_signal_3845) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_0_1_U1 ( .A0_t (MCOutput[33]), .A0_f (new_AGEMA_signal_3810), .A1_t (new_AGEMA_signal_3811), .A1_f (new_AGEMA_signal_3812), .B0_t (ShiftRowsOutput[17]), .B0_f (new_AGEMA_signal_3654), .B1_t (new_AGEMA_signal_3655), .B1_f (new_AGEMA_signal_3656), .Z0_t (MCOutput[1]), .Z0_f (new_AGEMA_signal_3978), .Z1_t (new_AGEMA_signal_3979), .Z1_f (new_AGEMA_signal_3980) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_0_2_U1 ( .A0_t (MCOutput[34]), .A0_f (new_AGEMA_signal_3008), .A1_t (new_AGEMA_signal_3009), .A1_f (new_AGEMA_signal_3010), .B0_t (SubCellInst_SboxInst_6_YY[0]), .B0_f (new_AGEMA_signal_2761), .B1_t (new_AGEMA_signal_2762), .B1_f (new_AGEMA_signal_2763), .Z0_t (MCOutput[2]), .Z0_f (new_AGEMA_signal_3206), .Z1_t (new_AGEMA_signal_3207), .Z1_f (new_AGEMA_signal_3208) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_0_3_U1 ( .A0_t (MCOutput[35]), .A0_f (new_AGEMA_signal_3338), .A1_t (new_AGEMA_signal_3339), .A1_f (new_AGEMA_signal_3340), .B0_t (SubCellInst_SboxInst_6_YY[1]), .B0_f (new_AGEMA_signal_3098), .B1_t (new_AGEMA_signal_3099), .B1_f (new_AGEMA_signal_3100), .Z0_t (MCOutput[3]), .Z0_f (new_AGEMA_signal_3552), .Z1_t (new_AGEMA_signal_3553), .Z1_f (new_AGEMA_signal_3554) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_1_0_U1 ( .A0_t (MCOutput[36]), .A0_f (new_AGEMA_signal_3702), .A1_t (new_AGEMA_signal_3703), .A1_f (new_AGEMA_signal_3704), .B0_t (ShiftRowsOutput[20]), .B0_f (new_AGEMA_signal_3474), .B1_t (new_AGEMA_signal_3475), .B1_f (new_AGEMA_signal_3476), .Z0_t (MCOutput[4]), .Z0_f (new_AGEMA_signal_3846), .Z1_t (new_AGEMA_signal_3847), .Z1_f (new_AGEMA_signal_3848) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_1_1_U1 ( .A0_t (MCOutput[37]), .A0_f (new_AGEMA_signal_3813), .A1_t (new_AGEMA_signal_3814), .A1_f (new_AGEMA_signal_3815), .B0_t (SubCellOutput[29]), .B0_f (new_AGEMA_signal_3657), .B1_t (new_AGEMA_signal_3658), .B1_f (new_AGEMA_signal_3659), .Z0_t (MCOutput[5]), .Z0_f (new_AGEMA_signal_3981), .Z1_t (new_AGEMA_signal_3982), .Z1_f (new_AGEMA_signal_3983) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_1_2_U1 ( .A0_t (MCOutput[38]), .A0_f (new_AGEMA_signal_3011), .A1_t (new_AGEMA_signal_3012), .A1_f (new_AGEMA_signal_3013), .B0_t (SubCellInst_SboxInst_7_YY[0]), .B0_f (new_AGEMA_signal_2770), .B1_t (new_AGEMA_signal_2771), .B1_f (new_AGEMA_signal_2772), .Z0_t (MCOutput[6]), .Z0_f (new_AGEMA_signal_3209), .Z1_t (new_AGEMA_signal_3210), .Z1_f (new_AGEMA_signal_3211) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_1_3_U1 ( .A0_t (MCOutput[39]), .A0_f (new_AGEMA_signal_3341), .A1_t (new_AGEMA_signal_3342), .A1_f (new_AGEMA_signal_3343), .B0_t (SubCellInst_SboxInst_7_YY[1]), .B0_f (new_AGEMA_signal_3107), .B1_t (new_AGEMA_signal_3108), .B1_f (new_AGEMA_signal_3109), .Z0_t (MCOutput[7]), .Z0_f (new_AGEMA_signal_3555), .Z1_t (new_AGEMA_signal_3556), .Z1_f (new_AGEMA_signal_3557) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_2_0_U1 ( .A0_t (MCOutput[40]), .A0_f (new_AGEMA_signal_3705), .A1_t (new_AGEMA_signal_3706), .A1_f (new_AGEMA_signal_3707), .B0_t (ShiftRowsOutput[24]), .B0_f (new_AGEMA_signal_3456), .B1_t (new_AGEMA_signal_3457), .B1_f (new_AGEMA_signal_3458), .Z0_t (MCOutput[8]), .Z0_f (new_AGEMA_signal_3849), .Z1_t (new_AGEMA_signal_3850), .Z1_f (new_AGEMA_signal_3851) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_2_1_U1 ( .A0_t (MCOutput[41]), .A0_f (new_AGEMA_signal_3816), .A1_t (new_AGEMA_signal_3817), .A1_f (new_AGEMA_signal_3818), .B0_t (ShiftRowsOutput[25]), .B0_f (new_AGEMA_signal_3648), .B1_t (new_AGEMA_signal_3649), .B1_f (new_AGEMA_signal_3650), .Z0_t (MCOutput[9]), .Z0_f (new_AGEMA_signal_3984), .Z1_t (new_AGEMA_signal_3985), .Z1_f (new_AGEMA_signal_3986) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_2_2_U1 ( .A0_t (MCOutput[42]), .A0_f (new_AGEMA_signal_3014), .A1_t (new_AGEMA_signal_3015), .A1_f (new_AGEMA_signal_3016), .B0_t (SubCellInst_SboxInst_4_YY[0]), .B0_f (new_AGEMA_signal_2743), .B1_t (new_AGEMA_signal_2744), .B1_f (new_AGEMA_signal_2745), .Z0_t (MCOutput[10]), .Z0_f (new_AGEMA_signal_3212), .Z1_t (new_AGEMA_signal_3213), .Z1_f (new_AGEMA_signal_3214) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_2_3_U1 ( .A0_t (MCOutput[43]), .A0_f (new_AGEMA_signal_3344), .A1_t (new_AGEMA_signal_3345), .A1_f (new_AGEMA_signal_3346), .B0_t (SubCellInst_SboxInst_4_YY[1]), .B0_f (new_AGEMA_signal_3080), .B1_t (new_AGEMA_signal_3081), .B1_f (new_AGEMA_signal_3082), .Z0_t (MCOutput[11]), .Z0_f (new_AGEMA_signal_3558), .Z1_t (new_AGEMA_signal_3559), .Z1_f (new_AGEMA_signal_3560) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_3_0_U1 ( .A0_t (MCOutput[44]), .A0_f (new_AGEMA_signal_3819), .A1_t (new_AGEMA_signal_3820), .A1_f (new_AGEMA_signal_3821), .B0_t (ShiftRowsOutput[28]), .B0_f (new_AGEMA_signal_3462), .B1_t (new_AGEMA_signal_3463), .B1_f (new_AGEMA_signal_3464), .Z0_t (MCOutput[12]), .Z0_f (new_AGEMA_signal_3987), .Z1_t (new_AGEMA_signal_3988), .Z1_f (new_AGEMA_signal_3989) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_3_1_U1 ( .A0_t (MCOutput[45]), .A0_f (new_AGEMA_signal_3942), .A1_t (new_AGEMA_signal_3943), .A1_f (new_AGEMA_signal_3944), .B0_t (ShiftRowsOutput[29]), .B0_f (new_AGEMA_signal_3651), .B1_t (new_AGEMA_signal_3652), .B1_f (new_AGEMA_signal_3653), .Z0_t (MCOutput[13]), .Z0_f (new_AGEMA_signal_4113), .Z1_t (new_AGEMA_signal_4114), .Z1_f (new_AGEMA_signal_4115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_3_2_U1 ( .A0_t (MCOutput[46]), .A0_f (new_AGEMA_signal_3182), .A1_t (new_AGEMA_signal_3183), .A1_f (new_AGEMA_signal_3184), .B0_t (SubCellInst_SboxInst_5_YY[0]), .B0_f (new_AGEMA_signal_2752), .B1_t (new_AGEMA_signal_2753), .B1_f (new_AGEMA_signal_2754), .Z0_t (MCOutput[14]), .Z0_f (new_AGEMA_signal_3359), .Z1_t (new_AGEMA_signal_3360), .Z1_f (new_AGEMA_signal_3361) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_3_3_U1 ( .A0_t (MCOutput[47]), .A0_f (new_AGEMA_signal_3525), .A1_t (new_AGEMA_signal_3526), .A1_f (new_AGEMA_signal_3527), .B0_t (SubCellInst_SboxInst_5_YY[1]), .B0_f (new_AGEMA_signal_3089), .B1_t (new_AGEMA_signal_3090), .B1_f (new_AGEMA_signal_3091), .Z0_t (MCOutput[15]), .Z0_f (new_AGEMA_signal_3720), .Z1_t (new_AGEMA_signal_3721), .Z1_f (new_AGEMA_signal_3722) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_0_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[0]), .A0_f (new_AGEMA_signal_1723), .A1_t (new_AGEMA_signal_1724), .A1_f (new_AGEMA_signal_1725), .B0_t (Key_s0_t[0]), .B0_f (Key_s0_f[0]), .B1_t (Key_s1_t[0]), .B1_f (Key_s1_f[0]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_0_U1_X), .Z0_f (new_AGEMA_signal_1729), .Z1_t (new_AGEMA_signal_1730), .Z1_f (new_AGEMA_signal_1731) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_0_U1_X), .B0_f (new_AGEMA_signal_1729), .B1_t (new_AGEMA_signal_1730), .B1_f (new_AGEMA_signal_1731), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_0_U1_Y), .Z0_f (new_AGEMA_signal_2505), .Z1_t (new_AGEMA_signal_2506), .Z1_f (new_AGEMA_signal_2507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_0_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_0_U1_Y), .A0_f (new_AGEMA_signal_2505), .A1_t (new_AGEMA_signal_2506), .A1_f (new_AGEMA_signal_2507), .B0_t (TweakeyGeneration_key_Feedback[0]), .B0_f (new_AGEMA_signal_1723), .B1_t (new_AGEMA_signal_1724), .B1_f (new_AGEMA_signal_1725), .Z0_t (TweakeyGeneration_key_Feedback[56]), .Z0_f (new_AGEMA_signal_2227), .Z1_t (new_AGEMA_signal_2228), .Z1_f (new_AGEMA_signal_2229) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_1_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[1]), .A0_f (new_AGEMA_signal_1732), .A1_t (new_AGEMA_signal_1733), .A1_f (new_AGEMA_signal_1734), .B0_t (Key_s0_t[1]), .B0_f (Key_s0_f[1]), .B1_t (Key_s1_t[1]), .B1_f (Key_s1_f[1]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_1_U1_X), .Z0_f (new_AGEMA_signal_1738), .Z1_t (new_AGEMA_signal_1739), .Z1_f (new_AGEMA_signal_1740) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_1_U1_X), .B0_f (new_AGEMA_signal_1738), .B1_t (new_AGEMA_signal_1739), .B1_f (new_AGEMA_signal_1740), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_1_U1_Y), .Z0_f (new_AGEMA_signal_2508), .Z1_t (new_AGEMA_signal_2509), .Z1_f (new_AGEMA_signal_2510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_1_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_1_U1_Y), .A0_f (new_AGEMA_signal_2508), .A1_t (new_AGEMA_signal_2509), .A1_f (new_AGEMA_signal_2510), .B0_t (TweakeyGeneration_key_Feedback[1]), .B0_f (new_AGEMA_signal_1732), .B1_t (new_AGEMA_signal_1733), .B1_f (new_AGEMA_signal_1734), .Z0_t (TweakeyGeneration_key_Feedback[57]), .Z0_f (new_AGEMA_signal_2236), .Z1_t (new_AGEMA_signal_2237), .Z1_f (new_AGEMA_signal_2238) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_2_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[2]), .A0_f (new_AGEMA_signal_1741), .A1_t (new_AGEMA_signal_1742), .A1_f (new_AGEMA_signal_1743), .B0_t (Key_s0_t[2]), .B0_f (Key_s0_f[2]), .B1_t (Key_s1_t[2]), .B1_f (Key_s1_f[2]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_2_U1_X), .Z0_f (new_AGEMA_signal_1747), .Z1_t (new_AGEMA_signal_1748), .Z1_f (new_AGEMA_signal_1749) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_2_U1_X), .B0_f (new_AGEMA_signal_1747), .B1_t (new_AGEMA_signal_1748), .B1_f (new_AGEMA_signal_1749), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_2_U1_Y), .Z0_f (new_AGEMA_signal_2511), .Z1_t (new_AGEMA_signal_2512), .Z1_f (new_AGEMA_signal_2513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_2_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_2_U1_Y), .A0_f (new_AGEMA_signal_2511), .A1_t (new_AGEMA_signal_2512), .A1_f (new_AGEMA_signal_2513), .B0_t (TweakeyGeneration_key_Feedback[2]), .B0_f (new_AGEMA_signal_1741), .B1_t (new_AGEMA_signal_1742), .B1_f (new_AGEMA_signal_1743), .Z0_t (TweakeyGeneration_key_Feedback[58]), .Z0_f (new_AGEMA_signal_2245), .Z1_t (new_AGEMA_signal_2246), .Z1_f (new_AGEMA_signal_2247) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_3_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[3]), .A0_f (new_AGEMA_signal_1750), .A1_t (new_AGEMA_signal_1751), .A1_f (new_AGEMA_signal_1752), .B0_t (Key_s0_t[3]), .B0_f (Key_s0_f[3]), .B1_t (Key_s1_t[3]), .B1_f (Key_s1_f[3]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_3_U1_X), .Z0_f (new_AGEMA_signal_1756), .Z1_t (new_AGEMA_signal_1757), .Z1_f (new_AGEMA_signal_1758) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_3_U1_X), .B0_f (new_AGEMA_signal_1756), .B1_t (new_AGEMA_signal_1757), .B1_f (new_AGEMA_signal_1758), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_3_U1_Y), .Z0_f (new_AGEMA_signal_2514), .Z1_t (new_AGEMA_signal_2515), .Z1_f (new_AGEMA_signal_2516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_3_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_3_U1_Y), .A0_f (new_AGEMA_signal_2514), .A1_t (new_AGEMA_signal_2515), .A1_f (new_AGEMA_signal_2516), .B0_t (TweakeyGeneration_key_Feedback[3]), .B0_f (new_AGEMA_signal_1750), .B1_t (new_AGEMA_signal_1751), .B1_f (new_AGEMA_signal_1752), .Z0_t (TweakeyGeneration_key_Feedback[59]), .Z0_f (new_AGEMA_signal_2254), .Z1_t (new_AGEMA_signal_2255), .Z1_f (new_AGEMA_signal_2256) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_4_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[4]), .A0_f (new_AGEMA_signal_1759), .A1_t (new_AGEMA_signal_1760), .A1_f (new_AGEMA_signal_1761), .B0_t (Key_s0_t[4]), .B0_f (Key_s0_f[4]), .B1_t (Key_s1_t[4]), .B1_f (Key_s1_f[4]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_4_U1_X), .Z0_f (new_AGEMA_signal_1765), .Z1_t (new_AGEMA_signal_1766), .Z1_f (new_AGEMA_signal_1767) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_4_U1_X), .B0_f (new_AGEMA_signal_1765), .B1_t (new_AGEMA_signal_1766), .B1_f (new_AGEMA_signal_1767), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_4_U1_Y), .Z0_f (new_AGEMA_signal_2517), .Z1_t (new_AGEMA_signal_2518), .Z1_f (new_AGEMA_signal_2519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_4_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_4_U1_Y), .A0_f (new_AGEMA_signal_2517), .A1_t (new_AGEMA_signal_2518), .A1_f (new_AGEMA_signal_2519), .B0_t (TweakeyGeneration_key_Feedback[4]), .B0_f (new_AGEMA_signal_1759), .B1_t (new_AGEMA_signal_1760), .B1_f (new_AGEMA_signal_1761), .Z0_t (TweakeyGeneration_key_Feedback[40]), .Z0_f (new_AGEMA_signal_2083), .Z1_t (new_AGEMA_signal_2084), .Z1_f (new_AGEMA_signal_2085) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_5_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[5]), .A0_f (new_AGEMA_signal_1768), .A1_t (new_AGEMA_signal_1769), .A1_f (new_AGEMA_signal_1770), .B0_t (Key_s0_t[5]), .B0_f (Key_s0_f[5]), .B1_t (Key_s1_t[5]), .B1_f (Key_s1_f[5]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_5_U1_X), .Z0_f (new_AGEMA_signal_1774), .Z1_t (new_AGEMA_signal_1775), .Z1_f (new_AGEMA_signal_1776) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_5_U1_X), .B0_f (new_AGEMA_signal_1774), .B1_t (new_AGEMA_signal_1775), .B1_f (new_AGEMA_signal_1776), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_5_U1_Y), .Z0_f (new_AGEMA_signal_2520), .Z1_t (new_AGEMA_signal_2521), .Z1_f (new_AGEMA_signal_2522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_5_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_5_U1_Y), .A0_f (new_AGEMA_signal_2520), .A1_t (new_AGEMA_signal_2521), .A1_f (new_AGEMA_signal_2522), .B0_t (TweakeyGeneration_key_Feedback[5]), .B0_f (new_AGEMA_signal_1768), .B1_t (new_AGEMA_signal_1769), .B1_f (new_AGEMA_signal_1770), .Z0_t (TweakeyGeneration_key_Feedback[41]), .Z0_f (new_AGEMA_signal_2092), .Z1_t (new_AGEMA_signal_2093), .Z1_f (new_AGEMA_signal_2094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_6_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[6]), .A0_f (new_AGEMA_signal_1777), .A1_t (new_AGEMA_signal_1778), .A1_f (new_AGEMA_signal_1779), .B0_t (Key_s0_t[6]), .B0_f (Key_s0_f[6]), .B1_t (Key_s1_t[6]), .B1_f (Key_s1_f[6]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_6_U1_X), .Z0_f (new_AGEMA_signal_1783), .Z1_t (new_AGEMA_signal_1784), .Z1_f (new_AGEMA_signal_1785) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_6_U1_X), .B0_f (new_AGEMA_signal_1783), .B1_t (new_AGEMA_signal_1784), .B1_f (new_AGEMA_signal_1785), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_6_U1_Y), .Z0_f (new_AGEMA_signal_2523), .Z1_t (new_AGEMA_signal_2524), .Z1_f (new_AGEMA_signal_2525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_6_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_6_U1_Y), .A0_f (new_AGEMA_signal_2523), .A1_t (new_AGEMA_signal_2524), .A1_f (new_AGEMA_signal_2525), .B0_t (TweakeyGeneration_key_Feedback[6]), .B0_f (new_AGEMA_signal_1777), .B1_t (new_AGEMA_signal_1778), .B1_f (new_AGEMA_signal_1779), .Z0_t (TweakeyGeneration_key_Feedback[42]), .Z0_f (new_AGEMA_signal_2101), .Z1_t (new_AGEMA_signal_2102), .Z1_f (new_AGEMA_signal_2103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_7_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[7]), .A0_f (new_AGEMA_signal_1786), .A1_t (new_AGEMA_signal_1787), .A1_f (new_AGEMA_signal_1788), .B0_t (Key_s0_t[7]), .B0_f (Key_s0_f[7]), .B1_t (Key_s1_t[7]), .B1_f (Key_s1_f[7]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_7_U1_X), .Z0_f (new_AGEMA_signal_1792), .Z1_t (new_AGEMA_signal_1793), .Z1_f (new_AGEMA_signal_1794) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_7_U1_X), .B0_f (new_AGEMA_signal_1792), .B1_t (new_AGEMA_signal_1793), .B1_f (new_AGEMA_signal_1794), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_7_U1_Y), .Z0_f (new_AGEMA_signal_2526), .Z1_t (new_AGEMA_signal_2527), .Z1_f (new_AGEMA_signal_2528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_7_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_7_U1_Y), .A0_f (new_AGEMA_signal_2526), .A1_t (new_AGEMA_signal_2527), .A1_f (new_AGEMA_signal_2528), .B0_t (TweakeyGeneration_key_Feedback[7]), .B0_f (new_AGEMA_signal_1786), .B1_t (new_AGEMA_signal_1787), .B1_f (new_AGEMA_signal_1788), .Z0_t (TweakeyGeneration_key_Feedback[43]), .Z0_f (new_AGEMA_signal_2110), .Z1_t (new_AGEMA_signal_2111), .Z1_f (new_AGEMA_signal_2112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_8_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[8]), .A0_f (new_AGEMA_signal_1795), .A1_t (new_AGEMA_signal_1796), .A1_f (new_AGEMA_signal_1797), .B0_t (Key_s0_t[8]), .B0_f (Key_s0_f[8]), .B1_t (Key_s1_t[8]), .B1_f (Key_s1_f[8]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_8_U1_X), .Z0_f (new_AGEMA_signal_1801), .Z1_t (new_AGEMA_signal_1802), .Z1_f (new_AGEMA_signal_1803) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_8_U1_X), .B0_f (new_AGEMA_signal_1801), .B1_t (new_AGEMA_signal_1802), .B1_f (new_AGEMA_signal_1803), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_8_U1_Y), .Z0_f (new_AGEMA_signal_2529), .Z1_t (new_AGEMA_signal_2530), .Z1_f (new_AGEMA_signal_2531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_8_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_8_U1_Y), .A0_f (new_AGEMA_signal_2529), .A1_t (new_AGEMA_signal_2530), .A1_f (new_AGEMA_signal_2531), .B0_t (TweakeyGeneration_key_Feedback[8]), .B0_f (new_AGEMA_signal_1795), .B1_t (new_AGEMA_signal_1796), .B1_f (new_AGEMA_signal_1797), .Z0_t (TweakeyGeneration_key_Feedback[48]), .Z0_f (new_AGEMA_signal_2155), .Z1_t (new_AGEMA_signal_2156), .Z1_f (new_AGEMA_signal_2157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_9_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[9]), .A0_f (new_AGEMA_signal_1804), .A1_t (new_AGEMA_signal_1805), .A1_f (new_AGEMA_signal_1806), .B0_t (Key_s0_t[9]), .B0_f (Key_s0_f[9]), .B1_t (Key_s1_t[9]), .B1_f (Key_s1_f[9]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_9_U1_X), .Z0_f (new_AGEMA_signal_1810), .Z1_t (new_AGEMA_signal_1811), .Z1_f (new_AGEMA_signal_1812) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_9_U1_X), .B0_f (new_AGEMA_signal_1810), .B1_t (new_AGEMA_signal_1811), .B1_f (new_AGEMA_signal_1812), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_9_U1_Y), .Z0_f (new_AGEMA_signal_2532), .Z1_t (new_AGEMA_signal_2533), .Z1_f (new_AGEMA_signal_2534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_9_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_9_U1_Y), .A0_f (new_AGEMA_signal_2532), .A1_t (new_AGEMA_signal_2533), .A1_f (new_AGEMA_signal_2534), .B0_t (TweakeyGeneration_key_Feedback[9]), .B0_f (new_AGEMA_signal_1804), .B1_t (new_AGEMA_signal_1805), .B1_f (new_AGEMA_signal_1806), .Z0_t (TweakeyGeneration_key_Feedback[49]), .Z0_f (new_AGEMA_signal_2164), .Z1_t (new_AGEMA_signal_2165), .Z1_f (new_AGEMA_signal_2166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_10_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[10]), .A0_f (new_AGEMA_signal_1813), .A1_t (new_AGEMA_signal_1814), .A1_f (new_AGEMA_signal_1815), .B0_t (Key_s0_t[10]), .B0_f (Key_s0_f[10]), .B1_t (Key_s1_t[10]), .B1_f (Key_s1_f[10]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_10_U1_X), .Z0_f (new_AGEMA_signal_1819), .Z1_t (new_AGEMA_signal_1820), .Z1_f (new_AGEMA_signal_1821) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_10_U1_X), .B0_f (new_AGEMA_signal_1819), .B1_t (new_AGEMA_signal_1820), .B1_f (new_AGEMA_signal_1821), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_10_U1_Y), .Z0_f (new_AGEMA_signal_2535), .Z1_t (new_AGEMA_signal_2536), .Z1_f (new_AGEMA_signal_2537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_10_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_10_U1_Y), .A0_f (new_AGEMA_signal_2535), .A1_t (new_AGEMA_signal_2536), .A1_f (new_AGEMA_signal_2537), .B0_t (TweakeyGeneration_key_Feedback[10]), .B0_f (new_AGEMA_signal_1813), .B1_t (new_AGEMA_signal_1814), .B1_f (new_AGEMA_signal_1815), .Z0_t (TweakeyGeneration_key_Feedback[50]), .Z0_f (new_AGEMA_signal_2173), .Z1_t (new_AGEMA_signal_2174), .Z1_f (new_AGEMA_signal_2175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_11_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[11]), .A0_f (new_AGEMA_signal_1822), .A1_t (new_AGEMA_signal_1823), .A1_f (new_AGEMA_signal_1824), .B0_t (Key_s0_t[11]), .B0_f (Key_s0_f[11]), .B1_t (Key_s1_t[11]), .B1_f (Key_s1_f[11]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_11_U1_X), .Z0_f (new_AGEMA_signal_1828), .Z1_t (new_AGEMA_signal_1829), .Z1_f (new_AGEMA_signal_1830) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_11_U1_X), .B0_f (new_AGEMA_signal_1828), .B1_t (new_AGEMA_signal_1829), .B1_f (new_AGEMA_signal_1830), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_11_U1_Y), .Z0_f (new_AGEMA_signal_2538), .Z1_t (new_AGEMA_signal_2539), .Z1_f (new_AGEMA_signal_2540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_11_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_11_U1_Y), .A0_f (new_AGEMA_signal_2538), .A1_t (new_AGEMA_signal_2539), .A1_f (new_AGEMA_signal_2540), .B0_t (TweakeyGeneration_key_Feedback[11]), .B0_f (new_AGEMA_signal_1822), .B1_t (new_AGEMA_signal_1823), .B1_f (new_AGEMA_signal_1824), .Z0_t (TweakeyGeneration_key_Feedback[51]), .Z0_f (new_AGEMA_signal_2182), .Z1_t (new_AGEMA_signal_2183), .Z1_f (new_AGEMA_signal_2184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_12_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[12]), .A0_f (new_AGEMA_signal_1831), .A1_t (new_AGEMA_signal_1832), .A1_f (new_AGEMA_signal_1833), .B0_t (Key_s0_t[12]), .B0_f (Key_s0_f[12]), .B1_t (Key_s1_t[12]), .B1_f (Key_s1_f[12]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_12_U1_X), .Z0_f (new_AGEMA_signal_1837), .Z1_t (new_AGEMA_signal_1838), .Z1_f (new_AGEMA_signal_1839) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_12_U1_X), .B0_f (new_AGEMA_signal_1837), .B1_t (new_AGEMA_signal_1838), .B1_f (new_AGEMA_signal_1839), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_12_U1_Y), .Z0_f (new_AGEMA_signal_2541), .Z1_t (new_AGEMA_signal_2542), .Z1_f (new_AGEMA_signal_2543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_12_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_12_U1_Y), .A0_f (new_AGEMA_signal_2541), .A1_t (new_AGEMA_signal_2542), .A1_f (new_AGEMA_signal_2543), .B0_t (TweakeyGeneration_key_Feedback[12]), .B0_f (new_AGEMA_signal_1831), .B1_t (new_AGEMA_signal_1832), .B1_f (new_AGEMA_signal_1833), .Z0_t (TweakeyGeneration_key_Feedback[36]), .Z0_f (new_AGEMA_signal_2047), .Z1_t (new_AGEMA_signal_2048), .Z1_f (new_AGEMA_signal_2049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_13_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[13]), .A0_f (new_AGEMA_signal_1840), .A1_t (new_AGEMA_signal_1841), .A1_f (new_AGEMA_signal_1842), .B0_t (Key_s0_t[13]), .B0_f (Key_s0_f[13]), .B1_t (Key_s1_t[13]), .B1_f (Key_s1_f[13]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_13_U1_X), .Z0_f (new_AGEMA_signal_1846), .Z1_t (new_AGEMA_signal_1847), .Z1_f (new_AGEMA_signal_1848) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_13_U1_X), .B0_f (new_AGEMA_signal_1846), .B1_t (new_AGEMA_signal_1847), .B1_f (new_AGEMA_signal_1848), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_13_U1_Y), .Z0_f (new_AGEMA_signal_2544), .Z1_t (new_AGEMA_signal_2545), .Z1_f (new_AGEMA_signal_2546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_13_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_13_U1_Y), .A0_f (new_AGEMA_signal_2544), .A1_t (new_AGEMA_signal_2545), .A1_f (new_AGEMA_signal_2546), .B0_t (TweakeyGeneration_key_Feedback[13]), .B0_f (new_AGEMA_signal_1840), .B1_t (new_AGEMA_signal_1841), .B1_f (new_AGEMA_signal_1842), .Z0_t (TweakeyGeneration_key_Feedback[37]), .Z0_f (new_AGEMA_signal_2056), .Z1_t (new_AGEMA_signal_2057), .Z1_f (new_AGEMA_signal_2058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_14_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[14]), .A0_f (new_AGEMA_signal_1849), .A1_t (new_AGEMA_signal_1850), .A1_f (new_AGEMA_signal_1851), .B0_t (Key_s0_t[14]), .B0_f (Key_s0_f[14]), .B1_t (Key_s1_t[14]), .B1_f (Key_s1_f[14]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_14_U1_X), .Z0_f (new_AGEMA_signal_1855), .Z1_t (new_AGEMA_signal_1856), .Z1_f (new_AGEMA_signal_1857) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_14_U1_X), .B0_f (new_AGEMA_signal_1855), .B1_t (new_AGEMA_signal_1856), .B1_f (new_AGEMA_signal_1857), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_14_U1_Y), .Z0_f (new_AGEMA_signal_2547), .Z1_t (new_AGEMA_signal_2548), .Z1_f (new_AGEMA_signal_2549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_14_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_14_U1_Y), .A0_f (new_AGEMA_signal_2547), .A1_t (new_AGEMA_signal_2548), .A1_f (new_AGEMA_signal_2549), .B0_t (TweakeyGeneration_key_Feedback[14]), .B0_f (new_AGEMA_signal_1849), .B1_t (new_AGEMA_signal_1850), .B1_f (new_AGEMA_signal_1851), .Z0_t (TweakeyGeneration_key_Feedback[38]), .Z0_f (new_AGEMA_signal_2065), .Z1_t (new_AGEMA_signal_2066), .Z1_f (new_AGEMA_signal_2067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_15_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[15]), .A0_f (new_AGEMA_signal_1858), .A1_t (new_AGEMA_signal_1859), .A1_f (new_AGEMA_signal_1860), .B0_t (Key_s0_t[15]), .B0_f (Key_s0_f[15]), .B1_t (Key_s1_t[15]), .B1_f (Key_s1_f[15]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_15_U1_X), .Z0_f (new_AGEMA_signal_1864), .Z1_t (new_AGEMA_signal_1865), .Z1_f (new_AGEMA_signal_1866) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_15_U1_X), .B0_f (new_AGEMA_signal_1864), .B1_t (new_AGEMA_signal_1865), .B1_f (new_AGEMA_signal_1866), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_15_U1_Y), .Z0_f (new_AGEMA_signal_2550), .Z1_t (new_AGEMA_signal_2551), .Z1_f (new_AGEMA_signal_2552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_15_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_15_U1_Y), .A0_f (new_AGEMA_signal_2550), .A1_t (new_AGEMA_signal_2551), .A1_f (new_AGEMA_signal_2552), .B0_t (TweakeyGeneration_key_Feedback[15]), .B0_f (new_AGEMA_signal_1858), .B1_t (new_AGEMA_signal_1859), .B1_f (new_AGEMA_signal_1860), .Z0_t (TweakeyGeneration_key_Feedback[39]), .Z0_f (new_AGEMA_signal_2074), .Z1_t (new_AGEMA_signal_2075), .Z1_f (new_AGEMA_signal_2076) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_16_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[16]), .A0_f (new_AGEMA_signal_1867), .A1_t (new_AGEMA_signal_1868), .A1_f (new_AGEMA_signal_1869), .B0_t (Key_s0_t[16]), .B0_f (Key_s0_f[16]), .B1_t (Key_s1_t[16]), .B1_f (Key_s1_f[16]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_16_U1_X), .Z0_f (new_AGEMA_signal_1873), .Z1_t (new_AGEMA_signal_1874), .Z1_f (new_AGEMA_signal_1875) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_16_U1_X), .B0_f (new_AGEMA_signal_1873), .B1_t (new_AGEMA_signal_1874), .B1_f (new_AGEMA_signal_1875), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_16_U1_Y), .Z0_f (new_AGEMA_signal_2553), .Z1_t (new_AGEMA_signal_2554), .Z1_f (new_AGEMA_signal_2555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_16_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_16_U1_Y), .A0_f (new_AGEMA_signal_2553), .A1_t (new_AGEMA_signal_2554), .A1_f (new_AGEMA_signal_2555), .B0_t (TweakeyGeneration_key_Feedback[16]), .B0_f (new_AGEMA_signal_1867), .B1_t (new_AGEMA_signal_1868), .B1_f (new_AGEMA_signal_1869), .Z0_t (TweakeyGeneration_key_Feedback[32]), .Z0_f (new_AGEMA_signal_2011), .Z1_t (new_AGEMA_signal_2012), .Z1_f (new_AGEMA_signal_2013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_17_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[17]), .A0_f (new_AGEMA_signal_1876), .A1_t (new_AGEMA_signal_1877), .A1_f (new_AGEMA_signal_1878), .B0_t (Key_s0_t[17]), .B0_f (Key_s0_f[17]), .B1_t (Key_s1_t[17]), .B1_f (Key_s1_f[17]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_17_U1_X), .Z0_f (new_AGEMA_signal_1882), .Z1_t (new_AGEMA_signal_1883), .Z1_f (new_AGEMA_signal_1884) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_17_U1_X), .B0_f (new_AGEMA_signal_1882), .B1_t (new_AGEMA_signal_1883), .B1_f (new_AGEMA_signal_1884), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_17_U1_Y), .Z0_f (new_AGEMA_signal_2556), .Z1_t (new_AGEMA_signal_2557), .Z1_f (new_AGEMA_signal_2558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_17_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_17_U1_Y), .A0_f (new_AGEMA_signal_2556), .A1_t (new_AGEMA_signal_2557), .A1_f (new_AGEMA_signal_2558), .B0_t (TweakeyGeneration_key_Feedback[17]), .B0_f (new_AGEMA_signal_1876), .B1_t (new_AGEMA_signal_1877), .B1_f (new_AGEMA_signal_1878), .Z0_t (TweakeyGeneration_key_Feedback[33]), .Z0_f (new_AGEMA_signal_2020), .Z1_t (new_AGEMA_signal_2021), .Z1_f (new_AGEMA_signal_2022) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_18_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[18]), .A0_f (new_AGEMA_signal_1885), .A1_t (new_AGEMA_signal_1886), .A1_f (new_AGEMA_signal_1887), .B0_t (Key_s0_t[18]), .B0_f (Key_s0_f[18]), .B1_t (Key_s1_t[18]), .B1_f (Key_s1_f[18]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_18_U1_X), .Z0_f (new_AGEMA_signal_1891), .Z1_t (new_AGEMA_signal_1892), .Z1_f (new_AGEMA_signal_1893) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_18_U1_X), .B0_f (new_AGEMA_signal_1891), .B1_t (new_AGEMA_signal_1892), .B1_f (new_AGEMA_signal_1893), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_18_U1_Y), .Z0_f (new_AGEMA_signal_2559), .Z1_t (new_AGEMA_signal_2560), .Z1_f (new_AGEMA_signal_2561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_18_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_18_U1_Y), .A0_f (new_AGEMA_signal_2559), .A1_t (new_AGEMA_signal_2560), .A1_f (new_AGEMA_signal_2561), .B0_t (TweakeyGeneration_key_Feedback[18]), .B0_f (new_AGEMA_signal_1885), .B1_t (new_AGEMA_signal_1886), .B1_f (new_AGEMA_signal_1887), .Z0_t (TweakeyGeneration_key_Feedback[34]), .Z0_f (new_AGEMA_signal_2029), .Z1_t (new_AGEMA_signal_2030), .Z1_f (new_AGEMA_signal_2031) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_19_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[19]), .A0_f (new_AGEMA_signal_1894), .A1_t (new_AGEMA_signal_1895), .A1_f (new_AGEMA_signal_1896), .B0_t (Key_s0_t[19]), .B0_f (Key_s0_f[19]), .B1_t (Key_s1_t[19]), .B1_f (Key_s1_f[19]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_19_U1_X), .Z0_f (new_AGEMA_signal_1900), .Z1_t (new_AGEMA_signal_1901), .Z1_f (new_AGEMA_signal_1902) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_19_U1_X), .B0_f (new_AGEMA_signal_1900), .B1_t (new_AGEMA_signal_1901), .B1_f (new_AGEMA_signal_1902), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_19_U1_Y), .Z0_f (new_AGEMA_signal_2562), .Z1_t (new_AGEMA_signal_2563), .Z1_f (new_AGEMA_signal_2564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_19_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_19_U1_Y), .A0_f (new_AGEMA_signal_2562), .A1_t (new_AGEMA_signal_2563), .A1_f (new_AGEMA_signal_2564), .B0_t (TweakeyGeneration_key_Feedback[19]), .B0_f (new_AGEMA_signal_1894), .B1_t (new_AGEMA_signal_1895), .B1_f (new_AGEMA_signal_1896), .Z0_t (TweakeyGeneration_key_Feedback[35]), .Z0_f (new_AGEMA_signal_2038), .Z1_t (new_AGEMA_signal_2039), .Z1_f (new_AGEMA_signal_2040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_20_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[20]), .A0_f (new_AGEMA_signal_1903), .A1_t (new_AGEMA_signal_1904), .A1_f (new_AGEMA_signal_1905), .B0_t (Key_s0_t[20]), .B0_f (Key_s0_f[20]), .B1_t (Key_s1_t[20]), .B1_f (Key_s1_f[20]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_20_U1_X), .Z0_f (new_AGEMA_signal_1909), .Z1_t (new_AGEMA_signal_1910), .Z1_f (new_AGEMA_signal_1911) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_20_U1_X), .B0_f (new_AGEMA_signal_1909), .B1_t (new_AGEMA_signal_1910), .B1_f (new_AGEMA_signal_1911), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_20_U1_Y), .Z0_f (new_AGEMA_signal_2565), .Z1_t (new_AGEMA_signal_2566), .Z1_f (new_AGEMA_signal_2567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_20_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_20_U1_Y), .A0_f (new_AGEMA_signal_2565), .A1_t (new_AGEMA_signal_2566), .A1_f (new_AGEMA_signal_2567), .B0_t (TweakeyGeneration_key_Feedback[20]), .B0_f (new_AGEMA_signal_1903), .B1_t (new_AGEMA_signal_1904), .B1_f (new_AGEMA_signal_1905), .Z0_t (TweakeyGeneration_key_Feedback[44]), .Z0_f (new_AGEMA_signal_2119), .Z1_t (new_AGEMA_signal_2120), .Z1_f (new_AGEMA_signal_2121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_21_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[21]), .A0_f (new_AGEMA_signal_1912), .A1_t (new_AGEMA_signal_1913), .A1_f (new_AGEMA_signal_1914), .B0_t (Key_s0_t[21]), .B0_f (Key_s0_f[21]), .B1_t (Key_s1_t[21]), .B1_f (Key_s1_f[21]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_21_U1_X), .Z0_f (new_AGEMA_signal_1918), .Z1_t (new_AGEMA_signal_1919), .Z1_f (new_AGEMA_signal_1920) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_21_U1_X), .B0_f (new_AGEMA_signal_1918), .B1_t (new_AGEMA_signal_1919), .B1_f (new_AGEMA_signal_1920), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_21_U1_Y), .Z0_f (new_AGEMA_signal_2568), .Z1_t (new_AGEMA_signal_2569), .Z1_f (new_AGEMA_signal_2570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_21_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_21_U1_Y), .A0_f (new_AGEMA_signal_2568), .A1_t (new_AGEMA_signal_2569), .A1_f (new_AGEMA_signal_2570), .B0_t (TweakeyGeneration_key_Feedback[21]), .B0_f (new_AGEMA_signal_1912), .B1_t (new_AGEMA_signal_1913), .B1_f (new_AGEMA_signal_1914), .Z0_t (TweakeyGeneration_key_Feedback[45]), .Z0_f (new_AGEMA_signal_2128), .Z1_t (new_AGEMA_signal_2129), .Z1_f (new_AGEMA_signal_2130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_22_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[22]), .A0_f (new_AGEMA_signal_1921), .A1_t (new_AGEMA_signal_1922), .A1_f (new_AGEMA_signal_1923), .B0_t (Key_s0_t[22]), .B0_f (Key_s0_f[22]), .B1_t (Key_s1_t[22]), .B1_f (Key_s1_f[22]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_22_U1_X), .Z0_f (new_AGEMA_signal_1927), .Z1_t (new_AGEMA_signal_1928), .Z1_f (new_AGEMA_signal_1929) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_22_U1_X), .B0_f (new_AGEMA_signal_1927), .B1_t (new_AGEMA_signal_1928), .B1_f (new_AGEMA_signal_1929), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_22_U1_Y), .Z0_f (new_AGEMA_signal_2571), .Z1_t (new_AGEMA_signal_2572), .Z1_f (new_AGEMA_signal_2573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_22_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_22_U1_Y), .A0_f (new_AGEMA_signal_2571), .A1_t (new_AGEMA_signal_2572), .A1_f (new_AGEMA_signal_2573), .B0_t (TweakeyGeneration_key_Feedback[22]), .B0_f (new_AGEMA_signal_1921), .B1_t (new_AGEMA_signal_1922), .B1_f (new_AGEMA_signal_1923), .Z0_t (TweakeyGeneration_key_Feedback[46]), .Z0_f (new_AGEMA_signal_2137), .Z1_t (new_AGEMA_signal_2138), .Z1_f (new_AGEMA_signal_2139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_23_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[23]), .A0_f (new_AGEMA_signal_1930), .A1_t (new_AGEMA_signal_1931), .A1_f (new_AGEMA_signal_1932), .B0_t (Key_s0_t[23]), .B0_f (Key_s0_f[23]), .B1_t (Key_s1_t[23]), .B1_f (Key_s1_f[23]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_23_U1_X), .Z0_f (new_AGEMA_signal_1936), .Z1_t (new_AGEMA_signal_1937), .Z1_f (new_AGEMA_signal_1938) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_23_U1_X), .B0_f (new_AGEMA_signal_1936), .B1_t (new_AGEMA_signal_1937), .B1_f (new_AGEMA_signal_1938), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_23_U1_Y), .Z0_f (new_AGEMA_signal_2574), .Z1_t (new_AGEMA_signal_2575), .Z1_f (new_AGEMA_signal_2576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_23_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_23_U1_Y), .A0_f (new_AGEMA_signal_2574), .A1_t (new_AGEMA_signal_2575), .A1_f (new_AGEMA_signal_2576), .B0_t (TweakeyGeneration_key_Feedback[23]), .B0_f (new_AGEMA_signal_1930), .B1_t (new_AGEMA_signal_1931), .B1_f (new_AGEMA_signal_1932), .Z0_t (TweakeyGeneration_key_Feedback[47]), .Z0_f (new_AGEMA_signal_2146), .Z1_t (new_AGEMA_signal_2147), .Z1_f (new_AGEMA_signal_2148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_24_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[24]), .A0_f (new_AGEMA_signal_1939), .A1_t (new_AGEMA_signal_1940), .A1_f (new_AGEMA_signal_1941), .B0_t (Key_s0_t[24]), .B0_f (Key_s0_f[24]), .B1_t (Key_s1_t[24]), .B1_f (Key_s1_f[24]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_24_U1_X), .Z0_f (new_AGEMA_signal_1945), .Z1_t (new_AGEMA_signal_1946), .Z1_f (new_AGEMA_signal_1947) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_24_U1_X), .B0_f (new_AGEMA_signal_1945), .B1_t (new_AGEMA_signal_1946), .B1_f (new_AGEMA_signal_1947), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_24_U1_Y), .Z0_f (new_AGEMA_signal_2577), .Z1_t (new_AGEMA_signal_2578), .Z1_f (new_AGEMA_signal_2579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_24_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_24_U1_Y), .A0_f (new_AGEMA_signal_2577), .A1_t (new_AGEMA_signal_2578), .A1_f (new_AGEMA_signal_2579), .B0_t (TweakeyGeneration_key_Feedback[24]), .B0_f (new_AGEMA_signal_1939), .B1_t (new_AGEMA_signal_1940), .B1_f (new_AGEMA_signal_1941), .Z0_t (TweakeyGeneration_key_Feedback[60]), .Z0_f (new_AGEMA_signal_2263), .Z1_t (new_AGEMA_signal_2264), .Z1_f (new_AGEMA_signal_2265) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_25_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[25]), .A0_f (new_AGEMA_signal_1948), .A1_t (new_AGEMA_signal_1949), .A1_f (new_AGEMA_signal_1950), .B0_t (Key_s0_t[25]), .B0_f (Key_s0_f[25]), .B1_t (Key_s1_t[25]), .B1_f (Key_s1_f[25]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_25_U1_X), .Z0_f (new_AGEMA_signal_1954), .Z1_t (new_AGEMA_signal_1955), .Z1_f (new_AGEMA_signal_1956) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_25_U1_X), .B0_f (new_AGEMA_signal_1954), .B1_t (new_AGEMA_signal_1955), .B1_f (new_AGEMA_signal_1956), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_25_U1_Y), .Z0_f (new_AGEMA_signal_2580), .Z1_t (new_AGEMA_signal_2581), .Z1_f (new_AGEMA_signal_2582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_25_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_25_U1_Y), .A0_f (new_AGEMA_signal_2580), .A1_t (new_AGEMA_signal_2581), .A1_f (new_AGEMA_signal_2582), .B0_t (TweakeyGeneration_key_Feedback[25]), .B0_f (new_AGEMA_signal_1948), .B1_t (new_AGEMA_signal_1949), .B1_f (new_AGEMA_signal_1950), .Z0_t (TweakeyGeneration_key_Feedback[61]), .Z0_f (new_AGEMA_signal_2272), .Z1_t (new_AGEMA_signal_2273), .Z1_f (new_AGEMA_signal_2274) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_26_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[26]), .A0_f (new_AGEMA_signal_1957), .A1_t (new_AGEMA_signal_1958), .A1_f (new_AGEMA_signal_1959), .B0_t (Key_s0_t[26]), .B0_f (Key_s0_f[26]), .B1_t (Key_s1_t[26]), .B1_f (Key_s1_f[26]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_26_U1_X), .Z0_f (new_AGEMA_signal_1963), .Z1_t (new_AGEMA_signal_1964), .Z1_f (new_AGEMA_signal_1965) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_26_U1_X), .B0_f (new_AGEMA_signal_1963), .B1_t (new_AGEMA_signal_1964), .B1_f (new_AGEMA_signal_1965), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_26_U1_Y), .Z0_f (new_AGEMA_signal_2583), .Z1_t (new_AGEMA_signal_2584), .Z1_f (new_AGEMA_signal_2585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_26_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_26_U1_Y), .A0_f (new_AGEMA_signal_2583), .A1_t (new_AGEMA_signal_2584), .A1_f (new_AGEMA_signal_2585), .B0_t (TweakeyGeneration_key_Feedback[26]), .B0_f (new_AGEMA_signal_1957), .B1_t (new_AGEMA_signal_1958), .B1_f (new_AGEMA_signal_1959), .Z0_t (TweakeyGeneration_key_Feedback[62]), .Z0_f (new_AGEMA_signal_2281), .Z1_t (new_AGEMA_signal_2282), .Z1_f (new_AGEMA_signal_2283) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_27_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[27]), .A0_f (new_AGEMA_signal_1966), .A1_t (new_AGEMA_signal_1967), .A1_f (new_AGEMA_signal_1968), .B0_t (Key_s0_t[27]), .B0_f (Key_s0_f[27]), .B1_t (Key_s1_t[27]), .B1_f (Key_s1_f[27]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_27_U1_X), .Z0_f (new_AGEMA_signal_1972), .Z1_t (new_AGEMA_signal_1973), .Z1_f (new_AGEMA_signal_1974) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_27_U1_X), .B0_f (new_AGEMA_signal_1972), .B1_t (new_AGEMA_signal_1973), .B1_f (new_AGEMA_signal_1974), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_27_U1_Y), .Z0_f (new_AGEMA_signal_2586), .Z1_t (new_AGEMA_signal_2587), .Z1_f (new_AGEMA_signal_2588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_27_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_27_U1_Y), .A0_f (new_AGEMA_signal_2586), .A1_t (new_AGEMA_signal_2587), .A1_f (new_AGEMA_signal_2588), .B0_t (TweakeyGeneration_key_Feedback[27]), .B0_f (new_AGEMA_signal_1966), .B1_t (new_AGEMA_signal_1967), .B1_f (new_AGEMA_signal_1968), .Z0_t (TweakeyGeneration_key_Feedback[63]), .Z0_f (new_AGEMA_signal_2290), .Z1_t (new_AGEMA_signal_2291), .Z1_f (new_AGEMA_signal_2292) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_28_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[28]), .A0_f (new_AGEMA_signal_1975), .A1_t (new_AGEMA_signal_1976), .A1_f (new_AGEMA_signal_1977), .B0_t (Key_s0_t[28]), .B0_f (Key_s0_f[28]), .B1_t (Key_s1_t[28]), .B1_f (Key_s1_f[28]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_28_U1_X), .Z0_f (new_AGEMA_signal_1981), .Z1_t (new_AGEMA_signal_1982), .Z1_f (new_AGEMA_signal_1983) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_28_U1_X), .B0_f (new_AGEMA_signal_1981), .B1_t (new_AGEMA_signal_1982), .B1_f (new_AGEMA_signal_1983), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_28_U1_Y), .Z0_f (new_AGEMA_signal_2589), .Z1_t (new_AGEMA_signal_2590), .Z1_f (new_AGEMA_signal_2591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_28_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_28_U1_Y), .A0_f (new_AGEMA_signal_2589), .A1_t (new_AGEMA_signal_2590), .A1_f (new_AGEMA_signal_2591), .B0_t (TweakeyGeneration_key_Feedback[28]), .B0_f (new_AGEMA_signal_1975), .B1_t (new_AGEMA_signal_1976), .B1_f (new_AGEMA_signal_1977), .Z0_t (TweakeyGeneration_key_Feedback[52]), .Z0_f (new_AGEMA_signal_2191), .Z1_t (new_AGEMA_signal_2192), .Z1_f (new_AGEMA_signal_2193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_29_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[29]), .A0_f (new_AGEMA_signal_1984), .A1_t (new_AGEMA_signal_1985), .A1_f (new_AGEMA_signal_1986), .B0_t (Key_s0_t[29]), .B0_f (Key_s0_f[29]), .B1_t (Key_s1_t[29]), .B1_f (Key_s1_f[29]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_29_U1_X), .Z0_f (new_AGEMA_signal_1990), .Z1_t (new_AGEMA_signal_1991), .Z1_f (new_AGEMA_signal_1992) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_29_U1_X), .B0_f (new_AGEMA_signal_1990), .B1_t (new_AGEMA_signal_1991), .B1_f (new_AGEMA_signal_1992), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_29_U1_Y), .Z0_f (new_AGEMA_signal_2592), .Z1_t (new_AGEMA_signal_2593), .Z1_f (new_AGEMA_signal_2594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_29_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_29_U1_Y), .A0_f (new_AGEMA_signal_2592), .A1_t (new_AGEMA_signal_2593), .A1_f (new_AGEMA_signal_2594), .B0_t (TweakeyGeneration_key_Feedback[29]), .B0_f (new_AGEMA_signal_1984), .B1_t (new_AGEMA_signal_1985), .B1_f (new_AGEMA_signal_1986), .Z0_t (TweakeyGeneration_key_Feedback[53]), .Z0_f (new_AGEMA_signal_2200), .Z1_t (new_AGEMA_signal_2201), .Z1_f (new_AGEMA_signal_2202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_30_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[30]), .A0_f (new_AGEMA_signal_1993), .A1_t (new_AGEMA_signal_1994), .A1_f (new_AGEMA_signal_1995), .B0_t (Key_s0_t[30]), .B0_f (Key_s0_f[30]), .B1_t (Key_s1_t[30]), .B1_f (Key_s1_f[30]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_30_U1_X), .Z0_f (new_AGEMA_signal_1999), .Z1_t (new_AGEMA_signal_2000), .Z1_f (new_AGEMA_signal_2001) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_30_U1_X), .B0_f (new_AGEMA_signal_1999), .B1_t (new_AGEMA_signal_2000), .B1_f (new_AGEMA_signal_2001), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_30_U1_Y), .Z0_f (new_AGEMA_signal_2595), .Z1_t (new_AGEMA_signal_2596), .Z1_f (new_AGEMA_signal_2597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_30_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_30_U1_Y), .A0_f (new_AGEMA_signal_2595), .A1_t (new_AGEMA_signal_2596), .A1_f (new_AGEMA_signal_2597), .B0_t (TweakeyGeneration_key_Feedback[30]), .B0_f (new_AGEMA_signal_1993), .B1_t (new_AGEMA_signal_1994), .B1_f (new_AGEMA_signal_1995), .Z0_t (TweakeyGeneration_key_Feedback[54]), .Z0_f (new_AGEMA_signal_2209), .Z1_t (new_AGEMA_signal_2210), .Z1_f (new_AGEMA_signal_2211) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_31_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[31]), .A0_f (new_AGEMA_signal_2002), .A1_t (new_AGEMA_signal_2003), .A1_f (new_AGEMA_signal_2004), .B0_t (Key_s0_t[31]), .B0_f (Key_s0_f[31]), .B1_t (Key_s1_t[31]), .B1_f (Key_s1_f[31]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_31_U1_X), .Z0_f (new_AGEMA_signal_2008), .Z1_t (new_AGEMA_signal_2009), .Z1_f (new_AGEMA_signal_2010) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_31_U1_X), .B0_f (new_AGEMA_signal_2008), .B1_t (new_AGEMA_signal_2009), .B1_f (new_AGEMA_signal_2010), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_31_U1_Y), .Z0_f (new_AGEMA_signal_2598), .Z1_t (new_AGEMA_signal_2599), .Z1_f (new_AGEMA_signal_2600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_31_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_31_U1_Y), .A0_f (new_AGEMA_signal_2598), .A1_t (new_AGEMA_signal_2599), .A1_f (new_AGEMA_signal_2600), .B0_t (TweakeyGeneration_key_Feedback[31]), .B0_f (new_AGEMA_signal_2002), .B1_t (new_AGEMA_signal_2003), .B1_f (new_AGEMA_signal_2004), .Z0_t (TweakeyGeneration_key_Feedback[55]), .Z0_f (new_AGEMA_signal_2218), .Z1_t (new_AGEMA_signal_2219), .Z1_f (new_AGEMA_signal_2220) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_32_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[32]), .A0_f (new_AGEMA_signal_2011), .A1_t (new_AGEMA_signal_2012), .A1_f (new_AGEMA_signal_2013), .B0_t (Key_s0_t[32]), .B0_f (Key_s0_f[32]), .B1_t (Key_s1_t[32]), .B1_f (Key_s1_f[32]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_32_U1_X), .Z0_f (new_AGEMA_signal_2017), .Z1_t (new_AGEMA_signal_2018), .Z1_f (new_AGEMA_signal_2019) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_32_U1_X), .B0_f (new_AGEMA_signal_2017), .B1_t (new_AGEMA_signal_2018), .B1_f (new_AGEMA_signal_2019), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_32_U1_Y), .Z0_f (new_AGEMA_signal_2601), .Z1_t (new_AGEMA_signal_2602), .Z1_f (new_AGEMA_signal_2603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_32_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_32_U1_Y), .A0_f (new_AGEMA_signal_2601), .A1_t (new_AGEMA_signal_2602), .A1_f (new_AGEMA_signal_2603), .B0_t (TweakeyGeneration_key_Feedback[32]), .B0_f (new_AGEMA_signal_2011), .B1_t (new_AGEMA_signal_2012), .B1_f (new_AGEMA_signal_2013), .Z0_t (TweakeyGeneration_key_Feedback[0]), .Z0_f (new_AGEMA_signal_1723), .Z1_t (new_AGEMA_signal_1724), .Z1_f (new_AGEMA_signal_1725) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_33_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[33]), .A0_f (new_AGEMA_signal_2020), .A1_t (new_AGEMA_signal_2021), .A1_f (new_AGEMA_signal_2022), .B0_t (Key_s0_t[33]), .B0_f (Key_s0_f[33]), .B1_t (Key_s1_t[33]), .B1_f (Key_s1_f[33]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_33_U1_X), .Z0_f (new_AGEMA_signal_2026), .Z1_t (new_AGEMA_signal_2027), .Z1_f (new_AGEMA_signal_2028) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_33_U1_X), .B0_f (new_AGEMA_signal_2026), .B1_t (new_AGEMA_signal_2027), .B1_f (new_AGEMA_signal_2028), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_33_U1_Y), .Z0_f (new_AGEMA_signal_2604), .Z1_t (new_AGEMA_signal_2605), .Z1_f (new_AGEMA_signal_2606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_33_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_33_U1_Y), .A0_f (new_AGEMA_signal_2604), .A1_t (new_AGEMA_signal_2605), .A1_f (new_AGEMA_signal_2606), .B0_t (TweakeyGeneration_key_Feedback[33]), .B0_f (new_AGEMA_signal_2020), .B1_t (new_AGEMA_signal_2021), .B1_f (new_AGEMA_signal_2022), .Z0_t (TweakeyGeneration_key_Feedback[1]), .Z0_f (new_AGEMA_signal_1732), .Z1_t (new_AGEMA_signal_1733), .Z1_f (new_AGEMA_signal_1734) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_34_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[34]), .A0_f (new_AGEMA_signal_2029), .A1_t (new_AGEMA_signal_2030), .A1_f (new_AGEMA_signal_2031), .B0_t (Key_s0_t[34]), .B0_f (Key_s0_f[34]), .B1_t (Key_s1_t[34]), .B1_f (Key_s1_f[34]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_34_U1_X), .Z0_f (new_AGEMA_signal_2035), .Z1_t (new_AGEMA_signal_2036), .Z1_f (new_AGEMA_signal_2037) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_34_U1_X), .B0_f (new_AGEMA_signal_2035), .B1_t (new_AGEMA_signal_2036), .B1_f (new_AGEMA_signal_2037), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_34_U1_Y), .Z0_f (new_AGEMA_signal_2607), .Z1_t (new_AGEMA_signal_2608), .Z1_f (new_AGEMA_signal_2609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_34_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_34_U1_Y), .A0_f (new_AGEMA_signal_2607), .A1_t (new_AGEMA_signal_2608), .A1_f (new_AGEMA_signal_2609), .B0_t (TweakeyGeneration_key_Feedback[34]), .B0_f (new_AGEMA_signal_2029), .B1_t (new_AGEMA_signal_2030), .B1_f (new_AGEMA_signal_2031), .Z0_t (TweakeyGeneration_key_Feedback[2]), .Z0_f (new_AGEMA_signal_1741), .Z1_t (new_AGEMA_signal_1742), .Z1_f (new_AGEMA_signal_1743) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_35_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[35]), .A0_f (new_AGEMA_signal_2038), .A1_t (new_AGEMA_signal_2039), .A1_f (new_AGEMA_signal_2040), .B0_t (Key_s0_t[35]), .B0_f (Key_s0_f[35]), .B1_t (Key_s1_t[35]), .B1_f (Key_s1_f[35]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_35_U1_X), .Z0_f (new_AGEMA_signal_2044), .Z1_t (new_AGEMA_signal_2045), .Z1_f (new_AGEMA_signal_2046) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_35_U1_X), .B0_f (new_AGEMA_signal_2044), .B1_t (new_AGEMA_signal_2045), .B1_f (new_AGEMA_signal_2046), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_35_U1_Y), .Z0_f (new_AGEMA_signal_2610), .Z1_t (new_AGEMA_signal_2611), .Z1_f (new_AGEMA_signal_2612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_35_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_35_U1_Y), .A0_f (new_AGEMA_signal_2610), .A1_t (new_AGEMA_signal_2611), .A1_f (new_AGEMA_signal_2612), .B0_t (TweakeyGeneration_key_Feedback[35]), .B0_f (new_AGEMA_signal_2038), .B1_t (new_AGEMA_signal_2039), .B1_f (new_AGEMA_signal_2040), .Z0_t (TweakeyGeneration_key_Feedback[3]), .Z0_f (new_AGEMA_signal_1750), .Z1_t (new_AGEMA_signal_1751), .Z1_f (new_AGEMA_signal_1752) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_36_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[36]), .A0_f (new_AGEMA_signal_2047), .A1_t (new_AGEMA_signal_2048), .A1_f (new_AGEMA_signal_2049), .B0_t (Key_s0_t[36]), .B0_f (Key_s0_f[36]), .B1_t (Key_s1_t[36]), .B1_f (Key_s1_f[36]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_36_U1_X), .Z0_f (new_AGEMA_signal_2053), .Z1_t (new_AGEMA_signal_2054), .Z1_f (new_AGEMA_signal_2055) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_36_U1_X), .B0_f (new_AGEMA_signal_2053), .B1_t (new_AGEMA_signal_2054), .B1_f (new_AGEMA_signal_2055), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_36_U1_Y), .Z0_f (new_AGEMA_signal_2613), .Z1_t (new_AGEMA_signal_2614), .Z1_f (new_AGEMA_signal_2615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_36_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_36_U1_Y), .A0_f (new_AGEMA_signal_2613), .A1_t (new_AGEMA_signal_2614), .A1_f (new_AGEMA_signal_2615), .B0_t (TweakeyGeneration_key_Feedback[36]), .B0_f (new_AGEMA_signal_2047), .B1_t (new_AGEMA_signal_2048), .B1_f (new_AGEMA_signal_2049), .Z0_t (TweakeyGeneration_key_Feedback[4]), .Z0_f (new_AGEMA_signal_1759), .Z1_t (new_AGEMA_signal_1760), .Z1_f (new_AGEMA_signal_1761) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_37_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[37]), .A0_f (new_AGEMA_signal_2056), .A1_t (new_AGEMA_signal_2057), .A1_f (new_AGEMA_signal_2058), .B0_t (Key_s0_t[37]), .B0_f (Key_s0_f[37]), .B1_t (Key_s1_t[37]), .B1_f (Key_s1_f[37]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_37_U1_X), .Z0_f (new_AGEMA_signal_2062), .Z1_t (new_AGEMA_signal_2063), .Z1_f (new_AGEMA_signal_2064) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_37_U1_X), .B0_f (new_AGEMA_signal_2062), .B1_t (new_AGEMA_signal_2063), .B1_f (new_AGEMA_signal_2064), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_37_U1_Y), .Z0_f (new_AGEMA_signal_2616), .Z1_t (new_AGEMA_signal_2617), .Z1_f (new_AGEMA_signal_2618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_37_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_37_U1_Y), .A0_f (new_AGEMA_signal_2616), .A1_t (new_AGEMA_signal_2617), .A1_f (new_AGEMA_signal_2618), .B0_t (TweakeyGeneration_key_Feedback[37]), .B0_f (new_AGEMA_signal_2056), .B1_t (new_AGEMA_signal_2057), .B1_f (new_AGEMA_signal_2058), .Z0_t (TweakeyGeneration_key_Feedback[5]), .Z0_f (new_AGEMA_signal_1768), .Z1_t (new_AGEMA_signal_1769), .Z1_f (new_AGEMA_signal_1770) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_38_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[38]), .A0_f (new_AGEMA_signal_2065), .A1_t (new_AGEMA_signal_2066), .A1_f (new_AGEMA_signal_2067), .B0_t (Key_s0_t[38]), .B0_f (Key_s0_f[38]), .B1_t (Key_s1_t[38]), .B1_f (Key_s1_f[38]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_38_U1_X), .Z0_f (new_AGEMA_signal_2071), .Z1_t (new_AGEMA_signal_2072), .Z1_f (new_AGEMA_signal_2073) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_38_U1_X), .B0_f (new_AGEMA_signal_2071), .B1_t (new_AGEMA_signal_2072), .B1_f (new_AGEMA_signal_2073), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_38_U1_Y), .Z0_f (new_AGEMA_signal_2619), .Z1_t (new_AGEMA_signal_2620), .Z1_f (new_AGEMA_signal_2621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_38_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_38_U1_Y), .A0_f (new_AGEMA_signal_2619), .A1_t (new_AGEMA_signal_2620), .A1_f (new_AGEMA_signal_2621), .B0_t (TweakeyGeneration_key_Feedback[38]), .B0_f (new_AGEMA_signal_2065), .B1_t (new_AGEMA_signal_2066), .B1_f (new_AGEMA_signal_2067), .Z0_t (TweakeyGeneration_key_Feedback[6]), .Z0_f (new_AGEMA_signal_1777), .Z1_t (new_AGEMA_signal_1778), .Z1_f (new_AGEMA_signal_1779) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_39_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[39]), .A0_f (new_AGEMA_signal_2074), .A1_t (new_AGEMA_signal_2075), .A1_f (new_AGEMA_signal_2076), .B0_t (Key_s0_t[39]), .B0_f (Key_s0_f[39]), .B1_t (Key_s1_t[39]), .B1_f (Key_s1_f[39]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_39_U1_X), .Z0_f (new_AGEMA_signal_2080), .Z1_t (new_AGEMA_signal_2081), .Z1_f (new_AGEMA_signal_2082) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_39_U1_X), .B0_f (new_AGEMA_signal_2080), .B1_t (new_AGEMA_signal_2081), .B1_f (new_AGEMA_signal_2082), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_39_U1_Y), .Z0_f (new_AGEMA_signal_2622), .Z1_t (new_AGEMA_signal_2623), .Z1_f (new_AGEMA_signal_2624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_39_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_39_U1_Y), .A0_f (new_AGEMA_signal_2622), .A1_t (new_AGEMA_signal_2623), .A1_f (new_AGEMA_signal_2624), .B0_t (TweakeyGeneration_key_Feedback[39]), .B0_f (new_AGEMA_signal_2074), .B1_t (new_AGEMA_signal_2075), .B1_f (new_AGEMA_signal_2076), .Z0_t (TweakeyGeneration_key_Feedback[7]), .Z0_f (new_AGEMA_signal_1786), .Z1_t (new_AGEMA_signal_1787), .Z1_f (new_AGEMA_signal_1788) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_40_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[40]), .A0_f (new_AGEMA_signal_2083), .A1_t (new_AGEMA_signal_2084), .A1_f (new_AGEMA_signal_2085), .B0_t (Key_s0_t[40]), .B0_f (Key_s0_f[40]), .B1_t (Key_s1_t[40]), .B1_f (Key_s1_f[40]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_40_U1_X), .Z0_f (new_AGEMA_signal_2089), .Z1_t (new_AGEMA_signal_2090), .Z1_f (new_AGEMA_signal_2091) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_40_U1_X), .B0_f (new_AGEMA_signal_2089), .B1_t (new_AGEMA_signal_2090), .B1_f (new_AGEMA_signal_2091), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_40_U1_Y), .Z0_f (new_AGEMA_signal_2625), .Z1_t (new_AGEMA_signal_2626), .Z1_f (new_AGEMA_signal_2627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_40_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_40_U1_Y), .A0_f (new_AGEMA_signal_2625), .A1_t (new_AGEMA_signal_2626), .A1_f (new_AGEMA_signal_2627), .B0_t (TweakeyGeneration_key_Feedback[40]), .B0_f (new_AGEMA_signal_2083), .B1_t (new_AGEMA_signal_2084), .B1_f (new_AGEMA_signal_2085), .Z0_t (TweakeyGeneration_key_Feedback[8]), .Z0_f (new_AGEMA_signal_1795), .Z1_t (new_AGEMA_signal_1796), .Z1_f (new_AGEMA_signal_1797) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_41_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[41]), .A0_f (new_AGEMA_signal_2092), .A1_t (new_AGEMA_signal_2093), .A1_f (new_AGEMA_signal_2094), .B0_t (Key_s0_t[41]), .B0_f (Key_s0_f[41]), .B1_t (Key_s1_t[41]), .B1_f (Key_s1_f[41]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_41_U1_X), .Z0_f (new_AGEMA_signal_2098), .Z1_t (new_AGEMA_signal_2099), .Z1_f (new_AGEMA_signal_2100) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_41_U1_X), .B0_f (new_AGEMA_signal_2098), .B1_t (new_AGEMA_signal_2099), .B1_f (new_AGEMA_signal_2100), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_41_U1_Y), .Z0_f (new_AGEMA_signal_2628), .Z1_t (new_AGEMA_signal_2629), .Z1_f (new_AGEMA_signal_2630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_41_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_41_U1_Y), .A0_f (new_AGEMA_signal_2628), .A1_t (new_AGEMA_signal_2629), .A1_f (new_AGEMA_signal_2630), .B0_t (TweakeyGeneration_key_Feedback[41]), .B0_f (new_AGEMA_signal_2092), .B1_t (new_AGEMA_signal_2093), .B1_f (new_AGEMA_signal_2094), .Z0_t (TweakeyGeneration_key_Feedback[9]), .Z0_f (new_AGEMA_signal_1804), .Z1_t (new_AGEMA_signal_1805), .Z1_f (new_AGEMA_signal_1806) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_42_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[42]), .A0_f (new_AGEMA_signal_2101), .A1_t (new_AGEMA_signal_2102), .A1_f (new_AGEMA_signal_2103), .B0_t (Key_s0_t[42]), .B0_f (Key_s0_f[42]), .B1_t (Key_s1_t[42]), .B1_f (Key_s1_f[42]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_42_U1_X), .Z0_f (new_AGEMA_signal_2107), .Z1_t (new_AGEMA_signal_2108), .Z1_f (new_AGEMA_signal_2109) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_42_U1_X), .B0_f (new_AGEMA_signal_2107), .B1_t (new_AGEMA_signal_2108), .B1_f (new_AGEMA_signal_2109), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_42_U1_Y), .Z0_f (new_AGEMA_signal_2631), .Z1_t (new_AGEMA_signal_2632), .Z1_f (new_AGEMA_signal_2633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_42_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_42_U1_Y), .A0_f (new_AGEMA_signal_2631), .A1_t (new_AGEMA_signal_2632), .A1_f (new_AGEMA_signal_2633), .B0_t (TweakeyGeneration_key_Feedback[42]), .B0_f (new_AGEMA_signal_2101), .B1_t (new_AGEMA_signal_2102), .B1_f (new_AGEMA_signal_2103), .Z0_t (TweakeyGeneration_key_Feedback[10]), .Z0_f (new_AGEMA_signal_1813), .Z1_t (new_AGEMA_signal_1814), .Z1_f (new_AGEMA_signal_1815) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_43_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[43]), .A0_f (new_AGEMA_signal_2110), .A1_t (new_AGEMA_signal_2111), .A1_f (new_AGEMA_signal_2112), .B0_t (Key_s0_t[43]), .B0_f (Key_s0_f[43]), .B1_t (Key_s1_t[43]), .B1_f (Key_s1_f[43]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_43_U1_X), .Z0_f (new_AGEMA_signal_2116), .Z1_t (new_AGEMA_signal_2117), .Z1_f (new_AGEMA_signal_2118) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_43_U1_X), .B0_f (new_AGEMA_signal_2116), .B1_t (new_AGEMA_signal_2117), .B1_f (new_AGEMA_signal_2118), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_43_U1_Y), .Z0_f (new_AGEMA_signal_2634), .Z1_t (new_AGEMA_signal_2635), .Z1_f (new_AGEMA_signal_2636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_43_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_43_U1_Y), .A0_f (new_AGEMA_signal_2634), .A1_t (new_AGEMA_signal_2635), .A1_f (new_AGEMA_signal_2636), .B0_t (TweakeyGeneration_key_Feedback[43]), .B0_f (new_AGEMA_signal_2110), .B1_t (new_AGEMA_signal_2111), .B1_f (new_AGEMA_signal_2112), .Z0_t (TweakeyGeneration_key_Feedback[11]), .Z0_f (new_AGEMA_signal_1822), .Z1_t (new_AGEMA_signal_1823), .Z1_f (new_AGEMA_signal_1824) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_44_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[44]), .A0_f (new_AGEMA_signal_2119), .A1_t (new_AGEMA_signal_2120), .A1_f (new_AGEMA_signal_2121), .B0_t (Key_s0_t[44]), .B0_f (Key_s0_f[44]), .B1_t (Key_s1_t[44]), .B1_f (Key_s1_f[44]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_44_U1_X), .Z0_f (new_AGEMA_signal_2125), .Z1_t (new_AGEMA_signal_2126), .Z1_f (new_AGEMA_signal_2127) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_44_U1_X), .B0_f (new_AGEMA_signal_2125), .B1_t (new_AGEMA_signal_2126), .B1_f (new_AGEMA_signal_2127), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_44_U1_Y), .Z0_f (new_AGEMA_signal_2637), .Z1_t (new_AGEMA_signal_2638), .Z1_f (new_AGEMA_signal_2639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_44_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_44_U1_Y), .A0_f (new_AGEMA_signal_2637), .A1_t (new_AGEMA_signal_2638), .A1_f (new_AGEMA_signal_2639), .B0_t (TweakeyGeneration_key_Feedback[44]), .B0_f (new_AGEMA_signal_2119), .B1_t (new_AGEMA_signal_2120), .B1_f (new_AGEMA_signal_2121), .Z0_t (TweakeyGeneration_key_Feedback[12]), .Z0_f (new_AGEMA_signal_1831), .Z1_t (new_AGEMA_signal_1832), .Z1_f (new_AGEMA_signal_1833) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_45_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[45]), .A0_f (new_AGEMA_signal_2128), .A1_t (new_AGEMA_signal_2129), .A1_f (new_AGEMA_signal_2130), .B0_t (Key_s0_t[45]), .B0_f (Key_s0_f[45]), .B1_t (Key_s1_t[45]), .B1_f (Key_s1_f[45]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_45_U1_X), .Z0_f (new_AGEMA_signal_2134), .Z1_t (new_AGEMA_signal_2135), .Z1_f (new_AGEMA_signal_2136) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_45_U1_X), .B0_f (new_AGEMA_signal_2134), .B1_t (new_AGEMA_signal_2135), .B1_f (new_AGEMA_signal_2136), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_45_U1_Y), .Z0_f (new_AGEMA_signal_2640), .Z1_t (new_AGEMA_signal_2641), .Z1_f (new_AGEMA_signal_2642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_45_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_45_U1_Y), .A0_f (new_AGEMA_signal_2640), .A1_t (new_AGEMA_signal_2641), .A1_f (new_AGEMA_signal_2642), .B0_t (TweakeyGeneration_key_Feedback[45]), .B0_f (new_AGEMA_signal_2128), .B1_t (new_AGEMA_signal_2129), .B1_f (new_AGEMA_signal_2130), .Z0_t (TweakeyGeneration_key_Feedback[13]), .Z0_f (new_AGEMA_signal_1840), .Z1_t (new_AGEMA_signal_1841), .Z1_f (new_AGEMA_signal_1842) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_46_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[46]), .A0_f (new_AGEMA_signal_2137), .A1_t (new_AGEMA_signal_2138), .A1_f (new_AGEMA_signal_2139), .B0_t (Key_s0_t[46]), .B0_f (Key_s0_f[46]), .B1_t (Key_s1_t[46]), .B1_f (Key_s1_f[46]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_46_U1_X), .Z0_f (new_AGEMA_signal_2143), .Z1_t (new_AGEMA_signal_2144), .Z1_f (new_AGEMA_signal_2145) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_46_U1_X), .B0_f (new_AGEMA_signal_2143), .B1_t (new_AGEMA_signal_2144), .B1_f (new_AGEMA_signal_2145), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_46_U1_Y), .Z0_f (new_AGEMA_signal_2643), .Z1_t (new_AGEMA_signal_2644), .Z1_f (new_AGEMA_signal_2645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_46_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_46_U1_Y), .A0_f (new_AGEMA_signal_2643), .A1_t (new_AGEMA_signal_2644), .A1_f (new_AGEMA_signal_2645), .B0_t (TweakeyGeneration_key_Feedback[46]), .B0_f (new_AGEMA_signal_2137), .B1_t (new_AGEMA_signal_2138), .B1_f (new_AGEMA_signal_2139), .Z0_t (TweakeyGeneration_key_Feedback[14]), .Z0_f (new_AGEMA_signal_1849), .Z1_t (new_AGEMA_signal_1850), .Z1_f (new_AGEMA_signal_1851) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_47_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[47]), .A0_f (new_AGEMA_signal_2146), .A1_t (new_AGEMA_signal_2147), .A1_f (new_AGEMA_signal_2148), .B0_t (Key_s0_t[47]), .B0_f (Key_s0_f[47]), .B1_t (Key_s1_t[47]), .B1_f (Key_s1_f[47]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_47_U1_X), .Z0_f (new_AGEMA_signal_2152), .Z1_t (new_AGEMA_signal_2153), .Z1_f (new_AGEMA_signal_2154) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_47_U1_X), .B0_f (new_AGEMA_signal_2152), .B1_t (new_AGEMA_signal_2153), .B1_f (new_AGEMA_signal_2154), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_47_U1_Y), .Z0_f (new_AGEMA_signal_2646), .Z1_t (new_AGEMA_signal_2647), .Z1_f (new_AGEMA_signal_2648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_47_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_47_U1_Y), .A0_f (new_AGEMA_signal_2646), .A1_t (new_AGEMA_signal_2647), .A1_f (new_AGEMA_signal_2648), .B0_t (TweakeyGeneration_key_Feedback[47]), .B0_f (new_AGEMA_signal_2146), .B1_t (new_AGEMA_signal_2147), .B1_f (new_AGEMA_signal_2148), .Z0_t (TweakeyGeneration_key_Feedback[15]), .Z0_f (new_AGEMA_signal_1858), .Z1_t (new_AGEMA_signal_1859), .Z1_f (new_AGEMA_signal_1860) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_48_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[48]), .A0_f (new_AGEMA_signal_2155), .A1_t (new_AGEMA_signal_2156), .A1_f (new_AGEMA_signal_2157), .B0_t (Key_s0_t[48]), .B0_f (Key_s0_f[48]), .B1_t (Key_s1_t[48]), .B1_f (Key_s1_f[48]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_48_U1_X), .Z0_f (new_AGEMA_signal_2161), .Z1_t (new_AGEMA_signal_2162), .Z1_f (new_AGEMA_signal_2163) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_48_U1_X), .B0_f (new_AGEMA_signal_2161), .B1_t (new_AGEMA_signal_2162), .B1_f (new_AGEMA_signal_2163), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_48_U1_Y), .Z0_f (new_AGEMA_signal_2649), .Z1_t (new_AGEMA_signal_2650), .Z1_f (new_AGEMA_signal_2651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_48_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_48_U1_Y), .A0_f (new_AGEMA_signal_2649), .A1_t (new_AGEMA_signal_2650), .A1_f (new_AGEMA_signal_2651), .B0_t (TweakeyGeneration_key_Feedback[48]), .B0_f (new_AGEMA_signal_2155), .B1_t (new_AGEMA_signal_2156), .B1_f (new_AGEMA_signal_2157), .Z0_t (TweakeyGeneration_key_Feedback[16]), .Z0_f (new_AGEMA_signal_1867), .Z1_t (new_AGEMA_signal_1868), .Z1_f (new_AGEMA_signal_1869) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_49_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[49]), .A0_f (new_AGEMA_signal_2164), .A1_t (new_AGEMA_signal_2165), .A1_f (new_AGEMA_signal_2166), .B0_t (Key_s0_t[49]), .B0_f (Key_s0_f[49]), .B1_t (Key_s1_t[49]), .B1_f (Key_s1_f[49]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_49_U1_X), .Z0_f (new_AGEMA_signal_2170), .Z1_t (new_AGEMA_signal_2171), .Z1_f (new_AGEMA_signal_2172) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_49_U1_X), .B0_f (new_AGEMA_signal_2170), .B1_t (new_AGEMA_signal_2171), .B1_f (new_AGEMA_signal_2172), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_49_U1_Y), .Z0_f (new_AGEMA_signal_2652), .Z1_t (new_AGEMA_signal_2653), .Z1_f (new_AGEMA_signal_2654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_49_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_49_U1_Y), .A0_f (new_AGEMA_signal_2652), .A1_t (new_AGEMA_signal_2653), .A1_f (new_AGEMA_signal_2654), .B0_t (TweakeyGeneration_key_Feedback[49]), .B0_f (new_AGEMA_signal_2164), .B1_t (new_AGEMA_signal_2165), .B1_f (new_AGEMA_signal_2166), .Z0_t (TweakeyGeneration_key_Feedback[17]), .Z0_f (new_AGEMA_signal_1876), .Z1_t (new_AGEMA_signal_1877), .Z1_f (new_AGEMA_signal_1878) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_50_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[50]), .A0_f (new_AGEMA_signal_2173), .A1_t (new_AGEMA_signal_2174), .A1_f (new_AGEMA_signal_2175), .B0_t (Key_s0_t[50]), .B0_f (Key_s0_f[50]), .B1_t (Key_s1_t[50]), .B1_f (Key_s1_f[50]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_50_U1_X), .Z0_f (new_AGEMA_signal_2179), .Z1_t (new_AGEMA_signal_2180), .Z1_f (new_AGEMA_signal_2181) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_50_U1_X), .B0_f (new_AGEMA_signal_2179), .B1_t (new_AGEMA_signal_2180), .B1_f (new_AGEMA_signal_2181), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_50_U1_Y), .Z0_f (new_AGEMA_signal_2655), .Z1_t (new_AGEMA_signal_2656), .Z1_f (new_AGEMA_signal_2657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_50_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_50_U1_Y), .A0_f (new_AGEMA_signal_2655), .A1_t (new_AGEMA_signal_2656), .A1_f (new_AGEMA_signal_2657), .B0_t (TweakeyGeneration_key_Feedback[50]), .B0_f (new_AGEMA_signal_2173), .B1_t (new_AGEMA_signal_2174), .B1_f (new_AGEMA_signal_2175), .Z0_t (TweakeyGeneration_key_Feedback[18]), .Z0_f (new_AGEMA_signal_1885), .Z1_t (new_AGEMA_signal_1886), .Z1_f (new_AGEMA_signal_1887) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_51_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[51]), .A0_f (new_AGEMA_signal_2182), .A1_t (new_AGEMA_signal_2183), .A1_f (new_AGEMA_signal_2184), .B0_t (Key_s0_t[51]), .B0_f (Key_s0_f[51]), .B1_t (Key_s1_t[51]), .B1_f (Key_s1_f[51]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_51_U1_X), .Z0_f (new_AGEMA_signal_2188), .Z1_t (new_AGEMA_signal_2189), .Z1_f (new_AGEMA_signal_2190) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_51_U1_X), .B0_f (new_AGEMA_signal_2188), .B1_t (new_AGEMA_signal_2189), .B1_f (new_AGEMA_signal_2190), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_51_U1_Y), .Z0_f (new_AGEMA_signal_2658), .Z1_t (new_AGEMA_signal_2659), .Z1_f (new_AGEMA_signal_2660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_51_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_51_U1_Y), .A0_f (new_AGEMA_signal_2658), .A1_t (new_AGEMA_signal_2659), .A1_f (new_AGEMA_signal_2660), .B0_t (TweakeyGeneration_key_Feedback[51]), .B0_f (new_AGEMA_signal_2182), .B1_t (new_AGEMA_signal_2183), .B1_f (new_AGEMA_signal_2184), .Z0_t (TweakeyGeneration_key_Feedback[19]), .Z0_f (new_AGEMA_signal_1894), .Z1_t (new_AGEMA_signal_1895), .Z1_f (new_AGEMA_signal_1896) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_52_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[52]), .A0_f (new_AGEMA_signal_2191), .A1_t (new_AGEMA_signal_2192), .A1_f (new_AGEMA_signal_2193), .B0_t (Key_s0_t[52]), .B0_f (Key_s0_f[52]), .B1_t (Key_s1_t[52]), .B1_f (Key_s1_f[52]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_52_U1_X), .Z0_f (new_AGEMA_signal_2197), .Z1_t (new_AGEMA_signal_2198), .Z1_f (new_AGEMA_signal_2199) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_52_U1_X), .B0_f (new_AGEMA_signal_2197), .B1_t (new_AGEMA_signal_2198), .B1_f (new_AGEMA_signal_2199), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_52_U1_Y), .Z0_f (new_AGEMA_signal_2661), .Z1_t (new_AGEMA_signal_2662), .Z1_f (new_AGEMA_signal_2663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_52_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_52_U1_Y), .A0_f (new_AGEMA_signal_2661), .A1_t (new_AGEMA_signal_2662), .A1_f (new_AGEMA_signal_2663), .B0_t (TweakeyGeneration_key_Feedback[52]), .B0_f (new_AGEMA_signal_2191), .B1_t (new_AGEMA_signal_2192), .B1_f (new_AGEMA_signal_2193), .Z0_t (TweakeyGeneration_key_Feedback[20]), .Z0_f (new_AGEMA_signal_1903), .Z1_t (new_AGEMA_signal_1904), .Z1_f (new_AGEMA_signal_1905) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_53_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[53]), .A0_f (new_AGEMA_signal_2200), .A1_t (new_AGEMA_signal_2201), .A1_f (new_AGEMA_signal_2202), .B0_t (Key_s0_t[53]), .B0_f (Key_s0_f[53]), .B1_t (Key_s1_t[53]), .B1_f (Key_s1_f[53]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_53_U1_X), .Z0_f (new_AGEMA_signal_2206), .Z1_t (new_AGEMA_signal_2207), .Z1_f (new_AGEMA_signal_2208) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_53_U1_X), .B0_f (new_AGEMA_signal_2206), .B1_t (new_AGEMA_signal_2207), .B1_f (new_AGEMA_signal_2208), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_53_U1_Y), .Z0_f (new_AGEMA_signal_2664), .Z1_t (new_AGEMA_signal_2665), .Z1_f (new_AGEMA_signal_2666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_53_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_53_U1_Y), .A0_f (new_AGEMA_signal_2664), .A1_t (new_AGEMA_signal_2665), .A1_f (new_AGEMA_signal_2666), .B0_t (TweakeyGeneration_key_Feedback[53]), .B0_f (new_AGEMA_signal_2200), .B1_t (new_AGEMA_signal_2201), .B1_f (new_AGEMA_signal_2202), .Z0_t (TweakeyGeneration_key_Feedback[21]), .Z0_f (new_AGEMA_signal_1912), .Z1_t (new_AGEMA_signal_1913), .Z1_f (new_AGEMA_signal_1914) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_54_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[54]), .A0_f (new_AGEMA_signal_2209), .A1_t (new_AGEMA_signal_2210), .A1_f (new_AGEMA_signal_2211), .B0_t (Key_s0_t[54]), .B0_f (Key_s0_f[54]), .B1_t (Key_s1_t[54]), .B1_f (Key_s1_f[54]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_54_U1_X), .Z0_f (new_AGEMA_signal_2215), .Z1_t (new_AGEMA_signal_2216), .Z1_f (new_AGEMA_signal_2217) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_54_U1_X), .B0_f (new_AGEMA_signal_2215), .B1_t (new_AGEMA_signal_2216), .B1_f (new_AGEMA_signal_2217), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_54_U1_Y), .Z0_f (new_AGEMA_signal_2667), .Z1_t (new_AGEMA_signal_2668), .Z1_f (new_AGEMA_signal_2669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_54_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_54_U1_Y), .A0_f (new_AGEMA_signal_2667), .A1_t (new_AGEMA_signal_2668), .A1_f (new_AGEMA_signal_2669), .B0_t (TweakeyGeneration_key_Feedback[54]), .B0_f (new_AGEMA_signal_2209), .B1_t (new_AGEMA_signal_2210), .B1_f (new_AGEMA_signal_2211), .Z0_t (TweakeyGeneration_key_Feedback[22]), .Z0_f (new_AGEMA_signal_1921), .Z1_t (new_AGEMA_signal_1922), .Z1_f (new_AGEMA_signal_1923) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_55_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[55]), .A0_f (new_AGEMA_signal_2218), .A1_t (new_AGEMA_signal_2219), .A1_f (new_AGEMA_signal_2220), .B0_t (Key_s0_t[55]), .B0_f (Key_s0_f[55]), .B1_t (Key_s1_t[55]), .B1_f (Key_s1_f[55]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_55_U1_X), .Z0_f (new_AGEMA_signal_2224), .Z1_t (new_AGEMA_signal_2225), .Z1_f (new_AGEMA_signal_2226) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_55_U1_X), .B0_f (new_AGEMA_signal_2224), .B1_t (new_AGEMA_signal_2225), .B1_f (new_AGEMA_signal_2226), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_55_U1_Y), .Z0_f (new_AGEMA_signal_2670), .Z1_t (new_AGEMA_signal_2671), .Z1_f (new_AGEMA_signal_2672) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_55_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_55_U1_Y), .A0_f (new_AGEMA_signal_2670), .A1_t (new_AGEMA_signal_2671), .A1_f (new_AGEMA_signal_2672), .B0_t (TweakeyGeneration_key_Feedback[55]), .B0_f (new_AGEMA_signal_2218), .B1_t (new_AGEMA_signal_2219), .B1_f (new_AGEMA_signal_2220), .Z0_t (TweakeyGeneration_key_Feedback[23]), .Z0_f (new_AGEMA_signal_1930), .Z1_t (new_AGEMA_signal_1931), .Z1_f (new_AGEMA_signal_1932) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_56_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[56]), .A0_f (new_AGEMA_signal_2227), .A1_t (new_AGEMA_signal_2228), .A1_f (new_AGEMA_signal_2229), .B0_t (Key_s0_t[56]), .B0_f (Key_s0_f[56]), .B1_t (Key_s1_t[56]), .B1_f (Key_s1_f[56]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_56_U1_X), .Z0_f (new_AGEMA_signal_2233), .Z1_t (new_AGEMA_signal_2234), .Z1_f (new_AGEMA_signal_2235) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_56_U1_X), .B0_f (new_AGEMA_signal_2233), .B1_t (new_AGEMA_signal_2234), .B1_f (new_AGEMA_signal_2235), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_56_U1_Y), .Z0_f (new_AGEMA_signal_2673), .Z1_t (new_AGEMA_signal_2674), .Z1_f (new_AGEMA_signal_2675) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_56_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_56_U1_Y), .A0_f (new_AGEMA_signal_2673), .A1_t (new_AGEMA_signal_2674), .A1_f (new_AGEMA_signal_2675), .B0_t (TweakeyGeneration_key_Feedback[56]), .B0_f (new_AGEMA_signal_2227), .B1_t (new_AGEMA_signal_2228), .B1_f (new_AGEMA_signal_2229), .Z0_t (TweakeyGeneration_key_Feedback[24]), .Z0_f (new_AGEMA_signal_1939), .Z1_t (new_AGEMA_signal_1940), .Z1_f (new_AGEMA_signal_1941) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_57_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[57]), .A0_f (new_AGEMA_signal_2236), .A1_t (new_AGEMA_signal_2237), .A1_f (new_AGEMA_signal_2238), .B0_t (Key_s0_t[57]), .B0_f (Key_s0_f[57]), .B1_t (Key_s1_t[57]), .B1_f (Key_s1_f[57]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_57_U1_X), .Z0_f (new_AGEMA_signal_2242), .Z1_t (new_AGEMA_signal_2243), .Z1_f (new_AGEMA_signal_2244) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_57_U1_X), .B0_f (new_AGEMA_signal_2242), .B1_t (new_AGEMA_signal_2243), .B1_f (new_AGEMA_signal_2244), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_57_U1_Y), .Z0_f (new_AGEMA_signal_2676), .Z1_t (new_AGEMA_signal_2677), .Z1_f (new_AGEMA_signal_2678) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_57_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_57_U1_Y), .A0_f (new_AGEMA_signal_2676), .A1_t (new_AGEMA_signal_2677), .A1_f (new_AGEMA_signal_2678), .B0_t (TweakeyGeneration_key_Feedback[57]), .B0_f (new_AGEMA_signal_2236), .B1_t (new_AGEMA_signal_2237), .B1_f (new_AGEMA_signal_2238), .Z0_t (TweakeyGeneration_key_Feedback[25]), .Z0_f (new_AGEMA_signal_1948), .Z1_t (new_AGEMA_signal_1949), .Z1_f (new_AGEMA_signal_1950) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_58_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[58]), .A0_f (new_AGEMA_signal_2245), .A1_t (new_AGEMA_signal_2246), .A1_f (new_AGEMA_signal_2247), .B0_t (Key_s0_t[58]), .B0_f (Key_s0_f[58]), .B1_t (Key_s1_t[58]), .B1_f (Key_s1_f[58]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_58_U1_X), .Z0_f (new_AGEMA_signal_2251), .Z1_t (new_AGEMA_signal_2252), .Z1_f (new_AGEMA_signal_2253) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_58_U1_X), .B0_f (new_AGEMA_signal_2251), .B1_t (new_AGEMA_signal_2252), .B1_f (new_AGEMA_signal_2253), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_58_U1_Y), .Z0_f (new_AGEMA_signal_2679), .Z1_t (new_AGEMA_signal_2680), .Z1_f (new_AGEMA_signal_2681) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_58_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_58_U1_Y), .A0_f (new_AGEMA_signal_2679), .A1_t (new_AGEMA_signal_2680), .A1_f (new_AGEMA_signal_2681), .B0_t (TweakeyGeneration_key_Feedback[58]), .B0_f (new_AGEMA_signal_2245), .B1_t (new_AGEMA_signal_2246), .B1_f (new_AGEMA_signal_2247), .Z0_t (TweakeyGeneration_key_Feedback[26]), .Z0_f (new_AGEMA_signal_1957), .Z1_t (new_AGEMA_signal_1958), .Z1_f (new_AGEMA_signal_1959) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_59_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[59]), .A0_f (new_AGEMA_signal_2254), .A1_t (new_AGEMA_signal_2255), .A1_f (new_AGEMA_signal_2256), .B0_t (Key_s0_t[59]), .B0_f (Key_s0_f[59]), .B1_t (Key_s1_t[59]), .B1_f (Key_s1_f[59]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_59_U1_X), .Z0_f (new_AGEMA_signal_2260), .Z1_t (new_AGEMA_signal_2261), .Z1_f (new_AGEMA_signal_2262) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_59_U1_X), .B0_f (new_AGEMA_signal_2260), .B1_t (new_AGEMA_signal_2261), .B1_f (new_AGEMA_signal_2262), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_59_U1_Y), .Z0_f (new_AGEMA_signal_2682), .Z1_t (new_AGEMA_signal_2683), .Z1_f (new_AGEMA_signal_2684) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_59_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_59_U1_Y), .A0_f (new_AGEMA_signal_2682), .A1_t (new_AGEMA_signal_2683), .A1_f (new_AGEMA_signal_2684), .B0_t (TweakeyGeneration_key_Feedback[59]), .B0_f (new_AGEMA_signal_2254), .B1_t (new_AGEMA_signal_2255), .B1_f (new_AGEMA_signal_2256), .Z0_t (TweakeyGeneration_key_Feedback[27]), .Z0_f (new_AGEMA_signal_1966), .Z1_t (new_AGEMA_signal_1967), .Z1_f (new_AGEMA_signal_1968) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_60_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[60]), .A0_f (new_AGEMA_signal_2263), .A1_t (new_AGEMA_signal_2264), .A1_f (new_AGEMA_signal_2265), .B0_t (Key_s0_t[60]), .B0_f (Key_s0_f[60]), .B1_t (Key_s1_t[60]), .B1_f (Key_s1_f[60]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_60_U1_X), .Z0_f (new_AGEMA_signal_2269), .Z1_t (new_AGEMA_signal_2270), .Z1_f (new_AGEMA_signal_2271) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_60_U1_X), .B0_f (new_AGEMA_signal_2269), .B1_t (new_AGEMA_signal_2270), .B1_f (new_AGEMA_signal_2271), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_60_U1_Y), .Z0_f (new_AGEMA_signal_2685), .Z1_t (new_AGEMA_signal_2686), .Z1_f (new_AGEMA_signal_2687) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_60_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_60_U1_Y), .A0_f (new_AGEMA_signal_2685), .A1_t (new_AGEMA_signal_2686), .A1_f (new_AGEMA_signal_2687), .B0_t (TweakeyGeneration_key_Feedback[60]), .B0_f (new_AGEMA_signal_2263), .B1_t (new_AGEMA_signal_2264), .B1_f (new_AGEMA_signal_2265), .Z0_t (TweakeyGeneration_key_Feedback[28]), .Z0_f (new_AGEMA_signal_1975), .Z1_t (new_AGEMA_signal_1976), .Z1_f (new_AGEMA_signal_1977) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_61_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[61]), .A0_f (new_AGEMA_signal_2272), .A1_t (new_AGEMA_signal_2273), .A1_f (new_AGEMA_signal_2274), .B0_t (Key_s0_t[61]), .B0_f (Key_s0_f[61]), .B1_t (Key_s1_t[61]), .B1_f (Key_s1_f[61]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_61_U1_X), .Z0_f (new_AGEMA_signal_2278), .Z1_t (new_AGEMA_signal_2279), .Z1_f (new_AGEMA_signal_2280) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_61_U1_X), .B0_f (new_AGEMA_signal_2278), .B1_t (new_AGEMA_signal_2279), .B1_f (new_AGEMA_signal_2280), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_61_U1_Y), .Z0_f (new_AGEMA_signal_2688), .Z1_t (new_AGEMA_signal_2689), .Z1_f (new_AGEMA_signal_2690) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_61_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_61_U1_Y), .A0_f (new_AGEMA_signal_2688), .A1_t (new_AGEMA_signal_2689), .A1_f (new_AGEMA_signal_2690), .B0_t (TweakeyGeneration_key_Feedback[61]), .B0_f (new_AGEMA_signal_2272), .B1_t (new_AGEMA_signal_2273), .B1_f (new_AGEMA_signal_2274), .Z0_t (TweakeyGeneration_key_Feedback[29]), .Z0_f (new_AGEMA_signal_1984), .Z1_t (new_AGEMA_signal_1985), .Z1_f (new_AGEMA_signal_1986) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_62_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[62]), .A0_f (new_AGEMA_signal_2281), .A1_t (new_AGEMA_signal_2282), .A1_f (new_AGEMA_signal_2283), .B0_t (Key_s0_t[62]), .B0_f (Key_s0_f[62]), .B1_t (Key_s1_t[62]), .B1_f (Key_s1_f[62]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_62_U1_X), .Z0_f (new_AGEMA_signal_2287), .Z1_t (new_AGEMA_signal_2288), .Z1_f (new_AGEMA_signal_2289) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_62_U1_X), .B0_f (new_AGEMA_signal_2287), .B1_t (new_AGEMA_signal_2288), .B1_f (new_AGEMA_signal_2289), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_62_U1_Y), .Z0_f (new_AGEMA_signal_2691), .Z1_t (new_AGEMA_signal_2692), .Z1_f (new_AGEMA_signal_2693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_62_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_62_U1_Y), .A0_f (new_AGEMA_signal_2691), .A1_t (new_AGEMA_signal_2692), .A1_f (new_AGEMA_signal_2693), .B0_t (TweakeyGeneration_key_Feedback[62]), .B0_f (new_AGEMA_signal_2281), .B1_t (new_AGEMA_signal_2282), .B1_f (new_AGEMA_signal_2283), .Z0_t (TweakeyGeneration_key_Feedback[30]), .Z0_f (new_AGEMA_signal_1993), .Z1_t (new_AGEMA_signal_1994), .Z1_f (new_AGEMA_signal_1995) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_63_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[63]), .A0_f (new_AGEMA_signal_2290), .A1_t (new_AGEMA_signal_2291), .A1_f (new_AGEMA_signal_2292), .B0_t (Key_s0_t[63]), .B0_f (Key_s0_f[63]), .B1_t (Key_s1_t[63]), .B1_f (Key_s1_f[63]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_63_U1_X), .Z0_f (new_AGEMA_signal_2296), .Z1_t (new_AGEMA_signal_2297), .Z1_f (new_AGEMA_signal_2298) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_63_U1_X), .B0_f (new_AGEMA_signal_2296), .B1_t (new_AGEMA_signal_2297), .B1_f (new_AGEMA_signal_2298), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_63_U1_Y), .Z0_f (new_AGEMA_signal_2694), .Z1_t (new_AGEMA_signal_2695), .Z1_f (new_AGEMA_signal_2696) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_63_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_63_U1_Y), .A0_f (new_AGEMA_signal_2694), .A1_t (new_AGEMA_signal_2695), .A1_f (new_AGEMA_signal_2696), .B0_t (TweakeyGeneration_key_Feedback[63]), .B0_f (new_AGEMA_signal_2290), .B1_t (new_AGEMA_signal_2291), .B1_f (new_AGEMA_signal_2292), .Z0_t (TweakeyGeneration_key_Feedback[31]), .Z0_f (new_AGEMA_signal_2002), .Z1_t (new_AGEMA_signal_2003), .Z1_f (new_AGEMA_signal_2004) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_0_U1 ( .A0_t (FSMUpdate[0]), .A0_f (new_AGEMA_signal_3362), .B0_t (rst_t), .B0_f (rst_f), .Z0_t (FSMUpdate[1]), .Z0_f (new_AGEMA_signal_2300) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_1_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (FSMUpdate[1]), .B0_f (new_AGEMA_signal_2300), .Z0_t (FSM[1]), .Z0_f (new_AGEMA_signal_2301) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_2_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (FSMUpdate[2]), .B0_f (new_AGEMA_signal_3216), .Z0_t (FSMUpdate[3]), .Z0_f (new_AGEMA_signal_2302) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_3_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (FSMUpdate[3]), .B0_f (new_AGEMA_signal_2302), .Z0_t (FSMUpdate[4]), .Z0_f (new_AGEMA_signal_2303) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_4_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (FSMUpdate[4]), .B0_f (new_AGEMA_signal_2303), .Z0_t (FSM[4]), .Z0_f (new_AGEMA_signal_2304) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_5_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (FSMUpdate[5]), .B0_f (new_AGEMA_signal_3217), .Z0_t (FSM[5]), .Z0_f (new_AGEMA_signal_2309) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_0_U4 ( .A0_t (FSM[5]), .A0_f (new_AGEMA_signal_2309), .B0_t (FSMUpdateInst_StateUpdateInst_0_n3), .B0_f (new_AGEMA_signal_2697), .Z0_t (FSMUpdateInst_StateUpdateInst_0_n4), .Z0_f (new_AGEMA_signal_2845) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_0_U3 ( .A0_t (FSMUpdateInst_StateUpdateInst_0_n2), .A0_f (new_AGEMA_signal_2306), .B0_t (FSMUpdateInst_StateUpdateInst_0_n1), .B0_f (new_AGEMA_signal_2305), .Z0_t (FSMUpdateInst_StateUpdateInst_0_n3), .Z0_f (new_AGEMA_signal_2697) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_0_U2 ( .A0_t (FSMUpdate[4]), .A0_f (new_AGEMA_signal_2303), .B0_t (FSMUpdate[3]), .B0_f (new_AGEMA_signal_2302), .Z0_t (FSMUpdateInst_StateUpdateInst_0_n1), .Z0_f (new_AGEMA_signal_2305) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_0_U1 ( .A0_t (FSMUpdate[1]), .A0_f (new_AGEMA_signal_2300), .B0_t (FSM[1]), .B0_f (new_AGEMA_signal_2301), .Z0_t (FSMUpdateInst_StateUpdateInst_0_n2), .Z0_f (new_AGEMA_signal_2306) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) FSMUpdateInst_StateUpdateInst_0_U7_XOR1_U1 ( .A0_t (FSMUpdateInst_StateUpdateInst_0_n4), .A0_f (new_AGEMA_signal_2845), .B0_t (FSM[5]), .B0_f (new_AGEMA_signal_2309), .Z0_t (FSMUpdateInst_StateUpdateInst_0_U7_X), .Z0_f (new_AGEMA_signal_3017) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_0_U7_AND1_U1 ( .A0_t (FSM[4]), .A0_f (new_AGEMA_signal_2304), .B0_t (FSMUpdateInst_StateUpdateInst_0_U7_X), .B0_f (new_AGEMA_signal_3017), .Z0_t (FSMUpdateInst_StateUpdateInst_0_U7_Y), .Z0_f (new_AGEMA_signal_3215) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) FSMUpdateInst_StateUpdateInst_0_U7_XOR2_U1 ( .A0_t (FSMUpdateInst_StateUpdateInst_0_U7_Y), .A0_f (new_AGEMA_signal_3215), .B0_t (FSMUpdateInst_StateUpdateInst_0_n4), .B0_f (new_AGEMA_signal_2845), .Z0_t (FSMUpdate[0]), .Z0_f (new_AGEMA_signal_3362) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_2_U5 ( .A0_t (FSMUpdateInst_StateUpdateInst_2_n4), .A0_f (new_AGEMA_signal_3018), .B0_t (FSM[1]), .B0_f (new_AGEMA_signal_2301), .Z0_t (FSMUpdate[2]), .Z0_f (new_AGEMA_signal_3216) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_2_U4 ( .A0_t (FSMUpdateInst_StateUpdateInst_2_n3), .A0_f (new_AGEMA_signal_2846), .B0_t (FSM[5]), .B0_f (new_AGEMA_signal_2309), .Z0_t (FSMUpdateInst_StateUpdateInst_2_n4), .Z0_f (new_AGEMA_signal_3018) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_2_U3 ( .A0_t (FSM[4]), .A0_f (new_AGEMA_signal_2304), .B0_t (FSMUpdateInst_StateUpdateInst_2_n2), .B0_f (new_AGEMA_signal_2698), .Z0_t (FSMUpdateInst_StateUpdateInst_2_n3), .Z0_f (new_AGEMA_signal_2846) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_2_U2 ( .A0_t (FSMUpdate[1]), .A0_f (new_AGEMA_signal_2300), .B0_t (FSMUpdateInst_StateUpdateInst_2_n1), .B0_f (new_AGEMA_signal_2307), .Z0_t (FSMUpdateInst_StateUpdateInst_2_n2), .Z0_f (new_AGEMA_signal_2698) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_2_U1 ( .A0_t (FSMUpdate[4]), .A0_f (new_AGEMA_signal_2303), .B0_t (FSMUpdate[3]), .B0_f (new_AGEMA_signal_2302), .Z0_t (FSMUpdateInst_StateUpdateInst_2_n1), .Z0_f (new_AGEMA_signal_2307) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_5_U5 ( .A0_t (FSM[4]), .A0_f (new_AGEMA_signal_2304), .B0_t (FSMUpdateInst_StateUpdateInst_5_n4), .B0_f (new_AGEMA_signal_3019), .Z0_t (FSMUpdate[5]), .Z0_f (new_AGEMA_signal_3217) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_5_U4 ( .A0_t (FSMUpdate[4]), .A0_f (new_AGEMA_signal_2303), .B0_t (FSMUpdateInst_StateUpdateInst_5_n3), .B0_f (new_AGEMA_signal_2847), .Z0_t (FSMUpdateInst_StateUpdateInst_5_n4), .Z0_f (new_AGEMA_signal_3019) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_5_U3 ( .A0_t (FSM[5]), .A0_f (new_AGEMA_signal_2309), .B0_t (FSMUpdateInst_StateUpdateInst_5_n2), .B0_f (new_AGEMA_signal_2699), .Z0_t (FSMUpdateInst_StateUpdateInst_5_n3), .Z0_f (new_AGEMA_signal_2847) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_5_U2 ( .A0_t (FSMUpdate[3]), .A0_f (new_AGEMA_signal_2302), .B0_t (FSMUpdateInst_StateUpdateInst_5_n1), .B0_f (new_AGEMA_signal_2308), .Z0_t (FSMUpdateInst_StateUpdateInst_5_n2), .Z0_f (new_AGEMA_signal_2699) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_5_U1 ( .A0_t (FSMUpdate[1]), .A0_f (new_AGEMA_signal_2300), .B0_t (FSM[1]), .B0_f (new_AGEMA_signal_2301), .Z0_t (FSMUpdateInst_StateUpdateInst_5_n1), .Z0_f (new_AGEMA_signal_2308) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_doneInst_U6 ( .A0_t (FSMSignalsInst_doneInst_n5), .A0_f (new_AGEMA_signal_2700), .B0_t (FSMSignalsInst_doneInst_n4), .B0_f (new_AGEMA_signal_2310), .Z0_t (done_t), .Z0_f (done_f) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_doneInst_U5 ( .A0_t (FSM[4]), .A0_f (new_AGEMA_signal_2304), .B0_t (FSM[5]), .B0_f (new_AGEMA_signal_2309), .Z0_t (FSMSignalsInst_doneInst_n4), .Z0_f (new_AGEMA_signal_2310) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_doneInst_U4 ( .A0_t (FSMSignalsInst_doneInst_n3), .A0_f (new_AGEMA_signal_2312), .B0_t (FSMSignalsInst_doneInst_n2), .B0_f (new_AGEMA_signal_2311), .Z0_t (FSMSignalsInst_doneInst_n5), .Z0_f (new_AGEMA_signal_2700) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_doneInst_U3 ( .A0_t (FSMUpdate[4]), .A0_f (new_AGEMA_signal_2303), .B0_t (FSMUpdate[1]), .B0_f (new_AGEMA_signal_2300), .Z0_t (FSMSignalsInst_doneInst_n2), .Z0_f (new_AGEMA_signal_2311) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_doneInst_U1 ( .A0_t (FSMUpdate[3]), .A0_f (new_AGEMA_signal_2302), .B0_t (FSM[1]), .B0_f (new_AGEMA_signal_2301), .Z0_t (FSMSignalsInst_doneInst_n3), .Z0_f (new_AGEMA_signal_2312) ) ;

    /* register cells */
endmodule
