 // NumberOfConfigBits: 192
module ctrl_to_sec_switch_matrix
    #(
        parameter NoConfigBits=192
    )
    (
        input from_EA0,
        input from_EA1,
        input from_EA2,
        input from_EA3,
        input from_EB0,
        input from_EB1,
        input from_EB2,
        input from_EB3,
        input from_EC0,
        input from_EC1,
        input from_EC2,
        input from_EC3,
        input from_ED0,
        input from_ED1,
        input from_ED2,
        input from_ED3,
        input from_EF0,
        input from_EF1,
        input from_EF2,
        input from_EF3,
        input from_EG0,
        input from_EG1,
        input from_EG2,
        input from_EG3,
        input from_EG4,
        input from_EG5,
        input from_EG6,
        input from_EG7,
        input from_EH0,
        input from_EH1,
        input from_EH2,
        input from_EH3,
        input from_EH4,
        input from_EH5,
        input from_EH6,
        input from_EH7,
        input from_EI0,
        input from_EI1,
        input from_EI2,
        input from_EI3,
        input from_EI4,
        input from_EI5,
        input from_EI6,
        input from_EI7,
        input from_EI8,
        input from_EI9,
        input from_EI10,
        input from_EI11,
        input from_WA_1s0,
        input from_WA_1s1,
        input from_WB_1s0,
        input from_WB_1s1,
        input from_WC_1s0,
        input from_WC_1s1,
        input from_WD_1s0,
        input from_WD_1s1,
        input from_WF_1s0,
        input from_WF_1s1,
        input from_WG_1s0,
        input from_WG_1s1,
        input from_WH_1s0,
        input from_WH_1s1,
        input from_WI_1s0,
        input from_WI_1s1,
        input from_NA0,
        input from_NA1,
        input from_NA2,
        input from_NA3,
        input from_NB0,
        input from_NB1,
        input from_NB2,
        input from_NB3,
        input from_NC0,
        input from_NC1,
        input from_NC2,
        input from_NC3,
        input from_ND0,
        input from_ND1,
        input from_ND2,
        input from_ND3,
        input from_NF0,
        input from_NF1,
        input from_NF2,
        input from_NF3,
        input from_NG0,
        input from_NG1,
        input from_NG2,
        input from_NG3,
        input from_NH0,
        input from_NH1,
        input from_NH2,
        input from_NH3,
        input from_NI0,
        input from_NI1,
        input from_NI2,
        input from_NI3,
        input from_SA0,
        input from_SA1,
        input from_SA2,
        input from_SA3,
        input from_SB0,
        input from_SB1,
        input from_SB2,
        input from_SB3,
        input from_SC0,
        input from_SC1,
        input from_SC2,
        input from_SC3,
        input from_SD0,
        input from_SD1,
        input from_SD2,
        input from_SD3,
        input from_SF0,
        input from_SF1,
        input from_SF2,
        input from_SF3,
        input from_SG0,
        input from_SG1,
        input from_SG2,
        input from_SG3,
        input from_SH0,
        input from_SH1,
        input from_SH2,
        input from_SH3,
        input from_SI0,
        input from_SI1,
        input from_SI2,
        input from_SI3,
        output to_WA0,
        output to_WA1,
        output to_WA2,
        output to_WA3,
        output to_WB0,
        output to_WB1,
        output to_WB2,
        output to_WB3,
        output to_WC0,
        output to_WC1,
        output to_WC2,
        output to_WC3,
        output to_WD0,
        output to_WD1,
        output to_WD2,
        output to_WD3,
        output to_WF0,
        output to_WF1,
        output to_WF2,
        output to_WF3,
        output to_WG0,
        output to_WG1,
        output to_WG2,
        output to_WG3,
        output to_WG4,
        output to_WG5,
        output to_WG6,
        output to_WG7,
        output to_WH0,
        output to_WH1,
        output to_WH2,
        output to_WH3,
        output to_WH4,
        output to_WH5,
        output to_WH6,
        output to_WH7,
        output to_WI0,
        output to_WI1,
        output to_WI2,
        output to_WI3,
        output to_WI4,
        output to_WI5,
        output to_WI6,
        output to_WI7,
        output to_WI8,
        output to_WI9,
        output to_WI10,
        output to_WI11,
        output to_NA0,
        output to_NA1,
        output to_NA2,
        output to_NA3,
        output to_NB0,
        output to_NB1,
        output to_NB2,
        output to_NB3,
        output to_NC0,
        output to_NC1,
        output to_NC2,
        output to_NC3,
        output to_ND0,
        output to_ND1,
        output to_ND2,
        output to_ND3,
        output to_NF0,
        output to_NF1,
        output to_NF2,
        output to_NF3,
        output to_NG0,
        output to_NG1,
        output to_NG2,
        output to_NG3,
        output to_NH0,
        output to_NH1,
        output to_NH2,
        output to_NH3,
        output to_NI0,
        output to_NI1,
        output to_NI2,
        output to_NI3,
        output to_SA0,
        output to_SA1,
        output to_SA2,
        output to_SA3,
        output to_SB0,
        output to_SB1,
        output to_SB2,
        output to_SB3,
        output to_SC0,
        output to_SC1,
        output to_SC2,
        output to_SC3,
        output to_SD0,
        output to_SD1,
        output to_SD2,
        output to_SD3,
        output to_SF0,
        output to_SF1,
        output to_SF2,
        output to_SF3,
        output to_SG0,
        output to_SG1,
        output to_SG2,
        output to_SG3,
        output to_SH0,
        output to_SH1,
        output to_SH2,
        output to_SH3,
        output to_SI0,
        output to_SI1,
        output to_SI2,
        output to_SI3,
 //global
        input [NoConfigBits-1:0] ConfigBits,
        input [NoConfigBits-1:0] ConfigBits_N
);
parameter GND0 = 1'b0;
parameter GND = 1'b0;
parameter VCC0 = 1'b1;
parameter VCC = 1'b1;
parameter VDD0 = 1'b1;
parameter VDD = 1'b1;

wire[4-1:0] to_WA0_input;
wire[4-1:0] to_WA1_input;
wire[4-1:0] to_WA2_input;
wire[4-1:0] to_WA3_input;
wire[4-1:0] to_WB0_input;
wire[4-1:0] to_WB1_input;
wire[4-1:0] to_WB2_input;
wire[4-1:0] to_WB3_input;
wire[4-1:0] to_WC0_input;
wire[4-1:0] to_WC1_input;
wire[4-1:0] to_WC2_input;
wire[4-1:0] to_WC3_input;
wire[4-1:0] to_WD0_input;
wire[4-1:0] to_WD1_input;
wire[4-1:0] to_WD2_input;
wire[4-1:0] to_WD3_input;
wire[4-1:0] to_WF0_input;
wire[4-1:0] to_WF1_input;
wire[4-1:0] to_WF2_input;
wire[4-1:0] to_WF3_input;
wire[4-1:0] to_WG0_input;
wire[4-1:0] to_WG1_input;
wire[4-1:0] to_WG2_input;
wire[4-1:0] to_WG3_input;
wire[1-1:0] to_WG4_input;
wire[1-1:0] to_WG5_input;
wire[1-1:0] to_WG6_input;
wire[1-1:0] to_WG7_input;
wire[4-1:0] to_WH0_input;
wire[4-1:0] to_WH1_input;
wire[4-1:0] to_WH2_input;
wire[4-1:0] to_WH3_input;
wire[1-1:0] to_WH4_input;
wire[1-1:0] to_WH5_input;
wire[1-1:0] to_WH6_input;
wire[1-1:0] to_WH7_input;
wire[4-1:0] to_WI0_input;
wire[4-1:0] to_WI1_input;
wire[4-1:0] to_WI2_input;
wire[4-1:0] to_WI3_input;
wire[1-1:0] to_WI4_input;
wire[1-1:0] to_WI5_input;
wire[1-1:0] to_WI6_input;
wire[1-1:0] to_WI7_input;
wire[1-1:0] to_WI8_input;
wire[1-1:0] to_WI9_input;
wire[1-1:0] to_WI10_input;
wire[1-1:0] to_WI11_input;
wire[4-1:0] to_NA0_input;
wire[4-1:0] to_NA1_input;
wire[4-1:0] to_NA2_input;
wire[4-1:0] to_NA3_input;
wire[4-1:0] to_NB0_input;
wire[4-1:0] to_NB1_input;
wire[4-1:0] to_NB2_input;
wire[4-1:0] to_NB3_input;
wire[4-1:0] to_NC0_input;
wire[4-1:0] to_NC1_input;
wire[4-1:0] to_NC2_input;
wire[4-1:0] to_NC3_input;
wire[4-1:0] to_ND0_input;
wire[4-1:0] to_ND1_input;
wire[4-1:0] to_ND2_input;
wire[4-1:0] to_ND3_input;
wire[4-1:0] to_NF0_input;
wire[4-1:0] to_NF1_input;
wire[4-1:0] to_NF2_input;
wire[4-1:0] to_NF3_input;
wire[4-1:0] to_NG0_input;
wire[4-1:0] to_NG1_input;
wire[4-1:0] to_NG2_input;
wire[4-1:0] to_NG3_input;
wire[4-1:0] to_NH0_input;
wire[4-1:0] to_NH1_input;
wire[4-1:0] to_NH2_input;
wire[4-1:0] to_NH3_input;
wire[4-1:0] to_NI0_input;
wire[4-1:0] to_NI1_input;
wire[4-1:0] to_NI2_input;
wire[4-1:0] to_NI3_input;
wire[4-1:0] to_SA0_input;
wire[4-1:0] to_SA1_input;
wire[4-1:0] to_SA2_input;
wire[4-1:0] to_SA3_input;
wire[4-1:0] to_SB0_input;
wire[4-1:0] to_SB1_input;
wire[4-1:0] to_SB2_input;
wire[4-1:0] to_SB3_input;
wire[4-1:0] to_SC0_input;
wire[4-1:0] to_SC1_input;
wire[4-1:0] to_SC2_input;
wire[4-1:0] to_SC3_input;
wire[4-1:0] to_SD0_input;
wire[4-1:0] to_SD1_input;
wire[4-1:0] to_SD2_input;
wire[4-1:0] to_SD3_input;
wire[4-1:0] to_SF0_input;
wire[4-1:0] to_SF1_input;
wire[4-1:0] to_SF2_input;
wire[4-1:0] to_SF3_input;
wire[4-1:0] to_SG0_input;
wire[4-1:0] to_SG1_input;
wire[4-1:0] to_SG2_input;
wire[4-1:0] to_SG3_input;
wire[4-1:0] to_SH0_input;
wire[4-1:0] to_SH1_input;
wire[4-1:0] to_SH2_input;
wire[4-1:0] to_SH3_input;
wire[4-1:0] to_SI0_input;
wire[4-1:0] to_SI1_input;
wire[4-1:0] to_SI2_input;
wire[4-1:0] to_SI3_input;
 //The configuration bits (if any) are just a long shift register
 //This shift register is padded to an even number of flops/latches
 //switch matrix multiplexer to_WA0 MUX-4
assign to_WA0_input = {GND0,from_SA0,from_NA0,from_EA0};
cus_mux41_buf inst_cus_mux41_buf_to_WA0 (
    .A0(to_WA0_input[0]),
    .A1(to_WA0_input[1]),
    .A2(to_WA0_input[2]),
    .A3(to_WA0_input[3]),
    .S0(ConfigBits[0+0]),
    .S0N(ConfigBits_N[0+0]),
    .S1(ConfigBits[0+1]),
    .S1N(ConfigBits_N[0+1]),
    .X(to_WA0)
);

 //switch matrix multiplexer to_WA1 MUX-4
assign to_WA1_input = {VCC0,from_SA1,from_NA1,from_EA1};
cus_mux41_buf inst_cus_mux41_buf_to_WA1 (
    .A0(to_WA1_input[0]),
    .A1(to_WA1_input[1]),
    .A2(to_WA1_input[2]),
    .A3(to_WA1_input[3]),
    .S0(ConfigBits[2+0]),
    .S0N(ConfigBits_N[2+0]),
    .S1(ConfigBits[2+1]),
    .S1N(ConfigBits_N[2+1]),
    .X(to_WA1)
);

 //switch matrix multiplexer to_WA2 MUX-4
assign to_WA2_input = {from_SA2,from_NA2,from_WA_1s0,from_EA2};
cus_mux41_buf inst_cus_mux41_buf_to_WA2 (
    .A0(to_WA2_input[0]),
    .A1(to_WA2_input[1]),
    .A2(to_WA2_input[2]),
    .A3(to_WA2_input[3]),
    .S0(ConfigBits[4+0]),
    .S0N(ConfigBits_N[4+0]),
    .S1(ConfigBits[4+1]),
    .S1N(ConfigBits_N[4+1]),
    .X(to_WA2)
);

 //switch matrix multiplexer to_WA3 MUX-4
assign to_WA3_input = {from_SA3,from_NA3,from_WA_1s1,from_EA3};
cus_mux41_buf inst_cus_mux41_buf_to_WA3 (
    .A0(to_WA3_input[0]),
    .A1(to_WA3_input[1]),
    .A2(to_WA3_input[2]),
    .A3(to_WA3_input[3]),
    .S0(ConfigBits[6+0]),
    .S0N(ConfigBits_N[6+0]),
    .S1(ConfigBits[6+1]),
    .S1N(ConfigBits_N[6+1]),
    .X(to_WA3)
);

 //switch matrix multiplexer to_WB0 MUX-4
assign to_WB0_input = {GND0,from_SB0,from_NB0,from_EB0};
cus_mux41_buf inst_cus_mux41_buf_to_WB0 (
    .A0(to_WB0_input[0]),
    .A1(to_WB0_input[1]),
    .A2(to_WB0_input[2]),
    .A3(to_WB0_input[3]),
    .S0(ConfigBits[8+0]),
    .S0N(ConfigBits_N[8+0]),
    .S1(ConfigBits[8+1]),
    .S1N(ConfigBits_N[8+1]),
    .X(to_WB0)
);

 //switch matrix multiplexer to_WB1 MUX-4
assign to_WB1_input = {VCC0,from_SB1,from_NB1,from_EB1};
cus_mux41_buf inst_cus_mux41_buf_to_WB1 (
    .A0(to_WB1_input[0]),
    .A1(to_WB1_input[1]),
    .A2(to_WB1_input[2]),
    .A3(to_WB1_input[3]),
    .S0(ConfigBits[10+0]),
    .S0N(ConfigBits_N[10+0]),
    .S1(ConfigBits[10+1]),
    .S1N(ConfigBits_N[10+1]),
    .X(to_WB1)
);

 //switch matrix multiplexer to_WB2 MUX-4
assign to_WB2_input = {from_SB2,from_NB2,from_WB_1s0,from_EB2};
cus_mux41_buf inst_cus_mux41_buf_to_WB2 (
    .A0(to_WB2_input[0]),
    .A1(to_WB2_input[1]),
    .A2(to_WB2_input[2]),
    .A3(to_WB2_input[3]),
    .S0(ConfigBits[12+0]),
    .S0N(ConfigBits_N[12+0]),
    .S1(ConfigBits[12+1]),
    .S1N(ConfigBits_N[12+1]),
    .X(to_WB2)
);

 //switch matrix multiplexer to_WB3 MUX-4
assign to_WB3_input = {from_SB3,from_NB3,from_WB_1s1,from_EB3};
cus_mux41_buf inst_cus_mux41_buf_to_WB3 (
    .A0(to_WB3_input[0]),
    .A1(to_WB3_input[1]),
    .A2(to_WB3_input[2]),
    .A3(to_WB3_input[3]),
    .S0(ConfigBits[14+0]),
    .S0N(ConfigBits_N[14+0]),
    .S1(ConfigBits[14+1]),
    .S1N(ConfigBits_N[14+1]),
    .X(to_WB3)
);

 //switch matrix multiplexer to_WC0 MUX-4
assign to_WC0_input = {GND0,from_SC0,from_NC0,from_EC0};
cus_mux41_buf inst_cus_mux41_buf_to_WC0 (
    .A0(to_WC0_input[0]),
    .A1(to_WC0_input[1]),
    .A2(to_WC0_input[2]),
    .A3(to_WC0_input[3]),
    .S0(ConfigBits[16+0]),
    .S0N(ConfigBits_N[16+0]),
    .S1(ConfigBits[16+1]),
    .S1N(ConfigBits_N[16+1]),
    .X(to_WC0)
);

 //switch matrix multiplexer to_WC1 MUX-4
assign to_WC1_input = {VCC0,from_SC1,from_NC1,from_EC1};
cus_mux41_buf inst_cus_mux41_buf_to_WC1 (
    .A0(to_WC1_input[0]),
    .A1(to_WC1_input[1]),
    .A2(to_WC1_input[2]),
    .A3(to_WC1_input[3]),
    .S0(ConfigBits[18+0]),
    .S0N(ConfigBits_N[18+0]),
    .S1(ConfigBits[18+1]),
    .S1N(ConfigBits_N[18+1]),
    .X(to_WC1)
);

 //switch matrix multiplexer to_WC2 MUX-4
assign to_WC2_input = {from_SC2,from_NC2,from_WC_1s0,from_EC2};
cus_mux41_buf inst_cus_mux41_buf_to_WC2 (
    .A0(to_WC2_input[0]),
    .A1(to_WC2_input[1]),
    .A2(to_WC2_input[2]),
    .A3(to_WC2_input[3]),
    .S0(ConfigBits[20+0]),
    .S0N(ConfigBits_N[20+0]),
    .S1(ConfigBits[20+1]),
    .S1N(ConfigBits_N[20+1]),
    .X(to_WC2)
);

 //switch matrix multiplexer to_WC3 MUX-4
assign to_WC3_input = {from_SC3,from_NC3,from_WC_1s1,from_EC3};
cus_mux41_buf inst_cus_mux41_buf_to_WC3 (
    .A0(to_WC3_input[0]),
    .A1(to_WC3_input[1]),
    .A2(to_WC3_input[2]),
    .A3(to_WC3_input[3]),
    .S0(ConfigBits[22+0]),
    .S0N(ConfigBits_N[22+0]),
    .S1(ConfigBits[22+1]),
    .S1N(ConfigBits_N[22+1]),
    .X(to_WC3)
);

 //switch matrix multiplexer to_WD0 MUX-4
assign to_WD0_input = {GND0,from_SD0,from_ND0,from_ED0};
cus_mux41_buf inst_cus_mux41_buf_to_WD0 (
    .A0(to_WD0_input[0]),
    .A1(to_WD0_input[1]),
    .A2(to_WD0_input[2]),
    .A3(to_WD0_input[3]),
    .S0(ConfigBits[24+0]),
    .S0N(ConfigBits_N[24+0]),
    .S1(ConfigBits[24+1]),
    .S1N(ConfigBits_N[24+1]),
    .X(to_WD0)
);

 //switch matrix multiplexer to_WD1 MUX-4
assign to_WD1_input = {VCC0,from_SD1,from_ND1,from_ED1};
cus_mux41_buf inst_cus_mux41_buf_to_WD1 (
    .A0(to_WD1_input[0]),
    .A1(to_WD1_input[1]),
    .A2(to_WD1_input[2]),
    .A3(to_WD1_input[3]),
    .S0(ConfigBits[26+0]),
    .S0N(ConfigBits_N[26+0]),
    .S1(ConfigBits[26+1]),
    .S1N(ConfigBits_N[26+1]),
    .X(to_WD1)
);

 //switch matrix multiplexer to_WD2 MUX-4
assign to_WD2_input = {from_SD2,from_ND2,from_WD_1s0,from_ED2};
cus_mux41_buf inst_cus_mux41_buf_to_WD2 (
    .A0(to_WD2_input[0]),
    .A1(to_WD2_input[1]),
    .A2(to_WD2_input[2]),
    .A3(to_WD2_input[3]),
    .S0(ConfigBits[28+0]),
    .S0N(ConfigBits_N[28+0]),
    .S1(ConfigBits[28+1]),
    .S1N(ConfigBits_N[28+1]),
    .X(to_WD2)
);

 //switch matrix multiplexer to_WD3 MUX-4
assign to_WD3_input = {from_SD3,from_ND3,from_WD_1s1,from_ED3};
cus_mux41_buf inst_cus_mux41_buf_to_WD3 (
    .A0(to_WD3_input[0]),
    .A1(to_WD3_input[1]),
    .A2(to_WD3_input[2]),
    .A3(to_WD3_input[3]),
    .S0(ConfigBits[30+0]),
    .S0N(ConfigBits_N[30+0]),
    .S1(ConfigBits[30+1]),
    .S1N(ConfigBits_N[30+1]),
    .X(to_WD3)
);

 //switch matrix multiplexer to_WF0 MUX-4
assign to_WF0_input = {GND0,from_SF0,from_NF0,from_EF0};
cus_mux41_buf inst_cus_mux41_buf_to_WF0 (
    .A0(to_WF0_input[0]),
    .A1(to_WF0_input[1]),
    .A2(to_WF0_input[2]),
    .A3(to_WF0_input[3]),
    .S0(ConfigBits[32+0]),
    .S0N(ConfigBits_N[32+0]),
    .S1(ConfigBits[32+1]),
    .S1N(ConfigBits_N[32+1]),
    .X(to_WF0)
);

 //switch matrix multiplexer to_WF1 MUX-4
assign to_WF1_input = {VCC0,from_SF1,from_NF1,from_EF1};
cus_mux41_buf inst_cus_mux41_buf_to_WF1 (
    .A0(to_WF1_input[0]),
    .A1(to_WF1_input[1]),
    .A2(to_WF1_input[2]),
    .A3(to_WF1_input[3]),
    .S0(ConfigBits[34+0]),
    .S0N(ConfigBits_N[34+0]),
    .S1(ConfigBits[34+1]),
    .S1N(ConfigBits_N[34+1]),
    .X(to_WF1)
);

 //switch matrix multiplexer to_WF2 MUX-4
assign to_WF2_input = {from_SF2,from_NF2,from_WF_1s0,from_EF2};
cus_mux41_buf inst_cus_mux41_buf_to_WF2 (
    .A0(to_WF2_input[0]),
    .A1(to_WF2_input[1]),
    .A2(to_WF2_input[2]),
    .A3(to_WF2_input[3]),
    .S0(ConfigBits[36+0]),
    .S0N(ConfigBits_N[36+0]),
    .S1(ConfigBits[36+1]),
    .S1N(ConfigBits_N[36+1]),
    .X(to_WF2)
);

 //switch matrix multiplexer to_WF3 MUX-4
assign to_WF3_input = {from_SF3,from_NF3,from_WF_1s1,from_EF3};
cus_mux41_buf inst_cus_mux41_buf_to_WF3 (
    .A0(to_WF3_input[0]),
    .A1(to_WF3_input[1]),
    .A2(to_WF3_input[2]),
    .A3(to_WF3_input[3]),
    .S0(ConfigBits[38+0]),
    .S0N(ConfigBits_N[38+0]),
    .S1(ConfigBits[38+1]),
    .S1N(ConfigBits_N[38+1]),
    .X(to_WF3)
);

 //switch matrix multiplexer to_WG0 MUX-4
assign to_WG0_input = {GND0,from_SG0,from_NG0,from_EG0};
cus_mux41_buf inst_cus_mux41_buf_to_WG0 (
    .A0(to_WG0_input[0]),
    .A1(to_WG0_input[1]),
    .A2(to_WG0_input[2]),
    .A3(to_WG0_input[3]),
    .S0(ConfigBits[40+0]),
    .S0N(ConfigBits_N[40+0]),
    .S1(ConfigBits[40+1]),
    .S1N(ConfigBits_N[40+1]),
    .X(to_WG0)
);

 //switch matrix multiplexer to_WG1 MUX-4
assign to_WG1_input = {VCC0,from_SG1,from_NG1,from_EG1};
cus_mux41_buf inst_cus_mux41_buf_to_WG1 (
    .A0(to_WG1_input[0]),
    .A1(to_WG1_input[1]),
    .A2(to_WG1_input[2]),
    .A3(to_WG1_input[3]),
    .S0(ConfigBits[42+0]),
    .S0N(ConfigBits_N[42+0]),
    .S1(ConfigBits[42+1]),
    .S1N(ConfigBits_N[42+1]),
    .X(to_WG1)
);

 //switch matrix multiplexer to_WG2 MUX-4
assign to_WG2_input = {from_SG2,from_NG2,from_WG_1s0,from_EG2};
cus_mux41_buf inst_cus_mux41_buf_to_WG2 (
    .A0(to_WG2_input[0]),
    .A1(to_WG2_input[1]),
    .A2(to_WG2_input[2]),
    .A3(to_WG2_input[3]),
    .S0(ConfigBits[44+0]),
    .S0N(ConfigBits_N[44+0]),
    .S1(ConfigBits[44+1]),
    .S1N(ConfigBits_N[44+1]),
    .X(to_WG2)
);

 //switch matrix multiplexer to_WG3 MUX-4
assign to_WG3_input = {from_SG3,from_NG3,from_WG_1s1,from_EG3};
cus_mux41_buf inst_cus_mux41_buf_to_WG3 (
    .A0(to_WG3_input[0]),
    .A1(to_WG3_input[1]),
    .A2(to_WG3_input[2]),
    .A3(to_WG3_input[3]),
    .S0(ConfigBits[46+0]),
    .S0N(ConfigBits_N[46+0]),
    .S1(ConfigBits[46+1]),
    .S1N(ConfigBits_N[46+1]),
    .X(to_WG3)
);

 //switch matrix multiplexer to_WG4 MUX-1
assign to_WG4 = from_EG4;

 //switch matrix multiplexer to_WG5 MUX-1
assign to_WG5 = from_EG5;

 //switch matrix multiplexer to_WG6 MUX-1
assign to_WG6 = from_EG6;

 //switch matrix multiplexer to_WG7 MUX-1
assign to_WG7 = from_EG7;

 //switch matrix multiplexer to_WH0 MUX-4
assign to_WH0_input = {GND0,from_SH0,from_NH0,from_EH0};
cus_mux41_buf inst_cus_mux41_buf_to_WH0 (
    .A0(to_WH0_input[0]),
    .A1(to_WH0_input[1]),
    .A2(to_WH0_input[2]),
    .A3(to_WH0_input[3]),
    .S0(ConfigBits[48+0]),
    .S0N(ConfigBits_N[48+0]),
    .S1(ConfigBits[48+1]),
    .S1N(ConfigBits_N[48+1]),
    .X(to_WH0)
);

 //switch matrix multiplexer to_WH1 MUX-4
assign to_WH1_input = {VCC0,from_SH1,from_NH1,from_EH1};
cus_mux41_buf inst_cus_mux41_buf_to_WH1 (
    .A0(to_WH1_input[0]),
    .A1(to_WH1_input[1]),
    .A2(to_WH1_input[2]),
    .A3(to_WH1_input[3]),
    .S0(ConfigBits[50+0]),
    .S0N(ConfigBits_N[50+0]),
    .S1(ConfigBits[50+1]),
    .S1N(ConfigBits_N[50+1]),
    .X(to_WH1)
);

 //switch matrix multiplexer to_WH2 MUX-4
assign to_WH2_input = {from_SH2,from_NH2,from_WH_1s0,from_EH2};
cus_mux41_buf inst_cus_mux41_buf_to_WH2 (
    .A0(to_WH2_input[0]),
    .A1(to_WH2_input[1]),
    .A2(to_WH2_input[2]),
    .A3(to_WH2_input[3]),
    .S0(ConfigBits[52+0]),
    .S0N(ConfigBits_N[52+0]),
    .S1(ConfigBits[52+1]),
    .S1N(ConfigBits_N[52+1]),
    .X(to_WH2)
);

 //switch matrix multiplexer to_WH3 MUX-4
assign to_WH3_input = {from_SH3,from_NH3,from_WH_1s1,from_EH3};
cus_mux41_buf inst_cus_mux41_buf_to_WH3 (
    .A0(to_WH3_input[0]),
    .A1(to_WH3_input[1]),
    .A2(to_WH3_input[2]),
    .A3(to_WH3_input[3]),
    .S0(ConfigBits[54+0]),
    .S0N(ConfigBits_N[54+0]),
    .S1(ConfigBits[54+1]),
    .S1N(ConfigBits_N[54+1]),
    .X(to_WH3)
);

 //switch matrix multiplexer to_WH4 MUX-1
assign to_WH4 = from_EH4;

 //switch matrix multiplexer to_WH5 MUX-1
assign to_WH5 = from_EH5;

 //switch matrix multiplexer to_WH6 MUX-1
assign to_WH6 = from_EH6;

 //switch matrix multiplexer to_WH7 MUX-1
assign to_WH7 = from_EH7;

 //switch matrix multiplexer to_WI0 MUX-4
assign to_WI0_input = {GND0,from_SI0,from_NI0,from_EI0};
cus_mux41_buf inst_cus_mux41_buf_to_WI0 (
    .A0(to_WI0_input[0]),
    .A1(to_WI0_input[1]),
    .A2(to_WI0_input[2]),
    .A3(to_WI0_input[3]),
    .S0(ConfigBits[56+0]),
    .S0N(ConfigBits_N[56+0]),
    .S1(ConfigBits[56+1]),
    .S1N(ConfigBits_N[56+1]),
    .X(to_WI0)
);

 //switch matrix multiplexer to_WI1 MUX-4
assign to_WI1_input = {VCC0,from_SI1,from_NI1,from_EI1};
cus_mux41_buf inst_cus_mux41_buf_to_WI1 (
    .A0(to_WI1_input[0]),
    .A1(to_WI1_input[1]),
    .A2(to_WI1_input[2]),
    .A3(to_WI1_input[3]),
    .S0(ConfigBits[58+0]),
    .S0N(ConfigBits_N[58+0]),
    .S1(ConfigBits[58+1]),
    .S1N(ConfigBits_N[58+1]),
    .X(to_WI1)
);

 //switch matrix multiplexer to_WI2 MUX-4
assign to_WI2_input = {from_SI2,from_NI2,from_WI_1s0,from_EI2};
cus_mux41_buf inst_cus_mux41_buf_to_WI2 (
    .A0(to_WI2_input[0]),
    .A1(to_WI2_input[1]),
    .A2(to_WI2_input[2]),
    .A3(to_WI2_input[3]),
    .S0(ConfigBits[60+0]),
    .S0N(ConfigBits_N[60+0]),
    .S1(ConfigBits[60+1]),
    .S1N(ConfigBits_N[60+1]),
    .X(to_WI2)
);

 //switch matrix multiplexer to_WI3 MUX-4
assign to_WI3_input = {from_SI3,from_NI3,from_WI_1s1,from_EI3};
cus_mux41_buf inst_cus_mux41_buf_to_WI3 (
    .A0(to_WI3_input[0]),
    .A1(to_WI3_input[1]),
    .A2(to_WI3_input[2]),
    .A3(to_WI3_input[3]),
    .S0(ConfigBits[62+0]),
    .S0N(ConfigBits_N[62+0]),
    .S1(ConfigBits[62+1]),
    .S1N(ConfigBits_N[62+1]),
    .X(to_WI3)
);

 //switch matrix multiplexer to_WI4 MUX-1
assign to_WI4 = from_EI4;

 //switch matrix multiplexer to_WI5 MUX-1
assign to_WI5 = from_EI5;

 //switch matrix multiplexer to_WI6 MUX-1
assign to_WI6 = from_EI6;

 //switch matrix multiplexer to_WI7 MUX-1
assign to_WI7 = from_EI7;

 //switch matrix multiplexer to_WI8 MUX-1
assign to_WI8 = from_EI8;

 //switch matrix multiplexer to_WI9 MUX-1
assign to_WI9 = from_EI9;

 //switch matrix multiplexer to_WI10 MUX-1
assign to_WI10 = from_EI10;

 //switch matrix multiplexer to_WI11 MUX-1
assign to_WI11 = from_EI11;

 //switch matrix multiplexer to_NA0 MUX-4
assign to_NA0_input = {GND0,from_SA0,from_NA0,from_EA0};
cus_mux41_buf inst_cus_mux41_buf_to_NA0 (
    .A0(to_NA0_input[0]),
    .A1(to_NA0_input[1]),
    .A2(to_NA0_input[2]),
    .A3(to_NA0_input[3]),
    .S0(ConfigBits[64+0]),
    .S0N(ConfigBits_N[64+0]),
    .S1(ConfigBits[64+1]),
    .S1N(ConfigBits_N[64+1]),
    .X(to_NA0)
);

 //switch matrix multiplexer to_NA1 MUX-4
assign to_NA1_input = {VCC0,from_SA1,from_NA1,from_EA1};
cus_mux41_buf inst_cus_mux41_buf_to_NA1 (
    .A0(to_NA1_input[0]),
    .A1(to_NA1_input[1]),
    .A2(to_NA1_input[2]),
    .A3(to_NA1_input[3]),
    .S0(ConfigBits[66+0]),
    .S0N(ConfigBits_N[66+0]),
    .S1(ConfigBits[66+1]),
    .S1N(ConfigBits_N[66+1]),
    .X(to_NA1)
);

 //switch matrix multiplexer to_NA2 MUX-4
assign to_NA2_input = {from_SA2,from_NA2,from_WA_1s0,from_EA2};
cus_mux41_buf inst_cus_mux41_buf_to_NA2 (
    .A0(to_NA2_input[0]),
    .A1(to_NA2_input[1]),
    .A2(to_NA2_input[2]),
    .A3(to_NA2_input[3]),
    .S0(ConfigBits[68+0]),
    .S0N(ConfigBits_N[68+0]),
    .S1(ConfigBits[68+1]),
    .S1N(ConfigBits_N[68+1]),
    .X(to_NA2)
);

 //switch matrix multiplexer to_NA3 MUX-4
assign to_NA3_input = {from_SA3,from_NA3,from_WA_1s1,from_EA3};
cus_mux41_buf inst_cus_mux41_buf_to_NA3 (
    .A0(to_NA3_input[0]),
    .A1(to_NA3_input[1]),
    .A2(to_NA3_input[2]),
    .A3(to_NA3_input[3]),
    .S0(ConfigBits[70+0]),
    .S0N(ConfigBits_N[70+0]),
    .S1(ConfigBits[70+1]),
    .S1N(ConfigBits_N[70+1]),
    .X(to_NA3)
);

 //switch matrix multiplexer to_NB0 MUX-4
assign to_NB0_input = {GND0,from_SB0,from_NB0,from_EB0};
cus_mux41_buf inst_cus_mux41_buf_to_NB0 (
    .A0(to_NB0_input[0]),
    .A1(to_NB0_input[1]),
    .A2(to_NB0_input[2]),
    .A3(to_NB0_input[3]),
    .S0(ConfigBits[72+0]),
    .S0N(ConfigBits_N[72+0]),
    .S1(ConfigBits[72+1]),
    .S1N(ConfigBits_N[72+1]),
    .X(to_NB0)
);

 //switch matrix multiplexer to_NB1 MUX-4
assign to_NB1_input = {VCC0,from_SB1,from_NB1,from_EB1};
cus_mux41_buf inst_cus_mux41_buf_to_NB1 (
    .A0(to_NB1_input[0]),
    .A1(to_NB1_input[1]),
    .A2(to_NB1_input[2]),
    .A3(to_NB1_input[3]),
    .S0(ConfigBits[74+0]),
    .S0N(ConfigBits_N[74+0]),
    .S1(ConfigBits[74+1]),
    .S1N(ConfigBits_N[74+1]),
    .X(to_NB1)
);

 //switch matrix multiplexer to_NB2 MUX-4
assign to_NB2_input = {from_SB2,from_NB2,from_WB_1s0,from_EB2};
cus_mux41_buf inst_cus_mux41_buf_to_NB2 (
    .A0(to_NB2_input[0]),
    .A1(to_NB2_input[1]),
    .A2(to_NB2_input[2]),
    .A3(to_NB2_input[3]),
    .S0(ConfigBits[76+0]),
    .S0N(ConfigBits_N[76+0]),
    .S1(ConfigBits[76+1]),
    .S1N(ConfigBits_N[76+1]),
    .X(to_NB2)
);

 //switch matrix multiplexer to_NB3 MUX-4
assign to_NB3_input = {from_SB3,from_NB3,from_WB_1s1,from_EB3};
cus_mux41_buf inst_cus_mux41_buf_to_NB3 (
    .A0(to_NB3_input[0]),
    .A1(to_NB3_input[1]),
    .A2(to_NB3_input[2]),
    .A3(to_NB3_input[3]),
    .S0(ConfigBits[78+0]),
    .S0N(ConfigBits_N[78+0]),
    .S1(ConfigBits[78+1]),
    .S1N(ConfigBits_N[78+1]),
    .X(to_NB3)
);

 //switch matrix multiplexer to_NC0 MUX-4
assign to_NC0_input = {GND0,from_SC0,from_NC0,from_EC0};
cus_mux41_buf inst_cus_mux41_buf_to_NC0 (
    .A0(to_NC0_input[0]),
    .A1(to_NC0_input[1]),
    .A2(to_NC0_input[2]),
    .A3(to_NC0_input[3]),
    .S0(ConfigBits[80+0]),
    .S0N(ConfigBits_N[80+0]),
    .S1(ConfigBits[80+1]),
    .S1N(ConfigBits_N[80+1]),
    .X(to_NC0)
);

 //switch matrix multiplexer to_NC1 MUX-4
assign to_NC1_input = {VCC0,from_SC1,from_NC1,from_EC1};
cus_mux41_buf inst_cus_mux41_buf_to_NC1 (
    .A0(to_NC1_input[0]),
    .A1(to_NC1_input[1]),
    .A2(to_NC1_input[2]),
    .A3(to_NC1_input[3]),
    .S0(ConfigBits[82+0]),
    .S0N(ConfigBits_N[82+0]),
    .S1(ConfigBits[82+1]),
    .S1N(ConfigBits_N[82+1]),
    .X(to_NC1)
);

 //switch matrix multiplexer to_NC2 MUX-4
assign to_NC2_input = {from_SC2,from_NC2,from_WC_1s0,from_EC2};
cus_mux41_buf inst_cus_mux41_buf_to_NC2 (
    .A0(to_NC2_input[0]),
    .A1(to_NC2_input[1]),
    .A2(to_NC2_input[2]),
    .A3(to_NC2_input[3]),
    .S0(ConfigBits[84+0]),
    .S0N(ConfigBits_N[84+0]),
    .S1(ConfigBits[84+1]),
    .S1N(ConfigBits_N[84+1]),
    .X(to_NC2)
);

 //switch matrix multiplexer to_NC3 MUX-4
assign to_NC3_input = {from_SC3,from_NC3,from_WC_1s1,from_EC3};
cus_mux41_buf inst_cus_mux41_buf_to_NC3 (
    .A0(to_NC3_input[0]),
    .A1(to_NC3_input[1]),
    .A2(to_NC3_input[2]),
    .A3(to_NC3_input[3]),
    .S0(ConfigBits[86+0]),
    .S0N(ConfigBits_N[86+0]),
    .S1(ConfigBits[86+1]),
    .S1N(ConfigBits_N[86+1]),
    .X(to_NC3)
);

 //switch matrix multiplexer to_ND0 MUX-4
assign to_ND0_input = {GND0,from_SD0,from_ND0,from_ED0};
cus_mux41_buf inst_cus_mux41_buf_to_ND0 (
    .A0(to_ND0_input[0]),
    .A1(to_ND0_input[1]),
    .A2(to_ND0_input[2]),
    .A3(to_ND0_input[3]),
    .S0(ConfigBits[88+0]),
    .S0N(ConfigBits_N[88+0]),
    .S1(ConfigBits[88+1]),
    .S1N(ConfigBits_N[88+1]),
    .X(to_ND0)
);

 //switch matrix multiplexer to_ND1 MUX-4
assign to_ND1_input = {VCC0,from_SD1,from_ND1,from_ED1};
cus_mux41_buf inst_cus_mux41_buf_to_ND1 (
    .A0(to_ND1_input[0]),
    .A1(to_ND1_input[1]),
    .A2(to_ND1_input[2]),
    .A3(to_ND1_input[3]),
    .S0(ConfigBits[90+0]),
    .S0N(ConfigBits_N[90+0]),
    .S1(ConfigBits[90+1]),
    .S1N(ConfigBits_N[90+1]),
    .X(to_ND1)
);

 //switch matrix multiplexer to_ND2 MUX-4
assign to_ND2_input = {from_SD2,from_ND2,from_WD_1s0,from_ED2};
cus_mux41_buf inst_cus_mux41_buf_to_ND2 (
    .A0(to_ND2_input[0]),
    .A1(to_ND2_input[1]),
    .A2(to_ND2_input[2]),
    .A3(to_ND2_input[3]),
    .S0(ConfigBits[92+0]),
    .S0N(ConfigBits_N[92+0]),
    .S1(ConfigBits[92+1]),
    .S1N(ConfigBits_N[92+1]),
    .X(to_ND2)
);

 //switch matrix multiplexer to_ND3 MUX-4
assign to_ND3_input = {from_SD3,from_ND3,from_WD_1s1,from_ED3};
cus_mux41_buf inst_cus_mux41_buf_to_ND3 (
    .A0(to_ND3_input[0]),
    .A1(to_ND3_input[1]),
    .A2(to_ND3_input[2]),
    .A3(to_ND3_input[3]),
    .S0(ConfigBits[94+0]),
    .S0N(ConfigBits_N[94+0]),
    .S1(ConfigBits[94+1]),
    .S1N(ConfigBits_N[94+1]),
    .X(to_ND3)
);

 //switch matrix multiplexer to_NF0 MUX-4
assign to_NF0_input = {GND0,from_SF0,from_NF0,from_EF0};
cus_mux41_buf inst_cus_mux41_buf_to_NF0 (
    .A0(to_NF0_input[0]),
    .A1(to_NF0_input[1]),
    .A2(to_NF0_input[2]),
    .A3(to_NF0_input[3]),
    .S0(ConfigBits[96+0]),
    .S0N(ConfigBits_N[96+0]),
    .S1(ConfigBits[96+1]),
    .S1N(ConfigBits_N[96+1]),
    .X(to_NF0)
);

 //switch matrix multiplexer to_NF1 MUX-4
assign to_NF1_input = {VCC0,from_SF1,from_NF1,from_EF1};
cus_mux41_buf inst_cus_mux41_buf_to_NF1 (
    .A0(to_NF1_input[0]),
    .A1(to_NF1_input[1]),
    .A2(to_NF1_input[2]),
    .A3(to_NF1_input[3]),
    .S0(ConfigBits[98+0]),
    .S0N(ConfigBits_N[98+0]),
    .S1(ConfigBits[98+1]),
    .S1N(ConfigBits_N[98+1]),
    .X(to_NF1)
);

 //switch matrix multiplexer to_NF2 MUX-4
assign to_NF2_input = {from_SF2,from_NF2,from_WF_1s0,from_EF2};
cus_mux41_buf inst_cus_mux41_buf_to_NF2 (
    .A0(to_NF2_input[0]),
    .A1(to_NF2_input[1]),
    .A2(to_NF2_input[2]),
    .A3(to_NF2_input[3]),
    .S0(ConfigBits[100+0]),
    .S0N(ConfigBits_N[100+0]),
    .S1(ConfigBits[100+1]),
    .S1N(ConfigBits_N[100+1]),
    .X(to_NF2)
);

 //switch matrix multiplexer to_NF3 MUX-4
assign to_NF3_input = {from_SF3,from_NF3,from_WF_1s1,from_EF3};
cus_mux41_buf inst_cus_mux41_buf_to_NF3 (
    .A0(to_NF3_input[0]),
    .A1(to_NF3_input[1]),
    .A2(to_NF3_input[2]),
    .A3(to_NF3_input[3]),
    .S0(ConfigBits[102+0]),
    .S0N(ConfigBits_N[102+0]),
    .S1(ConfigBits[102+1]),
    .S1N(ConfigBits_N[102+1]),
    .X(to_NF3)
);

 //switch matrix multiplexer to_NG0 MUX-4
assign to_NG0_input = {GND0,from_SG0,from_NG0,from_EG0};
cus_mux41_buf inst_cus_mux41_buf_to_NG0 (
    .A0(to_NG0_input[0]),
    .A1(to_NG0_input[1]),
    .A2(to_NG0_input[2]),
    .A3(to_NG0_input[3]),
    .S0(ConfigBits[104+0]),
    .S0N(ConfigBits_N[104+0]),
    .S1(ConfigBits[104+1]),
    .S1N(ConfigBits_N[104+1]),
    .X(to_NG0)
);

 //switch matrix multiplexer to_NG1 MUX-4
assign to_NG1_input = {VCC0,from_SG1,from_NG1,from_EG1};
cus_mux41_buf inst_cus_mux41_buf_to_NG1 (
    .A0(to_NG1_input[0]),
    .A1(to_NG1_input[1]),
    .A2(to_NG1_input[2]),
    .A3(to_NG1_input[3]),
    .S0(ConfigBits[106+0]),
    .S0N(ConfigBits_N[106+0]),
    .S1(ConfigBits[106+1]),
    .S1N(ConfigBits_N[106+1]),
    .X(to_NG1)
);

 //switch matrix multiplexer to_NG2 MUX-4
assign to_NG2_input = {from_SG2,from_NG2,from_WG_1s0,from_EG2};
cus_mux41_buf inst_cus_mux41_buf_to_NG2 (
    .A0(to_NG2_input[0]),
    .A1(to_NG2_input[1]),
    .A2(to_NG2_input[2]),
    .A3(to_NG2_input[3]),
    .S0(ConfigBits[108+0]),
    .S0N(ConfigBits_N[108+0]),
    .S1(ConfigBits[108+1]),
    .S1N(ConfigBits_N[108+1]),
    .X(to_NG2)
);

 //switch matrix multiplexer to_NG3 MUX-4
assign to_NG3_input = {from_SG3,from_NG3,from_WG_1s1,from_EG3};
cus_mux41_buf inst_cus_mux41_buf_to_NG3 (
    .A0(to_NG3_input[0]),
    .A1(to_NG3_input[1]),
    .A2(to_NG3_input[2]),
    .A3(to_NG3_input[3]),
    .S0(ConfigBits[110+0]),
    .S0N(ConfigBits_N[110+0]),
    .S1(ConfigBits[110+1]),
    .S1N(ConfigBits_N[110+1]),
    .X(to_NG3)
);

 //switch matrix multiplexer to_NH0 MUX-4
assign to_NH0_input = {GND0,from_SH0,from_NH0,from_EH0};
cus_mux41_buf inst_cus_mux41_buf_to_NH0 (
    .A0(to_NH0_input[0]),
    .A1(to_NH0_input[1]),
    .A2(to_NH0_input[2]),
    .A3(to_NH0_input[3]),
    .S0(ConfigBits[112+0]),
    .S0N(ConfigBits_N[112+0]),
    .S1(ConfigBits[112+1]),
    .S1N(ConfigBits_N[112+1]),
    .X(to_NH0)
);

 //switch matrix multiplexer to_NH1 MUX-4
assign to_NH1_input = {VCC0,from_SH1,from_NH1,from_EH1};
cus_mux41_buf inst_cus_mux41_buf_to_NH1 (
    .A0(to_NH1_input[0]),
    .A1(to_NH1_input[1]),
    .A2(to_NH1_input[2]),
    .A3(to_NH1_input[3]),
    .S0(ConfigBits[114+0]),
    .S0N(ConfigBits_N[114+0]),
    .S1(ConfigBits[114+1]),
    .S1N(ConfigBits_N[114+1]),
    .X(to_NH1)
);

 //switch matrix multiplexer to_NH2 MUX-4
assign to_NH2_input = {from_SH2,from_NH2,from_WH_1s0,from_EH2};
cus_mux41_buf inst_cus_mux41_buf_to_NH2 (
    .A0(to_NH2_input[0]),
    .A1(to_NH2_input[1]),
    .A2(to_NH2_input[2]),
    .A3(to_NH2_input[3]),
    .S0(ConfigBits[116+0]),
    .S0N(ConfigBits_N[116+0]),
    .S1(ConfigBits[116+1]),
    .S1N(ConfigBits_N[116+1]),
    .X(to_NH2)
);

 //switch matrix multiplexer to_NH3 MUX-4
assign to_NH3_input = {from_SH3,from_NH3,from_WH_1s1,from_EH3};
cus_mux41_buf inst_cus_mux41_buf_to_NH3 (
    .A0(to_NH3_input[0]),
    .A1(to_NH3_input[1]),
    .A2(to_NH3_input[2]),
    .A3(to_NH3_input[3]),
    .S0(ConfigBits[118+0]),
    .S0N(ConfigBits_N[118+0]),
    .S1(ConfigBits[118+1]),
    .S1N(ConfigBits_N[118+1]),
    .X(to_NH3)
);

 //switch matrix multiplexer to_NI0 MUX-4
assign to_NI0_input = {GND0,from_SI0,from_NI0,from_EI0};
cus_mux41_buf inst_cus_mux41_buf_to_NI0 (
    .A0(to_NI0_input[0]),
    .A1(to_NI0_input[1]),
    .A2(to_NI0_input[2]),
    .A3(to_NI0_input[3]),
    .S0(ConfigBits[120+0]),
    .S0N(ConfigBits_N[120+0]),
    .S1(ConfigBits[120+1]),
    .S1N(ConfigBits_N[120+1]),
    .X(to_NI0)
);

 //switch matrix multiplexer to_NI1 MUX-4
assign to_NI1_input = {VCC0,from_SI1,from_NI1,from_EI1};
cus_mux41_buf inst_cus_mux41_buf_to_NI1 (
    .A0(to_NI1_input[0]),
    .A1(to_NI1_input[1]),
    .A2(to_NI1_input[2]),
    .A3(to_NI1_input[3]),
    .S0(ConfigBits[122+0]),
    .S0N(ConfigBits_N[122+0]),
    .S1(ConfigBits[122+1]),
    .S1N(ConfigBits_N[122+1]),
    .X(to_NI1)
);

 //switch matrix multiplexer to_NI2 MUX-4
assign to_NI2_input = {from_SI2,from_NI2,from_WI_1s0,from_EI2};
cus_mux41_buf inst_cus_mux41_buf_to_NI2 (
    .A0(to_NI2_input[0]),
    .A1(to_NI2_input[1]),
    .A2(to_NI2_input[2]),
    .A3(to_NI2_input[3]),
    .S0(ConfigBits[124+0]),
    .S0N(ConfigBits_N[124+0]),
    .S1(ConfigBits[124+1]),
    .S1N(ConfigBits_N[124+1]),
    .X(to_NI2)
);

 //switch matrix multiplexer to_NI3 MUX-4
assign to_NI3_input = {from_SI3,from_NI3,from_WI_1s1,from_EI3};
cus_mux41_buf inst_cus_mux41_buf_to_NI3 (
    .A0(to_NI3_input[0]),
    .A1(to_NI3_input[1]),
    .A2(to_NI3_input[2]),
    .A3(to_NI3_input[3]),
    .S0(ConfigBits[126+0]),
    .S0N(ConfigBits_N[126+0]),
    .S1(ConfigBits[126+1]),
    .S1N(ConfigBits_N[126+1]),
    .X(to_NI3)
);

 //switch matrix multiplexer to_SA0 MUX-4
assign to_SA0_input = {GND0,from_SA0,from_NA0,from_EA0};
cus_mux41_buf inst_cus_mux41_buf_to_SA0 (
    .A0(to_SA0_input[0]),
    .A1(to_SA0_input[1]),
    .A2(to_SA0_input[2]),
    .A3(to_SA0_input[3]),
    .S0(ConfigBits[128+0]),
    .S0N(ConfigBits_N[128+0]),
    .S1(ConfigBits[128+1]),
    .S1N(ConfigBits_N[128+1]),
    .X(to_SA0)
);

 //switch matrix multiplexer to_SA1 MUX-4
assign to_SA1_input = {VCC0,from_SA1,from_NA1,from_EA1};
cus_mux41_buf inst_cus_mux41_buf_to_SA1 (
    .A0(to_SA1_input[0]),
    .A1(to_SA1_input[1]),
    .A2(to_SA1_input[2]),
    .A3(to_SA1_input[3]),
    .S0(ConfigBits[130+0]),
    .S0N(ConfigBits_N[130+0]),
    .S1(ConfigBits[130+1]),
    .S1N(ConfigBits_N[130+1]),
    .X(to_SA1)
);

 //switch matrix multiplexer to_SA2 MUX-4
assign to_SA2_input = {from_SA2,from_NA2,from_WA_1s0,from_EA2};
cus_mux41_buf inst_cus_mux41_buf_to_SA2 (
    .A0(to_SA2_input[0]),
    .A1(to_SA2_input[1]),
    .A2(to_SA2_input[2]),
    .A3(to_SA2_input[3]),
    .S0(ConfigBits[132+0]),
    .S0N(ConfigBits_N[132+0]),
    .S1(ConfigBits[132+1]),
    .S1N(ConfigBits_N[132+1]),
    .X(to_SA2)
);

 //switch matrix multiplexer to_SA3 MUX-4
assign to_SA3_input = {from_SA3,from_NA3,from_WA_1s1,from_EA3};
cus_mux41_buf inst_cus_mux41_buf_to_SA3 (
    .A0(to_SA3_input[0]),
    .A1(to_SA3_input[1]),
    .A2(to_SA3_input[2]),
    .A3(to_SA3_input[3]),
    .S0(ConfigBits[134+0]),
    .S0N(ConfigBits_N[134+0]),
    .S1(ConfigBits[134+1]),
    .S1N(ConfigBits_N[134+1]),
    .X(to_SA3)
);

 //switch matrix multiplexer to_SB0 MUX-4
assign to_SB0_input = {GND0,from_SB0,from_NB0,from_EB0};
cus_mux41_buf inst_cus_mux41_buf_to_SB0 (
    .A0(to_SB0_input[0]),
    .A1(to_SB0_input[1]),
    .A2(to_SB0_input[2]),
    .A3(to_SB0_input[3]),
    .S0(ConfigBits[136+0]),
    .S0N(ConfigBits_N[136+0]),
    .S1(ConfigBits[136+1]),
    .S1N(ConfigBits_N[136+1]),
    .X(to_SB0)
);

 //switch matrix multiplexer to_SB1 MUX-4
assign to_SB1_input = {VCC0,from_SB1,from_NB1,from_EB1};
cus_mux41_buf inst_cus_mux41_buf_to_SB1 (
    .A0(to_SB1_input[0]),
    .A1(to_SB1_input[1]),
    .A2(to_SB1_input[2]),
    .A3(to_SB1_input[3]),
    .S0(ConfigBits[138+0]),
    .S0N(ConfigBits_N[138+0]),
    .S1(ConfigBits[138+1]),
    .S1N(ConfigBits_N[138+1]),
    .X(to_SB1)
);

 //switch matrix multiplexer to_SB2 MUX-4
assign to_SB2_input = {from_SB2,from_NB2,from_WB_1s0,from_EB2};
cus_mux41_buf inst_cus_mux41_buf_to_SB2 (
    .A0(to_SB2_input[0]),
    .A1(to_SB2_input[1]),
    .A2(to_SB2_input[2]),
    .A3(to_SB2_input[3]),
    .S0(ConfigBits[140+0]),
    .S0N(ConfigBits_N[140+0]),
    .S1(ConfigBits[140+1]),
    .S1N(ConfigBits_N[140+1]),
    .X(to_SB2)
);

 //switch matrix multiplexer to_SB3 MUX-4
assign to_SB3_input = {from_SB3,from_NB3,from_WB_1s1,from_EB3};
cus_mux41_buf inst_cus_mux41_buf_to_SB3 (
    .A0(to_SB3_input[0]),
    .A1(to_SB3_input[1]),
    .A2(to_SB3_input[2]),
    .A3(to_SB3_input[3]),
    .S0(ConfigBits[142+0]),
    .S0N(ConfigBits_N[142+0]),
    .S1(ConfigBits[142+1]),
    .S1N(ConfigBits_N[142+1]),
    .X(to_SB3)
);

 //switch matrix multiplexer to_SC0 MUX-4
assign to_SC0_input = {GND0,from_SC0,from_NC0,from_EC0};
cus_mux41_buf inst_cus_mux41_buf_to_SC0 (
    .A0(to_SC0_input[0]),
    .A1(to_SC0_input[1]),
    .A2(to_SC0_input[2]),
    .A3(to_SC0_input[3]),
    .S0(ConfigBits[144+0]),
    .S0N(ConfigBits_N[144+0]),
    .S1(ConfigBits[144+1]),
    .S1N(ConfigBits_N[144+1]),
    .X(to_SC0)
);

 //switch matrix multiplexer to_SC1 MUX-4
assign to_SC1_input = {VCC0,from_SC1,from_NC1,from_EC1};
cus_mux41_buf inst_cus_mux41_buf_to_SC1 (
    .A0(to_SC1_input[0]),
    .A1(to_SC1_input[1]),
    .A2(to_SC1_input[2]),
    .A3(to_SC1_input[3]),
    .S0(ConfigBits[146+0]),
    .S0N(ConfigBits_N[146+0]),
    .S1(ConfigBits[146+1]),
    .S1N(ConfigBits_N[146+1]),
    .X(to_SC1)
);

 //switch matrix multiplexer to_SC2 MUX-4
assign to_SC2_input = {from_SC2,from_NC2,from_WC_1s0,from_EC2};
cus_mux41_buf inst_cus_mux41_buf_to_SC2 (
    .A0(to_SC2_input[0]),
    .A1(to_SC2_input[1]),
    .A2(to_SC2_input[2]),
    .A3(to_SC2_input[3]),
    .S0(ConfigBits[148+0]),
    .S0N(ConfigBits_N[148+0]),
    .S1(ConfigBits[148+1]),
    .S1N(ConfigBits_N[148+1]),
    .X(to_SC2)
);

 //switch matrix multiplexer to_SC3 MUX-4
assign to_SC3_input = {from_SC3,from_NC3,from_WC_1s1,from_EC3};
cus_mux41_buf inst_cus_mux41_buf_to_SC3 (
    .A0(to_SC3_input[0]),
    .A1(to_SC3_input[1]),
    .A2(to_SC3_input[2]),
    .A3(to_SC3_input[3]),
    .S0(ConfigBits[150+0]),
    .S0N(ConfigBits_N[150+0]),
    .S1(ConfigBits[150+1]),
    .S1N(ConfigBits_N[150+1]),
    .X(to_SC3)
);

 //switch matrix multiplexer to_SD0 MUX-4
assign to_SD0_input = {GND0,from_SD0,from_ND0,from_ED0};
cus_mux41_buf inst_cus_mux41_buf_to_SD0 (
    .A0(to_SD0_input[0]),
    .A1(to_SD0_input[1]),
    .A2(to_SD0_input[2]),
    .A3(to_SD0_input[3]),
    .S0(ConfigBits[152+0]),
    .S0N(ConfigBits_N[152+0]),
    .S1(ConfigBits[152+1]),
    .S1N(ConfigBits_N[152+1]),
    .X(to_SD0)
);

 //switch matrix multiplexer to_SD1 MUX-4
assign to_SD1_input = {VCC0,from_SD1,from_ND1,from_ED1};
cus_mux41_buf inst_cus_mux41_buf_to_SD1 (
    .A0(to_SD1_input[0]),
    .A1(to_SD1_input[1]),
    .A2(to_SD1_input[2]),
    .A3(to_SD1_input[3]),
    .S0(ConfigBits[154+0]),
    .S0N(ConfigBits_N[154+0]),
    .S1(ConfigBits[154+1]),
    .S1N(ConfigBits_N[154+1]),
    .X(to_SD1)
);

 //switch matrix multiplexer to_SD2 MUX-4
assign to_SD2_input = {from_SD2,from_ND2,from_WD_1s0,from_ED2};
cus_mux41_buf inst_cus_mux41_buf_to_SD2 (
    .A0(to_SD2_input[0]),
    .A1(to_SD2_input[1]),
    .A2(to_SD2_input[2]),
    .A3(to_SD2_input[3]),
    .S0(ConfigBits[156+0]),
    .S0N(ConfigBits_N[156+0]),
    .S1(ConfigBits[156+1]),
    .S1N(ConfigBits_N[156+1]),
    .X(to_SD2)
);

 //switch matrix multiplexer to_SD3 MUX-4
assign to_SD3_input = {from_SD3,from_ND3,from_WD_1s1,from_ED3};
cus_mux41_buf inst_cus_mux41_buf_to_SD3 (
    .A0(to_SD3_input[0]),
    .A1(to_SD3_input[1]),
    .A2(to_SD3_input[2]),
    .A3(to_SD3_input[3]),
    .S0(ConfigBits[158+0]),
    .S0N(ConfigBits_N[158+0]),
    .S1(ConfigBits[158+1]),
    .S1N(ConfigBits_N[158+1]),
    .X(to_SD3)
);

 //switch matrix multiplexer to_SF0 MUX-4
assign to_SF0_input = {GND0,from_SF0,from_NF0,from_EF0};
cus_mux41_buf inst_cus_mux41_buf_to_SF0 (
    .A0(to_SF0_input[0]),
    .A1(to_SF0_input[1]),
    .A2(to_SF0_input[2]),
    .A3(to_SF0_input[3]),
    .S0(ConfigBits[160+0]),
    .S0N(ConfigBits_N[160+0]),
    .S1(ConfigBits[160+1]),
    .S1N(ConfigBits_N[160+1]),
    .X(to_SF0)
);

 //switch matrix multiplexer to_SF1 MUX-4
assign to_SF1_input = {VCC0,from_SF1,from_NF1,from_EF1};
cus_mux41_buf inst_cus_mux41_buf_to_SF1 (
    .A0(to_SF1_input[0]),
    .A1(to_SF1_input[1]),
    .A2(to_SF1_input[2]),
    .A3(to_SF1_input[3]),
    .S0(ConfigBits[162+0]),
    .S0N(ConfigBits_N[162+0]),
    .S1(ConfigBits[162+1]),
    .S1N(ConfigBits_N[162+1]),
    .X(to_SF1)
);

 //switch matrix multiplexer to_SF2 MUX-4
assign to_SF2_input = {from_SF2,from_NF2,from_WF_1s0,from_EF2};
cus_mux41_buf inst_cus_mux41_buf_to_SF2 (
    .A0(to_SF2_input[0]),
    .A1(to_SF2_input[1]),
    .A2(to_SF2_input[2]),
    .A3(to_SF2_input[3]),
    .S0(ConfigBits[164+0]),
    .S0N(ConfigBits_N[164+0]),
    .S1(ConfigBits[164+1]),
    .S1N(ConfigBits_N[164+1]),
    .X(to_SF2)
);

 //switch matrix multiplexer to_SF3 MUX-4
assign to_SF3_input = {from_SF3,from_NF3,from_WF_1s1,from_EF3};
cus_mux41_buf inst_cus_mux41_buf_to_SF3 (
    .A0(to_SF3_input[0]),
    .A1(to_SF3_input[1]),
    .A2(to_SF3_input[2]),
    .A3(to_SF3_input[3]),
    .S0(ConfigBits[166+0]),
    .S0N(ConfigBits_N[166+0]),
    .S1(ConfigBits[166+1]),
    .S1N(ConfigBits_N[166+1]),
    .X(to_SF3)
);

 //switch matrix multiplexer to_SG0 MUX-4
assign to_SG0_input = {GND0,from_SG0,from_NG0,from_EG0};
cus_mux41_buf inst_cus_mux41_buf_to_SG0 (
    .A0(to_SG0_input[0]),
    .A1(to_SG0_input[1]),
    .A2(to_SG0_input[2]),
    .A3(to_SG0_input[3]),
    .S0(ConfigBits[168+0]),
    .S0N(ConfigBits_N[168+0]),
    .S1(ConfigBits[168+1]),
    .S1N(ConfigBits_N[168+1]),
    .X(to_SG0)
);

 //switch matrix multiplexer to_SG1 MUX-4
assign to_SG1_input = {VCC0,from_SG1,from_NG1,from_EG1};
cus_mux41_buf inst_cus_mux41_buf_to_SG1 (
    .A0(to_SG1_input[0]),
    .A1(to_SG1_input[1]),
    .A2(to_SG1_input[2]),
    .A3(to_SG1_input[3]),
    .S0(ConfigBits[170+0]),
    .S0N(ConfigBits_N[170+0]),
    .S1(ConfigBits[170+1]),
    .S1N(ConfigBits_N[170+1]),
    .X(to_SG1)
);

 //switch matrix multiplexer to_SG2 MUX-4
assign to_SG2_input = {from_SG2,from_NG2,from_WG_1s0,from_EG2};
cus_mux41_buf inst_cus_mux41_buf_to_SG2 (
    .A0(to_SG2_input[0]),
    .A1(to_SG2_input[1]),
    .A2(to_SG2_input[2]),
    .A3(to_SG2_input[3]),
    .S0(ConfigBits[172+0]),
    .S0N(ConfigBits_N[172+0]),
    .S1(ConfigBits[172+1]),
    .S1N(ConfigBits_N[172+1]),
    .X(to_SG2)
);

 //switch matrix multiplexer to_SG3 MUX-4
assign to_SG3_input = {from_SG3,from_NG3,from_WG_1s1,from_EG3};
cus_mux41_buf inst_cus_mux41_buf_to_SG3 (
    .A0(to_SG3_input[0]),
    .A1(to_SG3_input[1]),
    .A2(to_SG3_input[2]),
    .A3(to_SG3_input[3]),
    .S0(ConfigBits[174+0]),
    .S0N(ConfigBits_N[174+0]),
    .S1(ConfigBits[174+1]),
    .S1N(ConfigBits_N[174+1]),
    .X(to_SG3)
);

 //switch matrix multiplexer to_SH0 MUX-4
assign to_SH0_input = {GND0,from_SH0,from_NH0,from_EH0};
cus_mux41_buf inst_cus_mux41_buf_to_SH0 (
    .A0(to_SH0_input[0]),
    .A1(to_SH0_input[1]),
    .A2(to_SH0_input[2]),
    .A3(to_SH0_input[3]),
    .S0(ConfigBits[176+0]),
    .S0N(ConfigBits_N[176+0]),
    .S1(ConfigBits[176+1]),
    .S1N(ConfigBits_N[176+1]),
    .X(to_SH0)
);

 //switch matrix multiplexer to_SH1 MUX-4
assign to_SH1_input = {VCC0,from_SH1,from_NH1,from_EH1};
cus_mux41_buf inst_cus_mux41_buf_to_SH1 (
    .A0(to_SH1_input[0]),
    .A1(to_SH1_input[1]),
    .A2(to_SH1_input[2]),
    .A3(to_SH1_input[3]),
    .S0(ConfigBits[178+0]),
    .S0N(ConfigBits_N[178+0]),
    .S1(ConfigBits[178+1]),
    .S1N(ConfigBits_N[178+1]),
    .X(to_SH1)
);

 //switch matrix multiplexer to_SH2 MUX-4
assign to_SH2_input = {from_SH2,from_NH2,from_WH_1s0,from_EH2};
cus_mux41_buf inst_cus_mux41_buf_to_SH2 (
    .A0(to_SH2_input[0]),
    .A1(to_SH2_input[1]),
    .A2(to_SH2_input[2]),
    .A3(to_SH2_input[3]),
    .S0(ConfigBits[180+0]),
    .S0N(ConfigBits_N[180+0]),
    .S1(ConfigBits[180+1]),
    .S1N(ConfigBits_N[180+1]),
    .X(to_SH2)
);

 //switch matrix multiplexer to_SH3 MUX-4
assign to_SH3_input = {from_SH3,from_NH3,from_WH_1s1,from_EH3};
cus_mux41_buf inst_cus_mux41_buf_to_SH3 (
    .A0(to_SH3_input[0]),
    .A1(to_SH3_input[1]),
    .A2(to_SH3_input[2]),
    .A3(to_SH3_input[3]),
    .S0(ConfigBits[182+0]),
    .S0N(ConfigBits_N[182+0]),
    .S1(ConfigBits[182+1]),
    .S1N(ConfigBits_N[182+1]),
    .X(to_SH3)
);

 //switch matrix multiplexer to_SI0 MUX-4
assign to_SI0_input = {GND0,from_SI0,from_NI0,from_EI0};
cus_mux41_buf inst_cus_mux41_buf_to_SI0 (
    .A0(to_SI0_input[0]),
    .A1(to_SI0_input[1]),
    .A2(to_SI0_input[2]),
    .A3(to_SI0_input[3]),
    .S0(ConfigBits[184+0]),
    .S0N(ConfigBits_N[184+0]),
    .S1(ConfigBits[184+1]),
    .S1N(ConfigBits_N[184+1]),
    .X(to_SI0)
);

 //switch matrix multiplexer to_SI1 MUX-4
assign to_SI1_input = {VCC0,from_SI1,from_NI1,from_EI1};
cus_mux41_buf inst_cus_mux41_buf_to_SI1 (
    .A0(to_SI1_input[0]),
    .A1(to_SI1_input[1]),
    .A2(to_SI1_input[2]),
    .A3(to_SI1_input[3]),
    .S0(ConfigBits[186+0]),
    .S0N(ConfigBits_N[186+0]),
    .S1(ConfigBits[186+1]),
    .S1N(ConfigBits_N[186+1]),
    .X(to_SI1)
);

 //switch matrix multiplexer to_SI2 MUX-4
assign to_SI2_input = {from_SI2,from_NI2,from_WI_1s0,from_EI2};
cus_mux41_buf inst_cus_mux41_buf_to_SI2 (
    .A0(to_SI2_input[0]),
    .A1(to_SI2_input[1]),
    .A2(to_SI2_input[2]),
    .A3(to_SI2_input[3]),
    .S0(ConfigBits[188+0]),
    .S0N(ConfigBits_N[188+0]),
    .S1(ConfigBits[188+1]),
    .S1N(ConfigBits_N[188+1]),
    .X(to_SI2)
);

 //switch matrix multiplexer to_SI3 MUX-4
assign to_SI3_input = {from_SI3,from_NI3,from_WI_1s1,from_EI3};
cus_mux41_buf inst_cus_mux41_buf_to_SI3 (
    .A0(to_SI3_input[0]),
    .A1(to_SI3_input[1]),
    .A2(to_SI3_input[2]),
    .A3(to_SI3_input[3]),
    .S0(ConfigBits[190+0]),
    .S0N(ConfigBits_N[190+0]),
    .S1(ConfigBits[190+1]),
    .S1N(ConfigBits_N[190+1]),
    .X(to_SI3)
);

endmodule