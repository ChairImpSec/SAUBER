module top_wrapper;
wire [59:0] io_in_0t, io_in_0f, io_in_1t, io_in_1f, io_out_0t, io_out_0f, io_out_1t, io_out_1f, io_oeb, ctrl_io_in_0t, ctrl_io_in_0f, ctrl_io_out_0t, ctrl_io_out_0f, ctrl_io_oeb;
 
// IO
 
(* keep, BEL="X0Y1.A" *) IO_1_bidirectional_frame_config_pass io0_i (.Q0_t(io_in_0t[0]), .Q0_f(io_in_0f[0]), .Q1_t(io_in_1t[0]), .Q1_f(io_in_1f[0]), .I0_t(io_out_0t[0]), .I0_f(io_out_0f[0]), .I1_t(io_out_1t[0]), .I1_f(io_out_1f[0]), .T(io_oeb[0]));
(* keep, BEL="X0Y2.A" *) IO_1_bidirectional_frame_config_pass io1_i (.Q0_t(io_in_0t[1]), .Q0_f(io_in_0f[1]), .Q1_t(io_in_1t[1]), .Q1_f(io_in_1f[1]), .I0_t(io_out_0t[1]), .I0_f(io_out_0f[1]), .I1_t(io_out_1t[1]), .I1_f(io_out_1f[1]), .T(io_oeb[1]));
(* keep, BEL="X0Y3.A" *) IO_1_bidirectional_frame_config_pass io2_i (.Q0_t(io_in_0t[2]), .Q0_f(io_in_0f[2]), .Q1_t(io_in_1t[2]), .Q1_f(io_in_1f[2]), .I0_t(io_out_0t[2]), .I0_f(io_out_0f[2]), .I1_t(io_out_1t[2]), .I1_f(io_out_1f[2]), .T(io_oeb[2]));
(* keep, BEL="X0Y4.A" *) IO_1_bidirectional_frame_config_pass io3_i (.Q0_t(io_in_0t[3]), .Q0_f(io_in_0f[3]), .Q1_t(io_in_1t[3]), .Q1_f(io_in_1f[3]), .I0_t(io_out_0t[3]), .I0_f(io_out_0f[3]), .I1_t(io_out_1t[3]), .I1_f(io_out_1f[3]), .T(io_oeb[3]));
(* keep, BEL="X0Y5.A" *) IO_1_bidirectional_frame_config_pass io4_i (.Q0_t(io_in_0t[4]), .Q0_f(io_in_0f[4]), .Q1_t(io_in_1t[4]), .Q1_f(io_in_1f[4]), .I0_t(io_out_0t[4]), .I0_f(io_out_0f[4]), .I1_t(io_out_1t[4]), .I1_f(io_out_1f[4]), .T(io_oeb[4]));
(* keep, BEL="X0Y6.A" *) IO_1_bidirectional_frame_config_pass io5_i (.Q0_t(io_in_0t[5]), .Q0_f(io_in_0f[5]), .Q1_t(io_in_1t[5]), .Q1_f(io_in_1f[5]), .I0_t(io_out_0t[5]), .I0_f(io_out_0f[5]), .I1_t(io_out_1t[5]), .I1_f(io_out_1f[5]), .T(io_oeb[5]));
(* keep, BEL="X0Y7.A" *) IO_1_bidirectional_frame_config_pass io6_i (.Q0_t(io_in_0t[6]), .Q0_f(io_in_0f[6]), .Q1_t(io_in_1t[6]), .Q1_f(io_in_1f[6]), .I0_t(io_out_0t[6]), .I0_f(io_out_0f[6]), .I1_t(io_out_1t[6]), .I1_f(io_out_1f[6]), .T(io_oeb[6]));
(* keep, BEL="X0Y8.A" *) IO_1_bidirectional_frame_config_pass io7_i (.Q0_t(io_in_0t[7]), .Q0_f(io_in_0f[7]), .Q1_t(io_in_1t[7]), .Q1_f(io_in_1f[7]), .I0_t(io_out_0t[7]), .I0_f(io_out_0f[7]), .I1_t(io_out_1t[7]), .I1_f(io_out_1f[7]), .T(io_oeb[7]));
(* keep, BEL="X0Y9.A" *) IO_1_bidirectional_frame_config_pass io8_i (.Q0_t(io_in_0t[8]), .Q0_f(io_in_0f[8]), .Q1_t(io_in_1t[8]), .Q1_f(io_in_1f[8]), .I0_t(io_out_0t[8]), .I0_f(io_out_0f[8]), .I1_t(io_out_1t[8]), .I1_f(io_out_1f[8]), .T(io_oeb[8]));
(* keep, BEL="X0Y10.A" *) IO_1_bidirectional_frame_config_pass io9_i (.Q0_t(io_in_0t[9]), .Q0_f(io_in_0f[9]), .Q1_t(io_in_1t[9]), .Q1_f(io_in_1f[9]), .I0_t(io_out_0t[9]), .I0_f(io_out_0f[9]), .I1_t(io_out_1t[9]), .I1_f(io_out_1f[9]), .T(io_oeb[9]));
(* keep, BEL="X0Y11.A" *) IO_1_bidirectional_frame_config_pass io10_i (.Q0_t(io_in_0t[10]), .Q0_f(io_in_0f[10]), .Q1_t(io_in_1t[10]), .Q1_f(io_in_1f[10]), .I0_t(io_out_0t[10]), .I0_f(io_out_0f[10]), .I1_t(io_out_1t[10]), .I1_f(io_out_1f[10]), .T(io_oeb[10]));
(* keep, BEL="X0Y12.A" *) IO_1_bidirectional_frame_config_pass io11_i (.Q0_t(io_in_0t[11]), .Q0_f(io_in_0f[11]), .Q1_t(io_in_1t[11]), .Q1_f(io_in_1f[11]), .I0_t(io_out_0t[11]), .I0_f(io_out_0f[11]), .I1_t(io_out_1t[11]), .I1_f(io_out_1f[11]), .T(io_oeb[11]));
(* keep, BEL="X0Y13.A" *) IO_1_bidirectional_frame_config_pass io12_i (.Q0_t(io_in_0t[12]), .Q0_f(io_in_0f[12]), .Q1_t(io_in_1t[12]), .Q1_f(io_in_1f[12]), .I0_t(io_out_0t[12]), .I0_f(io_out_0f[12]), .I1_t(io_out_1t[12]), .I1_f(io_out_1f[12]), .T(io_oeb[12]));
(* keep, BEL="X0Y14.A" *) IO_1_bidirectional_frame_config_pass io13_i (.Q0_t(io_in_0t[13]), .Q0_f(io_in_0f[13]), .Q1_t(io_in_1t[13]), .Q1_f(io_in_1f[13]), .I0_t(io_out_0t[13]), .I0_f(io_out_0f[13]), .I1_t(io_out_1t[13]), .I1_f(io_out_1f[13]), .T(io_oeb[13]));
(* keep, BEL="X0Y15.A" *) IO_1_bidirectional_frame_config_pass io14_i (.Q0_t(io_in_0t[14]), .Q0_f(io_in_0f[14]), .Q1_t(io_in_1t[14]), .Q1_f(io_in_1f[14]), .I0_t(io_out_0t[14]), .I0_f(io_out_0f[14]), .I1_t(io_out_1t[14]), .I1_f(io_out_1f[14]), .T(io_oeb[14]));
(* keep, BEL="X0Y16.A" *) IO_1_bidirectional_frame_config_pass io15_i (.Q0_t(io_in_0t[15]), .Q0_f(io_in_0f[15]), .Q1_t(io_in_1t[15]), .Q1_f(io_in_1f[15]), .I0_t(io_out_0t[15]), .I0_f(io_out_0f[15]), .I1_t(io_out_1t[15]), .I1_f(io_out_1f[15]), .T(io_oeb[15]));
(* keep, BEL="X0Y17.A" *) IO_1_bidirectional_frame_config_pass io16_i (.Q0_t(io_in_0t[16]), .Q0_f(io_in_0f[16]), .Q1_t(io_in_1t[16]), .Q1_f(io_in_1f[16]), .I0_t(io_out_0t[16]), .I0_f(io_out_0f[16]), .I1_t(io_out_1t[16]), .I1_f(io_out_1f[16]), .T(io_oeb[16]));
(* keep, BEL="X0Y18.A" *) IO_1_bidirectional_frame_config_pass io17_i (.Q0_t(io_in_0t[17]), .Q0_f(io_in_0f[17]), .Q1_t(io_in_1t[17]), .Q1_f(io_in_1f[17]), .I0_t(io_out_0t[17]), .I0_f(io_out_0f[17]), .I1_t(io_out_1t[17]), .I1_f(io_out_1f[17]), .T(io_oeb[17]));
(* keep, BEL="X0Y19.A" *) IO_1_bidirectional_frame_config_pass io18_i (.Q0_t(io_in_0t[18]), .Q0_f(io_in_0f[18]), .Q1_t(io_in_1t[18]), .Q1_f(io_in_1f[18]), .I0_t(io_out_0t[18]), .I0_f(io_out_0f[18]), .I1_t(io_out_1t[18]), .I1_f(io_out_1f[18]), .T(io_oeb[18]));
(* keep, BEL="X0Y20.A" *) IO_1_bidirectional_frame_config_pass io19_i (.Q0_t(io_in_0t[19]), .Q0_f(io_in_0f[19]), .Q1_t(io_in_1t[19]), .Q1_f(io_in_1f[19]), .I0_t(io_out_0t[19]), .I0_f(io_out_0f[19]), .I1_t(io_out_1t[19]), .I1_f(io_out_1f[19]), .T(io_oeb[19]));
(* keep, BEL="X0Y21.A" *) IO_1_bidirectional_frame_config_pass io20_i (.Q0_t(io_in_0t[20]), .Q0_f(io_in_0f[20]), .Q1_t(io_in_1t[20]), .Q1_f(io_in_1f[20]), .I0_t(io_out_0t[20]), .I0_f(io_out_0f[20]), .I1_t(io_out_1t[20]), .I1_f(io_out_1f[20]), .T(io_oeb[20]));
(* keep, BEL="X0Y22.A" *) IO_1_bidirectional_frame_config_pass io21_i (.Q0_t(io_in_0t[21]), .Q0_f(io_in_0f[21]), .Q1_t(io_in_1t[21]), .Q1_f(io_in_1f[21]), .I0_t(io_out_0t[21]), .I0_f(io_out_0f[21]), .I1_t(io_out_1t[21]), .I1_f(io_out_1f[21]), .T(io_oeb[21]));
(* keep, BEL="X0Y23.A" *) IO_1_bidirectional_frame_config_pass io22_i (.Q0_t(io_in_0t[22]), .Q0_f(io_in_0f[22]), .Q1_t(io_in_1t[22]), .Q1_f(io_in_1f[22]), .I0_t(io_out_0t[22]), .I0_f(io_out_0f[22]), .I1_t(io_out_1t[22]), .I1_f(io_out_1f[22]), .T(io_oeb[22]));
(* keep, BEL="X0Y24.A" *) IO_1_bidirectional_frame_config_pass io23_i (.Q0_t(io_in_0t[23]), .Q0_f(io_in_0f[23]), .Q1_t(io_in_1t[23]), .Q1_f(io_in_1f[23]), .I0_t(io_out_0t[23]), .I0_f(io_out_0f[23]), .I1_t(io_out_1t[23]), .I1_f(io_out_1f[23]), .T(io_oeb[23]));
(* keep, BEL="X0Y25.A" *) IO_1_bidirectional_frame_config_pass io24_i (.Q0_t(io_in_0t[24]), .Q0_f(io_in_0f[24]), .Q1_t(io_in_1t[24]), .Q1_f(io_in_1f[24]), .I0_t(io_out_0t[24]), .I0_f(io_out_0f[24]), .I1_t(io_out_1t[24]), .I1_f(io_out_1f[24]), .T(io_oeb[24]));
(* keep, BEL="X0Y26.A" *) IO_1_bidirectional_frame_config_pass io25_i (.Q0_t(io_in_0t[25]), .Q0_f(io_in_0f[25]), .Q1_t(io_in_1t[25]), .Q1_f(io_in_1f[25]), .I0_t(io_out_0t[25]), .I0_f(io_out_0f[25]), .I1_t(io_out_1t[25]), .I1_f(io_out_1f[25]), .T(io_oeb[25]));
(* keep, BEL="X0Y27.A" *) IO_1_bidirectional_frame_config_pass io26_i (.Q0_t(io_in_0t[26]), .Q0_f(io_in_0f[26]), .Q1_t(io_in_1t[26]), .Q1_f(io_in_1f[26]), .I0_t(io_out_0t[26]), .I0_f(io_out_0f[26]), .I1_t(io_out_1t[26]), .I1_f(io_out_1f[26]), .T(io_oeb[26]));
(* keep, BEL="X0Y28.A" *) IO_1_bidirectional_frame_config_pass io27_i (.Q0_t(io_in_0t[27]), .Q0_f(io_in_0f[27]), .Q1_t(io_in_1t[27]), .Q1_f(io_in_1f[27]), .I0_t(io_out_0t[27]), .I0_f(io_out_0f[27]), .I1_t(io_out_1t[27]), .I1_f(io_out_1f[27]), .T(io_oeb[27]));
(* keep, BEL="X0Y29.A" *) IO_1_bidirectional_frame_config_pass io28_i (.Q0_t(io_in_0t[28]), .Q0_f(io_in_0f[28]), .Q1_t(io_in_1t[28]), .Q1_f(io_in_1f[28]), .I0_t(io_out_0t[28]), .I0_f(io_out_0f[28]), .I1_t(io_out_1t[28]), .I1_f(io_out_1f[28]), .T(io_oeb[28]));
(* keep, BEL="X0Y30.A" *) IO_1_bidirectional_frame_config_pass io29_i (.Q0_t(io_in_0t[29]), .Q0_f(io_in_0f[29]), .Q1_t(io_in_1t[29]), .Q1_f(io_in_1f[29]), .I0_t(io_out_0t[29]), .I0_f(io_out_0f[29]), .I1_t(io_out_1t[29]), .I1_f(io_out_1f[29]), .T(io_oeb[29]));
(* keep, BEL="X0Y31.A" *) IO_1_bidirectional_frame_config_pass io30_i (.Q0_t(io_in_0t[30]), .Q0_f(io_in_0f[30]), .Q1_t(io_in_1t[30]), .Q1_f(io_in_1f[30]), .I0_t(io_out_0t[30]), .I0_f(io_out_0f[30]), .I1_t(io_out_1t[30]), .I1_f(io_out_1f[30]), .T(io_oeb[30]));
(* keep, BEL="X0Y32.A" *) IO_1_bidirectional_frame_config_pass io31_i (.Q0_t(io_in_0t[31]), .Q0_f(io_in_0f[31]), .Q1_t(io_in_1t[31]), .Q1_f(io_in_1f[31]), .I0_t(io_out_0t[31]), .I0_f(io_out_0f[31]), .I1_t(io_out_1t[31]), .I1_f(io_out_1f[31]), .T(io_oeb[31]));
(* keep, BEL="X0Y33.A" *) IO_1_bidirectional_frame_config_pass io32_i (.Q0_t(io_in_0t[32]), .Q0_f(io_in_0f[32]), .Q1_t(io_in_1t[32]), .Q1_f(io_in_1f[32]), .I0_t(io_out_0t[32]), .I0_f(io_out_0f[32]), .I1_t(io_out_1t[32]), .I1_f(io_out_1f[32]), .T(io_oeb[32]));
(* keep, BEL="X0Y34.A" *) IO_1_bidirectional_frame_config_pass io33_i (.Q0_t(io_in_0t[33]), .Q0_f(io_in_0f[33]), .Q1_t(io_in_1t[33]), .Q1_f(io_in_1f[33]), .I0_t(io_out_0t[33]), .I0_f(io_out_0f[33]), .I1_t(io_out_1t[33]), .I1_f(io_out_1f[33]), .T(io_oeb[33]));
(* keep, BEL="X0Y35.A" *) IO_1_bidirectional_frame_config_pass io34_i (.Q0_t(io_in_0t[34]), .Q0_f(io_in_0f[34]), .Q1_t(io_in_1t[34]), .Q1_f(io_in_1f[34]), .I0_t(io_out_0t[34]), .I0_f(io_out_0f[34]), .I1_t(io_out_1t[34]), .I1_f(io_out_1f[34]), .T(io_oeb[34]));
(* keep, BEL="X0Y36.A" *) IO_1_bidirectional_frame_config_pass io35_i (.Q0_t(io_in_0t[35]), .Q0_f(io_in_0f[35]), .Q1_t(io_in_1t[35]), .Q1_f(io_in_1f[35]), .I0_t(io_out_0t[35]), .I0_f(io_out_0f[35]), .I1_t(io_out_1t[35]), .I1_f(io_out_1f[35]), .T(io_oeb[35]));
(* keep, BEL="X0Y37.A" *) IO_1_bidirectional_frame_config_pass io36_i (.Q0_t(io_in_0t[36]), .Q0_f(io_in_0f[36]), .Q1_t(io_in_1t[36]), .Q1_f(io_in_1f[36]), .I0_t(io_out_0t[36]), .I0_f(io_out_0f[36]), .I1_t(io_out_1t[36]), .I1_f(io_out_1f[36]), .T(io_oeb[36]));
(* keep, BEL="X0Y38.A" *) IO_1_bidirectional_frame_config_pass io37_i (.Q0_t(io_in_0t[37]), .Q0_f(io_in_0f[37]), .Q1_t(io_in_1t[37]), .Q1_f(io_in_1f[37]), .I0_t(io_out_0t[37]), .I0_f(io_out_0f[37]), .I1_t(io_out_1t[37]), .I1_f(io_out_1f[37]), .T(io_oeb[37]));
(* keep, BEL="X0Y39.A" *) IO_1_bidirectional_frame_config_pass io38_i (.Q0_t(io_in_0t[38]), .Q0_f(io_in_0f[38]), .Q1_t(io_in_1t[38]), .Q1_f(io_in_1f[38]), .I0_t(io_out_0t[38]), .I0_f(io_out_0f[38]), .I1_t(io_out_1t[38]), .I1_f(io_out_1f[38]), .T(io_oeb[38]));
(* keep, BEL="X0Y40.A" *) IO_1_bidirectional_frame_config_pass io39_i (.Q0_t(io_in_0t[39]), .Q0_f(io_in_0f[39]), .Q1_t(io_in_1t[39]), .Q1_f(io_in_1f[39]), .I0_t(io_out_0t[39]), .I0_f(io_out_0f[39]), .I1_t(io_out_1t[39]), .I1_f(io_out_1f[39]), .T(io_oeb[39]));
(* keep, BEL="X0Y41.A" *) IO_1_bidirectional_frame_config_pass io40_i (.Q0_t(io_in_0t[40]), .Q0_f(io_in_0f[40]), .Q1_t(io_in_1t[40]), .Q1_f(io_in_1f[40]), .I0_t(io_out_0t[40]), .I0_f(io_out_0f[40]), .I1_t(io_out_1t[40]), .I1_f(io_out_1f[40]), .T(io_oeb[40]));
(* keep, BEL="X0Y42.A" *) IO_1_bidirectional_frame_config_pass io41_i (.Q0_t(io_in_0t[41]), .Q0_f(io_in_0f[41]), .Q1_t(io_in_1t[41]), .Q1_f(io_in_1f[41]), .I0_t(io_out_0t[41]), .I0_f(io_out_0f[41]), .I1_t(io_out_1t[41]), .I1_f(io_out_1f[41]), .T(io_oeb[41]));
(* keep, BEL="X0Y43.A" *) IO_1_bidirectional_frame_config_pass io42_i (.Q0_t(io_in_0t[42]), .Q0_f(io_in_0f[42]), .Q1_t(io_in_1t[42]), .Q1_f(io_in_1f[42]), .I0_t(io_out_0t[42]), .I0_f(io_out_0f[42]), .I1_t(io_out_1t[42]), .I1_f(io_out_1f[42]), .T(io_oeb[42]));
(* keep, BEL="X0Y44.A" *) IO_1_bidirectional_frame_config_pass io43_i (.Q0_t(io_in_0t[43]), .Q0_f(io_in_0f[43]), .Q1_t(io_in_1t[43]), .Q1_f(io_in_1f[43]), .I0_t(io_out_0t[43]), .I0_f(io_out_0f[43]), .I1_t(io_out_1t[43]), .I1_f(io_out_1f[43]), .T(io_oeb[43]));
(* keep, BEL="X0Y45.A" *) IO_1_bidirectional_frame_config_pass io44_i (.Q0_t(io_in_0t[44]), .Q0_f(io_in_0f[44]), .Q1_t(io_in_1t[44]), .Q1_f(io_in_1f[44]), .I0_t(io_out_0t[44]), .I0_f(io_out_0f[44]), .I1_t(io_out_1t[44]), .I1_f(io_out_1f[44]), .T(io_oeb[44]));
(* keep, BEL="X0Y46.A" *) IO_1_bidirectional_frame_config_pass io45_i (.Q0_t(io_in_0t[45]), .Q0_f(io_in_0f[45]), .Q1_t(io_in_1t[45]), .Q1_f(io_in_1f[45]), .I0_t(io_out_0t[45]), .I0_f(io_out_0f[45]), .I1_t(io_out_1t[45]), .I1_f(io_out_1f[45]), .T(io_oeb[45]));
(* keep, BEL="X0Y47.A" *) IO_1_bidirectional_frame_config_pass io46_i (.Q0_t(io_in_0t[46]), .Q0_f(io_in_0f[46]), .Q1_t(io_in_1t[46]), .Q1_f(io_in_1f[46]), .I0_t(io_out_0t[46]), .I0_f(io_out_0f[46]), .I1_t(io_out_1t[46]), .I1_f(io_out_1f[46]), .T(io_oeb[46]));
(* keep, BEL="X0Y48.A" *) IO_1_bidirectional_frame_config_pass io47_i (.Q0_t(io_in_0t[47]), .Q0_f(io_in_0f[47]), .Q1_t(io_in_1t[47]), .Q1_f(io_in_1f[47]), .I0_t(io_out_0t[47]), .I0_f(io_out_0f[47]), .I1_t(io_out_1t[47]), .I1_f(io_out_1f[47]), .T(io_oeb[47]));
(* keep, BEL="X0Y49.A" *) IO_1_bidirectional_frame_config_pass io48_i (.Q0_t(io_in_0t[48]), .Q0_f(io_in_0f[48]), .Q1_t(io_in_1t[48]), .Q1_f(io_in_1f[48]), .I0_t(io_out_0t[48]), .I0_f(io_out_0f[48]), .I1_t(io_out_1t[48]), .I1_f(io_out_1f[48]), .T(io_oeb[48]));
(* keep, BEL="X0Y50.A" *) IO_1_bidirectional_frame_config_pass io49_i (.Q0_t(io_in_0t[49]), .Q0_f(io_in_0f[49]), .Q1_t(io_in_1t[49]), .Q1_f(io_in_1f[49]), .I0_t(io_out_0t[49]), .I0_f(io_out_0f[49]), .I1_t(io_out_1t[49]), .I1_f(io_out_1f[49]), .T(io_oeb[49]));
(* keep, BEL="X0Y51.A" *) IO_1_bidirectional_frame_config_pass io50_i (.Q0_t(io_in_0t[50]), .Q0_f(io_in_0f[50]), .Q1_t(io_in_1t[50]), .Q1_f(io_in_1f[50]), .I0_t(io_out_0t[50]), .I0_f(io_out_0f[50]), .I1_t(io_out_1t[50]), .I1_f(io_out_1f[50]), .T(io_oeb[50]));
(* keep, BEL="X0Y52.A" *) IO_1_bidirectional_frame_config_pass io51_i (.Q0_t(io_in_0t[51]), .Q0_f(io_in_0f[51]), .Q1_t(io_in_1t[51]), .Q1_f(io_in_1f[51]), .I0_t(io_out_0t[51]), .I0_f(io_out_0f[51]), .I1_t(io_out_1t[51]), .I1_f(io_out_1f[51]), .T(io_oeb[51]));
(* keep, BEL="X0Y53.A" *) IO_1_bidirectional_frame_config_pass io52_i (.Q0_t(io_in_0t[52]), .Q0_f(io_in_0f[52]), .Q1_t(io_in_1t[52]), .Q1_f(io_in_1f[52]), .I0_t(io_out_0t[52]), .I0_f(io_out_0f[52]), .I1_t(io_out_1t[52]), .I1_f(io_out_1f[52]), .T(io_oeb[52]));
(* keep, BEL="X0Y54.A" *) IO_1_bidirectional_frame_config_pass io53_i (.Q0_t(io_in_0t[53]), .Q0_f(io_in_0f[53]), .Q1_t(io_in_1t[53]), .Q1_f(io_in_1f[53]), .I0_t(io_out_0t[53]), .I0_f(io_out_0f[53]), .I1_t(io_out_1t[53]), .I1_f(io_out_1f[53]), .T(io_oeb[53]));
(* keep, BEL="X0Y55.A" *) IO_1_bidirectional_frame_config_pass io54_i (.Q0_t(io_in_0t[54]), .Q0_f(io_in_0f[54]), .Q1_t(io_in_1t[54]), .Q1_f(io_in_1f[54]), .I0_t(io_out_0t[54]), .I0_f(io_out_0f[54]), .I1_t(io_out_1t[54]), .I1_f(io_out_1f[54]), .T(io_oeb[54]));
(* keep, BEL="X0Y56.A" *) IO_1_bidirectional_frame_config_pass io55_i (.Q0_t(io_in_0t[55]), .Q0_f(io_in_0f[55]), .Q1_t(io_in_1t[55]), .Q1_f(io_in_1f[55]), .I0_t(io_out_0t[55]), .I0_f(io_out_0f[55]), .I1_t(io_out_1t[55]), .I1_f(io_out_1f[55]), .T(io_oeb[55]));
(* keep, BEL="X0Y57.A" *) IO_1_bidirectional_frame_config_pass io56_i (.Q0_t(io_in_0t[56]), .Q0_f(io_in_0f[56]), .Q1_t(io_in_1t[56]), .Q1_f(io_in_1f[56]), .I0_t(io_out_0t[56]), .I0_f(io_out_0f[56]), .I1_t(io_out_1t[56]), .I1_f(io_out_1f[56]), .T(io_oeb[56]));
(* keep, BEL="X0Y58.A" *) IO_1_bidirectional_frame_config_pass io57_i (.Q0_t(io_in_0t[57]), .Q0_f(io_in_0f[57]), .Q1_t(io_in_1t[57]), .Q1_f(io_in_1f[57]), .I0_t(io_out_0t[57]), .I0_f(io_out_0f[57]), .I1_t(io_out_1t[57]), .I1_f(io_out_1f[57]), .T(io_oeb[57]));
(* keep, BEL="X0Y59.A" *) IO_1_bidirectional_frame_config_pass io58_i (.Q0_t(io_in_0t[58]), .Q0_f(io_in_0f[58]), .Q1_t(io_in_1t[58]), .Q1_f(io_in_1f[58]), .I0_t(io_out_0t[58]), .I0_f(io_out_0f[58]), .I1_t(io_out_1t[58]), .I1_f(io_out_1f[58]), .T(io_oeb[58]));
(* keep, BEL="X0Y60.A" *) IO_1_bidirectional_frame_config_pass io59_i (.Q0_t(io_in_0t[59]), .Q0_f(io_in_0f[59]), .Q1_t(io_in_1t[59]), .Q1_f(io_in_1f[59]), .I0_t(io_out_0t[59]), .I0_f(io_out_0f[59]), .I1_t(io_out_1t[59]), .I1_f(io_out_1f[59]), .T(io_oeb[59]));
 
// ctrl IO
 
(* keep, BEL="X38Y1.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io0_i (.Q0_t(ctrl_io_in_0t[0]), .Q0_f(ctrl_io_in_0f[0]), .I0_t(ctrl_io_out_0t[0]), .I0_f(ctrl_io_out_0f[0]), .T(ctrl_io_oeb[0]));
(* keep, BEL="X38Y2.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io1_i (.Q0_t(ctrl_io_in_0t[1]), .Q0_f(ctrl_io_in_0f[1]), .I0_t(ctrl_io_out_0t[1]), .I0_f(ctrl_io_out_0f[1]), .T(ctrl_io_oeb[1]));
(* keep, BEL="X38Y3.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io2_i (.Q0_t(ctrl_io_in_0t[2]), .Q0_f(ctrl_io_in_0f[2]), .I0_t(ctrl_io_out_0t[2]), .I0_f(ctrl_io_out_0f[2]), .T(ctrl_io_oeb[2]));
(* keep, BEL="X38Y4.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io3_i (.Q0_t(ctrl_io_in_0t[3]), .Q0_f(ctrl_io_in_0f[3]), .I0_t(ctrl_io_out_0t[3]), .I0_f(ctrl_io_out_0f[3]), .T(ctrl_io_oeb[3]));
(* keep, BEL="X38Y5.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io4_i (.Q0_t(ctrl_io_in_0t[4]), .Q0_f(ctrl_io_in_0f[4]), .I0_t(ctrl_io_out_0t[4]), .I0_f(ctrl_io_out_0f[4]), .T(ctrl_io_oeb[4]));
(* keep, BEL="X38Y6.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io5_i (.Q0_t(ctrl_io_in_0t[5]), .Q0_f(ctrl_io_in_0f[5]), .I0_t(ctrl_io_out_0t[5]), .I0_f(ctrl_io_out_0f[5]), .T(ctrl_io_oeb[5]));
(* keep, BEL="X38Y7.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io6_i (.Q0_t(ctrl_io_in_0t[6]), .Q0_f(ctrl_io_in_0f[6]), .I0_t(ctrl_io_out_0t[6]), .I0_f(ctrl_io_out_0f[6]), .T(ctrl_io_oeb[6]));
(* keep, BEL="X38Y8.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io7_i (.Q0_t(ctrl_io_in_0t[7]), .Q0_f(ctrl_io_in_0f[7]), .I0_t(ctrl_io_out_0t[7]), .I0_f(ctrl_io_out_0f[7]), .T(ctrl_io_oeb[7]));
(* keep, BEL="X38Y9.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io8_i (.Q0_t(ctrl_io_in_0t[8]), .Q0_f(ctrl_io_in_0f[8]), .I0_t(ctrl_io_out_0t[8]), .I0_f(ctrl_io_out_0f[8]), .T(ctrl_io_oeb[8]));
(* keep, BEL="X38Y10.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io9_i (.Q0_t(ctrl_io_in_0t[9]), .Q0_f(ctrl_io_in_0f[9]), .I0_t(ctrl_io_out_0t[9]), .I0_f(ctrl_io_out_0f[9]), .T(ctrl_io_oeb[9]));
(* keep, BEL="X38Y11.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io10_i (.Q0_t(ctrl_io_in_0t[10]), .Q0_f(ctrl_io_in_0f[10]), .I0_t(ctrl_io_out_0t[10]), .I0_f(ctrl_io_out_0f[10]), .T(ctrl_io_oeb[10]));
(* keep, BEL="X38Y12.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io11_i (.Q0_t(ctrl_io_in_0t[11]), .Q0_f(ctrl_io_in_0f[11]), .I0_t(ctrl_io_out_0t[11]), .I0_f(ctrl_io_out_0f[11]), .T(ctrl_io_oeb[11]));
(* keep, BEL="X38Y13.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io12_i (.Q0_t(ctrl_io_in_0t[12]), .Q0_f(ctrl_io_in_0f[12]), .I0_t(ctrl_io_out_0t[12]), .I0_f(ctrl_io_out_0f[12]), .T(ctrl_io_oeb[12]));
(* keep, BEL="X38Y14.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io13_i (.Q0_t(ctrl_io_in_0t[13]), .Q0_f(ctrl_io_in_0f[13]), .I0_t(ctrl_io_out_0t[13]), .I0_f(ctrl_io_out_0f[13]), .T(ctrl_io_oeb[13]));
(* keep, BEL="X38Y15.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io14_i (.Q0_t(ctrl_io_in_0t[14]), .Q0_f(ctrl_io_in_0f[14]), .I0_t(ctrl_io_out_0t[14]), .I0_f(ctrl_io_out_0f[14]), .T(ctrl_io_oeb[14]));
(* keep, BEL="X38Y16.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io15_i (.Q0_t(ctrl_io_in_0t[15]), .Q0_f(ctrl_io_in_0f[15]), .I0_t(ctrl_io_out_0t[15]), .I0_f(ctrl_io_out_0f[15]), .T(ctrl_io_oeb[15]));
(* keep, BEL="X38Y17.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io16_i (.Q0_t(ctrl_io_in_0t[16]), .Q0_f(ctrl_io_in_0f[16]), .I0_t(ctrl_io_out_0t[16]), .I0_f(ctrl_io_out_0f[16]), .T(ctrl_io_oeb[16]));
(* keep, BEL="X38Y18.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io17_i (.Q0_t(ctrl_io_in_0t[17]), .Q0_f(ctrl_io_in_0f[17]), .I0_t(ctrl_io_out_0t[17]), .I0_f(ctrl_io_out_0f[17]), .T(ctrl_io_oeb[17]));
(* keep, BEL="X38Y19.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io18_i (.Q0_t(ctrl_io_in_0t[18]), .Q0_f(ctrl_io_in_0f[18]), .I0_t(ctrl_io_out_0t[18]), .I0_f(ctrl_io_out_0f[18]), .T(ctrl_io_oeb[18]));
(* keep, BEL="X38Y20.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io19_i (.Q0_t(ctrl_io_in_0t[19]), .Q0_f(ctrl_io_in_0f[19]), .I0_t(ctrl_io_out_0t[19]), .I0_f(ctrl_io_out_0f[19]), .T(ctrl_io_oeb[19]));
(* keep, BEL="X38Y21.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io20_i (.Q0_t(ctrl_io_in_0t[20]), .Q0_f(ctrl_io_in_0f[20]), .I0_t(ctrl_io_out_0t[20]), .I0_f(ctrl_io_out_0f[20]), .T(ctrl_io_oeb[20]));
(* keep, BEL="X38Y22.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io21_i (.Q0_t(ctrl_io_in_0t[21]), .Q0_f(ctrl_io_in_0f[21]), .I0_t(ctrl_io_out_0t[21]), .I0_f(ctrl_io_out_0f[21]), .T(ctrl_io_oeb[21]));
(* keep, BEL="X38Y23.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io22_i (.Q0_t(ctrl_io_in_0t[22]), .Q0_f(ctrl_io_in_0f[22]), .I0_t(ctrl_io_out_0t[22]), .I0_f(ctrl_io_out_0f[22]), .T(ctrl_io_oeb[22]));
(* keep, BEL="X38Y24.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io23_i (.Q0_t(ctrl_io_in_0t[23]), .Q0_f(ctrl_io_in_0f[23]), .I0_t(ctrl_io_out_0t[23]), .I0_f(ctrl_io_out_0f[23]), .T(ctrl_io_oeb[23]));
(* keep, BEL="X38Y25.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io24_i (.Q0_t(ctrl_io_in_0t[24]), .Q0_f(ctrl_io_in_0f[24]), .I0_t(ctrl_io_out_0t[24]), .I0_f(ctrl_io_out_0f[24]), .T(ctrl_io_oeb[24]));
(* keep, BEL="X38Y26.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io25_i (.Q0_t(ctrl_io_in_0t[25]), .Q0_f(ctrl_io_in_0f[25]), .I0_t(ctrl_io_out_0t[25]), .I0_f(ctrl_io_out_0f[25]), .T(ctrl_io_oeb[25]));
(* keep, BEL="X38Y27.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io26_i (.Q0_t(ctrl_io_in_0t[26]), .Q0_f(ctrl_io_in_0f[26]), .I0_t(ctrl_io_out_0t[26]), .I0_f(ctrl_io_out_0f[26]), .T(ctrl_io_oeb[26]));
(* keep, BEL="X38Y28.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io27_i (.Q0_t(ctrl_io_in_0t[27]), .Q0_f(ctrl_io_in_0f[27]), .I0_t(ctrl_io_out_0t[27]), .I0_f(ctrl_io_out_0f[27]), .T(ctrl_io_oeb[27]));
(* keep, BEL="X38Y29.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io28_i (.Q0_t(ctrl_io_in_0t[28]), .Q0_f(ctrl_io_in_0f[28]), .I0_t(ctrl_io_out_0t[28]), .I0_f(ctrl_io_out_0f[28]), .T(ctrl_io_oeb[28]));
(* keep, BEL="X38Y30.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io29_i (.Q0_t(ctrl_io_in_0t[29]), .Q0_f(ctrl_io_in_0f[29]), .I0_t(ctrl_io_out_0t[29]), .I0_f(ctrl_io_out_0f[29]), .T(ctrl_io_oeb[29]));
(* keep, BEL="X38Y31.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io30_i (.Q0_t(ctrl_io_in_0t[30]), .Q0_f(ctrl_io_in_0f[30]), .I0_t(ctrl_io_out_0t[30]), .I0_f(ctrl_io_out_0f[30]), .T(ctrl_io_oeb[30]));
(* keep, BEL="X38Y32.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io31_i (.Q0_t(ctrl_io_in_0t[31]), .Q0_f(ctrl_io_in_0f[31]), .I0_t(ctrl_io_out_0t[31]), .I0_f(ctrl_io_out_0f[31]), .T(ctrl_io_oeb[31]));
(* keep, BEL="X38Y33.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io32_i (.Q0_t(ctrl_io_in_0t[32]), .Q0_f(ctrl_io_in_0f[32]), .I0_t(ctrl_io_out_0t[32]), .I0_f(ctrl_io_out_0f[32]), .T(ctrl_io_oeb[32]));
(* keep, BEL="X38Y34.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io33_i (.Q0_t(ctrl_io_in_0t[33]), .Q0_f(ctrl_io_in_0f[33]), .I0_t(ctrl_io_out_0t[33]), .I0_f(ctrl_io_out_0f[33]), .T(ctrl_io_oeb[33]));
(* keep, BEL="X38Y35.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io34_i (.Q0_t(ctrl_io_in_0t[34]), .Q0_f(ctrl_io_in_0f[34]), .I0_t(ctrl_io_out_0t[34]), .I0_f(ctrl_io_out_0f[34]), .T(ctrl_io_oeb[34]));
(* keep, BEL="X38Y36.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io35_i (.Q0_t(ctrl_io_in_0t[35]), .Q0_f(ctrl_io_in_0f[35]), .I0_t(ctrl_io_out_0t[35]), .I0_f(ctrl_io_out_0f[35]), .T(ctrl_io_oeb[35]));
(* keep, BEL="X38Y37.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io36_i (.Q0_t(ctrl_io_in_0t[36]), .Q0_f(ctrl_io_in_0f[36]), .I0_t(ctrl_io_out_0t[36]), .I0_f(ctrl_io_out_0f[36]), .T(ctrl_io_oeb[36]));
(* keep, BEL="X38Y38.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io37_i (.Q0_t(ctrl_io_in_0t[37]), .Q0_f(ctrl_io_in_0f[37]), .I0_t(ctrl_io_out_0t[37]), .I0_f(ctrl_io_out_0f[37]), .T(ctrl_io_oeb[37]));
(* keep, BEL="X38Y39.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io38_i (.Q0_t(ctrl_io_in_0t[38]), .Q0_f(ctrl_io_in_0f[38]), .I0_t(ctrl_io_out_0t[38]), .I0_f(ctrl_io_out_0f[38]), .T(ctrl_io_oeb[38]));
(* keep, BEL="X38Y40.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io39_i (.Q0_t(ctrl_io_in_0t[39]), .Q0_f(ctrl_io_in_0f[39]), .I0_t(ctrl_io_out_0t[39]), .I0_f(ctrl_io_out_0f[39]), .T(ctrl_io_oeb[39]));
(* keep, BEL="X38Y41.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io40_i (.Q0_t(ctrl_io_in_0t[40]), .Q0_f(ctrl_io_in_0f[40]), .I0_t(ctrl_io_out_0t[40]), .I0_f(ctrl_io_out_0f[40]), .T(ctrl_io_oeb[40]));
(* keep, BEL="X38Y42.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io41_i (.Q0_t(ctrl_io_in_0t[41]), .Q0_f(ctrl_io_in_0f[41]), .I0_t(ctrl_io_out_0t[41]), .I0_f(ctrl_io_out_0f[41]), .T(ctrl_io_oeb[41]));
(* keep, BEL="X38Y43.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io42_i (.Q0_t(ctrl_io_in_0t[42]), .Q0_f(ctrl_io_in_0f[42]), .I0_t(ctrl_io_out_0t[42]), .I0_f(ctrl_io_out_0f[42]), .T(ctrl_io_oeb[42]));
(* keep, BEL="X38Y44.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io43_i (.Q0_t(ctrl_io_in_0t[43]), .Q0_f(ctrl_io_in_0f[43]), .I0_t(ctrl_io_out_0t[43]), .I0_f(ctrl_io_out_0f[43]), .T(ctrl_io_oeb[43]));
(* keep, BEL="X38Y45.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io44_i (.Q0_t(ctrl_io_in_0t[44]), .Q0_f(ctrl_io_in_0f[44]), .I0_t(ctrl_io_out_0t[44]), .I0_f(ctrl_io_out_0f[44]), .T(ctrl_io_oeb[44]));
(* keep, BEL="X38Y46.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io45_i (.Q0_t(ctrl_io_in_0t[45]), .Q0_f(ctrl_io_in_0f[45]), .I0_t(ctrl_io_out_0t[45]), .I0_f(ctrl_io_out_0f[45]), .T(ctrl_io_oeb[45]));
(* keep, BEL="X38Y47.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io46_i (.Q0_t(ctrl_io_in_0t[46]), .Q0_f(ctrl_io_in_0f[46]), .I0_t(ctrl_io_out_0t[46]), .I0_f(ctrl_io_out_0f[46]), .T(ctrl_io_oeb[46]));
(* keep, BEL="X38Y48.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io47_i (.Q0_t(ctrl_io_in_0t[47]), .Q0_f(ctrl_io_in_0f[47]), .I0_t(ctrl_io_out_0t[47]), .I0_f(ctrl_io_out_0f[47]), .T(ctrl_io_oeb[47]));
(* keep, BEL="X38Y49.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io48_i (.Q0_t(ctrl_io_in_0t[48]), .Q0_f(ctrl_io_in_0f[48]), .I0_t(ctrl_io_out_0t[48]), .I0_f(ctrl_io_out_0f[48]), .T(ctrl_io_oeb[48]));
(* keep, BEL="X38Y50.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io49_i (.Q0_t(ctrl_io_in_0t[49]), .Q0_f(ctrl_io_in_0f[49]), .I0_t(ctrl_io_out_0t[49]), .I0_f(ctrl_io_out_0f[49]), .T(ctrl_io_oeb[49]));
(* keep, BEL="X38Y51.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io50_i (.Q0_t(ctrl_io_in_0t[50]), .Q0_f(ctrl_io_in_0f[50]), .I0_t(ctrl_io_out_0t[50]), .I0_f(ctrl_io_out_0f[50]), .T(ctrl_io_oeb[50]));
(* keep, BEL="X38Y52.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io51_i (.Q0_t(ctrl_io_in_0t[51]), .Q0_f(ctrl_io_in_0f[51]), .I0_t(ctrl_io_out_0t[51]), .I0_f(ctrl_io_out_0f[51]), .T(ctrl_io_oeb[51]));
(* keep, BEL="X38Y53.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io52_i (.Q0_t(ctrl_io_in_0t[52]), .Q0_f(ctrl_io_in_0f[52]), .I0_t(ctrl_io_out_0t[52]), .I0_f(ctrl_io_out_0f[52]), .T(ctrl_io_oeb[52]));
(* keep, BEL="X38Y54.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io53_i (.Q0_t(ctrl_io_in_0t[53]), .Q0_f(ctrl_io_in_0f[53]), .I0_t(ctrl_io_out_0t[53]), .I0_f(ctrl_io_out_0f[53]), .T(ctrl_io_oeb[53]));
(* keep, BEL="X38Y55.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io54_i (.Q0_t(ctrl_io_in_0t[54]), .Q0_f(ctrl_io_in_0f[54]), .I0_t(ctrl_io_out_0t[54]), .I0_f(ctrl_io_out_0f[54]), .T(ctrl_io_oeb[54]));
(* keep, BEL="X38Y56.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io55_i (.Q0_t(ctrl_io_in_0t[55]), .Q0_f(ctrl_io_in_0f[55]), .I0_t(ctrl_io_out_0t[55]), .I0_f(ctrl_io_out_0f[55]), .T(ctrl_io_oeb[55]));
(* keep, BEL="X38Y57.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io56_i (.Q0_t(ctrl_io_in_0t[56]), .Q0_f(ctrl_io_in_0f[56]), .I0_t(ctrl_io_out_0t[56]), .I0_f(ctrl_io_out_0f[56]), .T(ctrl_io_oeb[56]));
(* keep, BEL="X38Y58.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io57_i (.Q0_t(ctrl_io_in_0t[57]), .Q0_f(ctrl_io_in_0f[57]), .I0_t(ctrl_io_out_0t[57]), .I0_f(ctrl_io_out_0f[57]), .T(ctrl_io_oeb[57]));
(* keep, BEL="X38Y59.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io58_i (.Q0_t(ctrl_io_in_0t[58]), .Q0_f(ctrl_io_in_0f[58]), .I0_t(ctrl_io_out_0t[58]), .I0_f(ctrl_io_out_0f[58]), .T(ctrl_io_oeb[58]));
(* keep, BEL="X38Y60.A" *) ctrl_IO_1_bidirectional_frame_config_pass ctrl_io59_i (.Q0_t(ctrl_io_in_0t[59]), .Q0_f(ctrl_io_in_0f[59]), .I0_t(ctrl_io_out_0t[59]), .I0_f(ctrl_io_out_0f[59]), .T(ctrl_io_oeb[59]));
 
 
top top_i(.io_in_0t(io_in_0t), .io_in_0f(io_in_0f), .io_in_1t(io_in_1t), .io_in_1f(io_in_1f), .io_out_0t(io_out_0t), .io_out_0f(io_out_0f), .io_out_1t(io_out_1t), .io_out_1f(io_out_1f), .io_oeb(io_oeb), .ctrl_io_in_0t(ctrl_io_in_0t), .ctrl_io_in_0f(ctrl_io_in_0f), .ctrl_io_out_0t(ctrl_io_out_0t), .ctrl_io_out_0f(ctrl_io_out_0f), .ctrl_io_oeb(ctrl_io_oeb));
endmodule
