/* modified netlist. Source: module Midori64 in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/13-Midori64_round_based_enc_dec_PortParallel/4-AGEMA/Midori64.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module Midori64_SAUBER_Pipeline_d1 (DataIn_s0_t, key_s0_t, reset_t, enc_dec_t, key_s0_f, key_s1_t, key_s1_f, reset_f, enc_dec_f, DataIn_s0_f, DataIn_s1_t, DataIn_s1_f, DataOut_s0_t, done_t, done_f, DataOut_s0_f, DataOut_s1_t, DataOut_s1_f);
    input [63:0] DataIn_s0_t ;
    input [127:0] key_s0_t ;
    input reset_t ;
    input enc_dec_t ;
    input [127:0] key_s0_f ;
    input [127:0] key_s1_t ;
    input [127:0] key_s1_f ;
    input reset_f ;
    input enc_dec_f ;
    input [63:0] DataIn_s0_f ;
    input [63:0] DataIn_s1_t ;
    input [63:0] DataIn_s1_f ;
    output [63:0] DataOut_s0_t ;
    output done_t ;
    output done_f ;
    output [63:0] DataOut_s0_f ;
    output [63:0] DataOut_s1_t ;
    output [63:0] DataOut_s1_f ;
    wire controller_n2 ;
    wire controller_n1 ;
    wire controller_roundCounter_n15 ;
    wire controller_roundCounter_n14 ;
    wire controller_roundCounter_n13 ;
    wire controller_roundCounter_n8 ;
    wire controller_roundCounter_n4 ;
    wire controller_roundCounter_n5 ;
    wire controller_roundCounter_n6 ;
    wire controller_roundCounter_N7 ;
    wire controller_roundCounter_U9_Y ;
    wire controller_roundCounter_U9_X ;
    wire controller_roundCounter_U11_Y ;
    wire controller_roundCounter_U11_X ;
    wire controller_roundCounter_U15_Y ;
    wire controller_roundCounter_U15_X ;
    wire Midori_rounds_n16 ;
    wire Midori_rounds_n15 ;
    wire Midori_rounds_n14 ;
    wire Midori_rounds_n13 ;
    wire Midori_rounds_n12 ;
    wire Midori_rounds_n11 ;
    wire Midori_rounds_n10 ;
    wire Midori_rounds_n9 ;
    wire Midori_rounds_n8 ;
    wire Midori_rounds_n7 ;
    wire Midori_rounds_n6 ;
    wire Midori_rounds_n5 ;
    wire Midori_rounds_n4 ;
    wire Midori_rounds_n3 ;
    wire Midori_rounds_n2 ;
    wire Midori_rounds_n1 ;
    wire Midori_rounds_constant_MUX_n139 ;
    wire Midori_rounds_constant_MUX_n138 ;
    wire Midori_rounds_constant_MUX_n137 ;
    wire Midori_rounds_constant_MUX_n136 ;
    wire Midori_rounds_constant_MUX_n134 ;
    wire Midori_rounds_constant_MUX_n133 ;
    wire Midori_rounds_constant_MUX_n132 ;
    wire Midori_rounds_constant_MUX_n131 ;
    wire Midori_rounds_constant_MUX_n130 ;
    wire Midori_rounds_constant_MUX_n129 ;
    wire Midori_rounds_constant_MUX_n128 ;
    wire Midori_rounds_constant_MUX_n126 ;
    wire Midori_rounds_constant_MUX_n125 ;
    wire Midori_rounds_constant_MUX_n124 ;
    wire Midori_rounds_constant_MUX_n123 ;
    wire Midori_rounds_constant_MUX_n122 ;
    wire Midori_rounds_constant_MUX_n120 ;
    wire Midori_rounds_constant_MUX_n119 ;
    wire Midori_rounds_constant_MUX_n118 ;
    wire Midori_rounds_constant_MUX_n117 ;
    wire Midori_rounds_constant_MUX_n116 ;
    wire Midori_rounds_constant_MUX_n115 ;
    wire Midori_rounds_constant_MUX_n114 ;
    wire Midori_rounds_constant_MUX_n113 ;
    wire Midori_rounds_constant_MUX_n110 ;
    wire Midori_rounds_constant_MUX_n109 ;
    wire Midori_rounds_constant_MUX_n108 ;
    wire Midori_rounds_constant_MUX_n107 ;
    wire Midori_rounds_constant_MUX_n106 ;
    wire Midori_rounds_constant_MUX_n104 ;
    wire Midori_rounds_constant_MUX_n103 ;
    wire Midori_rounds_constant_MUX_n102 ;
    wire Midori_rounds_constant_MUX_n101 ;
    wire Midori_rounds_constant_MUX_n100 ;
    wire Midori_rounds_constant_MUX_n99 ;
    wire Midori_rounds_constant_MUX_n98 ;
    wire Midori_rounds_constant_MUX_n97 ;
    wire Midori_rounds_constant_MUX_n96 ;
    wire Midori_rounds_constant_MUX_n95 ;
    wire Midori_rounds_constant_MUX_n94 ;
    wire Midori_rounds_constant_MUX_n93 ;
    wire Midori_rounds_constant_MUX_n92 ;
    wire Midori_rounds_constant_MUX_n91 ;
    wire Midori_rounds_constant_MUX_n88 ;
    wire Midori_rounds_constant_MUX_n86 ;
    wire Midori_rounds_constant_MUX_n85 ;
    wire Midori_rounds_constant_MUX_n84 ;
    wire Midori_rounds_constant_MUX_n83 ;
    wire Midori_rounds_constant_MUX_n82 ;
    wire Midori_rounds_constant_MUX_n81 ;
    wire Midori_rounds_constant_MUX_n80 ;
    wire Midori_rounds_constant_MUX_n79 ;
    wire Midori_rounds_constant_MUX_n78 ;
    wire Midori_rounds_constant_MUX_n77 ;
    wire Midori_rounds_constant_MUX_n76 ;
    wire Midori_rounds_constant_MUX_n75 ;
    wire Midori_rounds_constant_MUX_n74 ;
    wire Midori_rounds_constant_MUX_n73 ;
    wire Midori_rounds_constant_MUX_n72 ;
    wire Midori_rounds_constant_MUX_n70 ;
    wire Midori_rounds_constant_MUX_n69 ;
    wire Midori_rounds_constant_MUX_n68 ;
    wire Midori_rounds_constant_MUX_n66 ;
    wire Midori_rounds_constant_MUX_n64 ;
    wire Midori_rounds_constant_MUX_n62 ;
    wire Midori_rounds_constant_MUX_n61 ;
    wire Midori_rounds_constant_MUX_n60 ;
    wire Midori_rounds_constant_MUX_n59 ;
    wire Midori_rounds_constant_MUX_n58 ;
    wire Midori_rounds_constant_MUX_n57 ;
    wire Midori_rounds_constant_MUX_n56 ;
    wire Midori_rounds_constant_MUX_n55 ;
    wire Midori_rounds_constant_MUX_n54 ;
    wire Midori_rounds_constant_MUX_n53 ;
    wire Midori_rounds_constant_MUX_n52 ;
    wire Midori_rounds_constant_MUX_n51 ;
    wire Midori_rounds_constant_MUX_n50 ;
    wire Midori_rounds_constant_MUX_n49 ;
    wire Midori_rounds_constant_MUX_n48 ;
    wire Midori_rounds_constant_MUX_n47 ;
    wire Midori_rounds_constant_MUX_n46 ;
    wire Midori_rounds_constant_MUX_n42 ;
    wire Midori_rounds_constant_MUX_n40 ;
    wire Midori_rounds_constant_MUX_n37 ;
    wire Midori_rounds_constant_MUX_n36 ;
    wire Midori_rounds_constant_MUX_n35 ;
    wire Midori_rounds_constant_MUX_n34 ;
    wire Midori_rounds_constant_MUX_n33 ;
    wire Midori_rounds_constant_MUX_n32 ;
    wire Midori_rounds_constant_MUX_n31 ;
    wire Midori_rounds_constant_MUX_n30 ;
    wire Midori_rounds_constant_MUX_n29 ;
    wire Midori_rounds_constant_MUX_n28 ;
    wire Midori_rounds_constant_MUX_n27 ;
    wire Midori_rounds_constant_MUX_n25 ;
    wire Midori_rounds_constant_MUX_n24 ;
    wire Midori_rounds_constant_MUX_n23 ;
    wire Midori_rounds_constant_MUX_n22 ;
    wire Midori_rounds_constant_MUX_n121 ;
    wire Midori_rounds_constant_MUX_n112 ;
    wire Midori_rounds_constant_MUX_n43 ;
    wire Midori_rounds_constant_MUX_n111 ;
    wire Midori_rounds_constant_MUX_U53_Y ;
    wire Midori_rounds_constant_MUX_U53_X ;
    wire Midori_rounds_constant_MUX_U119_Y ;
    wire Midori_rounds_constant_MUX_U119_X ;
    wire Midori_rounds_MUXInst_mux_inst_0_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_0_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_1_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_1_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_2_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_2_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_3_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_3_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_4_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_4_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_5_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_5_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_6_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_6_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_7_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_7_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_8_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_8_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_9_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_9_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_10_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_10_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_11_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_11_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_12_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_12_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_13_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_13_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_14_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_14_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_15_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_15_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_16_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_16_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_17_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_17_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_18_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_18_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_19_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_19_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_20_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_20_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_21_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_21_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_22_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_22_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_23_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_23_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_24_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_24_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_25_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_25_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_26_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_26_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_27_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_27_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_28_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_28_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_29_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_29_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_30_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_30_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_31_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_31_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_32_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_32_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_33_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_33_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_34_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_34_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_35_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_35_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_36_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_36_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_37_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_37_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_38_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_38_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_39_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_39_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_40_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_40_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_41_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_41_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_42_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_42_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_43_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_43_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_44_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_44_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_45_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_45_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_46_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_46_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_47_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_47_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_48_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_48_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_49_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_49_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_50_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_50_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_51_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_51_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_52_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_52_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_53_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_53_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_54_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_54_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_55_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_55_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_56_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_56_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_57_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_57_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_58_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_58_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_59_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_59_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_60_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_60_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_61_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_61_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_62_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_62_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_63_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_63_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_X ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n1 ;
    wire Midori_rounds_mul_input_Inst_mux_inst_0_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_0_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_1_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_1_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_2_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_2_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_3_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_3_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_4_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_4_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_5_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_5_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_6_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_6_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_7_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_7_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_8_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_8_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_9_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_9_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_10_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_10_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_11_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_11_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_12_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_12_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_13_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_13_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_14_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_14_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_15_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_15_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_16_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_16_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_17_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_17_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_18_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_18_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_19_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_19_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_20_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_20_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_21_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_21_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_22_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_22_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_23_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_23_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_24_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_24_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_25_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_25_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_26_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_26_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_27_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_27_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_28_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_28_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_29_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_29_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_30_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_30_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_31_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_31_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_32_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_32_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_33_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_33_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_34_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_34_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_35_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_35_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_36_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_36_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_37_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_37_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_38_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_38_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_39_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_39_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_40_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_40_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_41_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_41_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_42_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_42_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_43_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_43_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_44_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_44_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_45_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_45_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_46_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_46_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_47_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_47_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_48_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_48_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_49_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_49_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_50_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_50_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_51_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_51_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_52_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_52_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_53_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_53_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_54_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_54_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_55_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_55_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_56_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_56_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_57_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_57_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_58_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_58_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_59_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_59_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_60_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_60_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_61_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_61_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_62_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_62_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_63_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_63_U1_X ;
    wire Midori_rounds_mul_MC1_n8 ;
    wire Midori_rounds_mul_MC1_n7 ;
    wire Midori_rounds_mul_MC1_n6 ;
    wire Midori_rounds_mul_MC1_n5 ;
    wire Midori_rounds_mul_MC1_n4 ;
    wire Midori_rounds_mul_MC1_n3 ;
    wire Midori_rounds_mul_MC1_n2 ;
    wire Midori_rounds_mul_MC1_n1 ;
    wire Midori_rounds_mul_MC2_n8 ;
    wire Midori_rounds_mul_MC2_n7 ;
    wire Midori_rounds_mul_MC2_n6 ;
    wire Midori_rounds_mul_MC2_n5 ;
    wire Midori_rounds_mul_MC2_n4 ;
    wire Midori_rounds_mul_MC2_n3 ;
    wire Midori_rounds_mul_MC2_n2 ;
    wire Midori_rounds_mul_MC2_n1 ;
    wire Midori_rounds_mul_MC3_n8 ;
    wire Midori_rounds_mul_MC3_n7 ;
    wire Midori_rounds_mul_MC3_n6 ;
    wire Midori_rounds_mul_MC3_n5 ;
    wire Midori_rounds_mul_MC3_n4 ;
    wire Midori_rounds_mul_MC3_n3 ;
    wire Midori_rounds_mul_MC3_n2 ;
    wire Midori_rounds_mul_MC3_n1 ;
    wire Midori_rounds_mul_MC4_n8 ;
    wire Midori_rounds_mul_MC4_n7 ;
    wire Midori_rounds_mul_MC4_n6 ;
    wire Midori_rounds_mul_MC4_n5 ;
    wire Midori_rounds_mul_MC4_n4 ;
    wire Midori_rounds_mul_MC4_n3 ;
    wire Midori_rounds_mul_MC4_n2 ;
    wire Midori_rounds_mul_MC4_n1 ;
    wire Midori_rounds_Res_Inst_mux_inst_0_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_0_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_1_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_1_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_2_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_2_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_3_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_3_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_4_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_4_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_5_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_5_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_6_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_6_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_7_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_7_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_8_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_8_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_9_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_9_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_10_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_10_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_11_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_11_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_12_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_12_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_13_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_13_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_14_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_14_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_15_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_15_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_16_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_16_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_17_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_17_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_18_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_18_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_19_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_19_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_20_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_20_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_21_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_21_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_22_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_22_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_23_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_23_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_24_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_24_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_25_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_25_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_26_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_26_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_27_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_27_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_28_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_28_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_29_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_29_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_30_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_30_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_31_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_31_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_32_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_32_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_33_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_33_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_34_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_34_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_35_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_35_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_36_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_36_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_37_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_37_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_38_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_38_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_39_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_39_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_40_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_40_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_41_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_41_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_42_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_42_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_43_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_43_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_44_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_44_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_45_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_45_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_46_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_46_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_47_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_47_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_48_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_48_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_49_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_49_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_50_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_50_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_51_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_51_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_52_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_52_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_53_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_53_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_54_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_54_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_55_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_55_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_56_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_56_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_57_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_57_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_58_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_58_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_59_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_59_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_60_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_60_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_61_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_61_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_62_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_62_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_63_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_63_U1_X ;
    wire [63:0] wk ;
    wire [3:0] round_Signal ;
    wire [63:0] Midori_add_Result_Start ;
    wire [63:0] Midori_rounds_mul_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Inv_Result ;
    wire [63:0] Midori_rounds_mul_input ;
    wire [63:0] Midori_rounds_sub_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Result ;
    wire [63:0] Midori_rounds_roundReg_out ;
    wire [63:0] Midori_rounds_round_Result ;
    wire [63:0] Midori_rounds_SelectedKey ;
    wire [15:0] Midori_rounds_round_Constant ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;

    /* cells in depth 0 */
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U64 ( .A0_t (key_s0_t[127]), .A0_f (key_s0_f[127]), .A1_t (key_s1_t[127]), .A1_f (key_s1_f[127]), .B0_t (key_s0_t[63]), .B0_f (key_s0_f[63]), .B1_t (key_s1_t[63]), .B1_f (key_s1_f[63]), .Z0_t (wk[63]), .Z0_f (new_AGEMA_signal_2011), .Z1_t (new_AGEMA_signal_2012), .Z1_f (new_AGEMA_signal_2013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U63 ( .A0_t (key_s0_t[126]), .A0_f (key_s0_f[126]), .A1_t (key_s1_t[126]), .A1_f (key_s1_f[126]), .B0_t (key_s0_t[62]), .B0_f (key_s0_f[62]), .B1_t (key_s1_t[62]), .B1_f (key_s1_f[62]), .Z0_t (wk[62]), .Z0_f (new_AGEMA_signal_2020), .Z1_t (new_AGEMA_signal_2021), .Z1_f (new_AGEMA_signal_2022) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U62 ( .A0_t (key_s0_t[125]), .A0_f (key_s0_f[125]), .A1_t (key_s1_t[125]), .A1_f (key_s1_f[125]), .B0_t (key_s0_t[61]), .B0_f (key_s0_f[61]), .B1_t (key_s1_t[61]), .B1_f (key_s1_f[61]), .Z0_t (wk[61]), .Z0_f (new_AGEMA_signal_2029), .Z1_t (new_AGEMA_signal_2030), .Z1_f (new_AGEMA_signal_2031) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U61 ( .A0_t (key_s0_t[124]), .A0_f (key_s0_f[124]), .A1_t (key_s1_t[124]), .A1_f (key_s1_f[124]), .B0_t (key_s0_t[60]), .B0_f (key_s0_f[60]), .B1_t (key_s1_t[60]), .B1_f (key_s1_f[60]), .Z0_t (wk[60]), .Z0_f (new_AGEMA_signal_2038), .Z1_t (new_AGEMA_signal_2039), .Z1_f (new_AGEMA_signal_2040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U60 ( .A0_t (key_s0_t[123]), .A0_f (key_s0_f[123]), .A1_t (key_s1_t[123]), .A1_f (key_s1_f[123]), .B0_t (key_s0_t[59]), .B0_f (key_s0_f[59]), .B1_t (key_s1_t[59]), .B1_f (key_s1_f[59]), .Z0_t (wk[59]), .Z0_f (new_AGEMA_signal_2047), .Z1_t (new_AGEMA_signal_2048), .Z1_f (new_AGEMA_signal_2049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U59 ( .A0_t (key_s0_t[122]), .A0_f (key_s0_f[122]), .A1_t (key_s1_t[122]), .A1_f (key_s1_f[122]), .B0_t (key_s0_t[58]), .B0_f (key_s0_f[58]), .B1_t (key_s1_t[58]), .B1_f (key_s1_f[58]), .Z0_t (wk[58]), .Z0_f (new_AGEMA_signal_2056), .Z1_t (new_AGEMA_signal_2057), .Z1_f (new_AGEMA_signal_2058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U58 ( .A0_t (key_s0_t[121]), .A0_f (key_s0_f[121]), .A1_t (key_s1_t[121]), .A1_f (key_s1_f[121]), .B0_t (key_s0_t[57]), .B0_f (key_s0_f[57]), .B1_t (key_s1_t[57]), .B1_f (key_s1_f[57]), .Z0_t (wk[57]), .Z0_f (new_AGEMA_signal_2065), .Z1_t (new_AGEMA_signal_2066), .Z1_f (new_AGEMA_signal_2067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U57 ( .A0_t (key_s0_t[120]), .A0_f (key_s0_f[120]), .A1_t (key_s1_t[120]), .A1_f (key_s1_f[120]), .B0_t (key_s0_t[56]), .B0_f (key_s0_f[56]), .B1_t (key_s1_t[56]), .B1_f (key_s1_f[56]), .Z0_t (wk[56]), .Z0_f (new_AGEMA_signal_2074), .Z1_t (new_AGEMA_signal_2075), .Z1_f (new_AGEMA_signal_2076) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U56 ( .A0_t (key_s0_t[119]), .A0_f (key_s0_f[119]), .A1_t (key_s1_t[119]), .A1_f (key_s1_f[119]), .B0_t (key_s0_t[55]), .B0_f (key_s0_f[55]), .B1_t (key_s1_t[55]), .B1_f (key_s1_f[55]), .Z0_t (wk[55]), .Z0_f (new_AGEMA_signal_2083), .Z1_t (new_AGEMA_signal_2084), .Z1_f (new_AGEMA_signal_2085) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U55 ( .A0_t (key_s0_t[118]), .A0_f (key_s0_f[118]), .A1_t (key_s1_t[118]), .A1_f (key_s1_f[118]), .B0_t (key_s0_t[54]), .B0_f (key_s0_f[54]), .B1_t (key_s1_t[54]), .B1_f (key_s1_f[54]), .Z0_t (wk[54]), .Z0_f (new_AGEMA_signal_2092), .Z1_t (new_AGEMA_signal_2093), .Z1_f (new_AGEMA_signal_2094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U54 ( .A0_t (key_s0_t[117]), .A0_f (key_s0_f[117]), .A1_t (key_s1_t[117]), .A1_f (key_s1_f[117]), .B0_t (key_s0_t[53]), .B0_f (key_s0_f[53]), .B1_t (key_s1_t[53]), .B1_f (key_s1_f[53]), .Z0_t (wk[53]), .Z0_f (new_AGEMA_signal_2101), .Z1_t (new_AGEMA_signal_2102), .Z1_f (new_AGEMA_signal_2103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U53 ( .A0_t (key_s0_t[116]), .A0_f (key_s0_f[116]), .A1_t (key_s1_t[116]), .A1_f (key_s1_f[116]), .B0_t (key_s0_t[52]), .B0_f (key_s0_f[52]), .B1_t (key_s1_t[52]), .B1_f (key_s1_f[52]), .Z0_t (wk[52]), .Z0_f (new_AGEMA_signal_2110), .Z1_t (new_AGEMA_signal_2111), .Z1_f (new_AGEMA_signal_2112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U52 ( .A0_t (key_s0_t[115]), .A0_f (key_s0_f[115]), .A1_t (key_s1_t[115]), .A1_f (key_s1_f[115]), .B0_t (key_s0_t[51]), .B0_f (key_s0_f[51]), .B1_t (key_s1_t[51]), .B1_f (key_s1_f[51]), .Z0_t (wk[51]), .Z0_f (new_AGEMA_signal_2119), .Z1_t (new_AGEMA_signal_2120), .Z1_f (new_AGEMA_signal_2121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U51 ( .A0_t (key_s0_t[114]), .A0_f (key_s0_f[114]), .A1_t (key_s1_t[114]), .A1_f (key_s1_f[114]), .B0_t (key_s0_t[50]), .B0_f (key_s0_f[50]), .B1_t (key_s1_t[50]), .B1_f (key_s1_f[50]), .Z0_t (wk[50]), .Z0_f (new_AGEMA_signal_2128), .Z1_t (new_AGEMA_signal_2129), .Z1_f (new_AGEMA_signal_2130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U50 ( .A0_t (key_s0_t[113]), .A0_f (key_s0_f[113]), .A1_t (key_s1_t[113]), .A1_f (key_s1_f[113]), .B0_t (key_s0_t[49]), .B0_f (key_s0_f[49]), .B1_t (key_s1_t[49]), .B1_f (key_s1_f[49]), .Z0_t (wk[49]), .Z0_f (new_AGEMA_signal_2137), .Z1_t (new_AGEMA_signal_2138), .Z1_f (new_AGEMA_signal_2139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U49 ( .A0_t (key_s0_t[112]), .A0_f (key_s0_f[112]), .A1_t (key_s1_t[112]), .A1_f (key_s1_f[112]), .B0_t (key_s0_t[48]), .B0_f (key_s0_f[48]), .B1_t (key_s1_t[48]), .B1_f (key_s1_f[48]), .Z0_t (wk[48]), .Z0_f (new_AGEMA_signal_2146), .Z1_t (new_AGEMA_signal_2147), .Z1_f (new_AGEMA_signal_2148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U48 ( .A0_t (key_s0_t[111]), .A0_f (key_s0_f[111]), .A1_t (key_s1_t[111]), .A1_f (key_s1_f[111]), .B0_t (key_s0_t[47]), .B0_f (key_s0_f[47]), .B1_t (key_s1_t[47]), .B1_f (key_s1_f[47]), .Z0_t (wk[47]), .Z0_f (new_AGEMA_signal_2155), .Z1_t (new_AGEMA_signal_2156), .Z1_f (new_AGEMA_signal_2157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U47 ( .A0_t (key_s0_t[110]), .A0_f (key_s0_f[110]), .A1_t (key_s1_t[110]), .A1_f (key_s1_f[110]), .B0_t (key_s0_t[46]), .B0_f (key_s0_f[46]), .B1_t (key_s1_t[46]), .B1_f (key_s1_f[46]), .Z0_t (wk[46]), .Z0_f (new_AGEMA_signal_2164), .Z1_t (new_AGEMA_signal_2165), .Z1_f (new_AGEMA_signal_2166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U46 ( .A0_t (key_s0_t[109]), .A0_f (key_s0_f[109]), .A1_t (key_s1_t[109]), .A1_f (key_s1_f[109]), .B0_t (key_s0_t[45]), .B0_f (key_s0_f[45]), .B1_t (key_s1_t[45]), .B1_f (key_s1_f[45]), .Z0_t (wk[45]), .Z0_f (new_AGEMA_signal_2173), .Z1_t (new_AGEMA_signal_2174), .Z1_f (new_AGEMA_signal_2175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U45 ( .A0_t (key_s0_t[108]), .A0_f (key_s0_f[108]), .A1_t (key_s1_t[108]), .A1_f (key_s1_f[108]), .B0_t (key_s0_t[44]), .B0_f (key_s0_f[44]), .B1_t (key_s1_t[44]), .B1_f (key_s1_f[44]), .Z0_t (wk[44]), .Z0_f (new_AGEMA_signal_2182), .Z1_t (new_AGEMA_signal_2183), .Z1_f (new_AGEMA_signal_2184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U44 ( .A0_t (key_s0_t[107]), .A0_f (key_s0_f[107]), .A1_t (key_s1_t[107]), .A1_f (key_s1_f[107]), .B0_t (key_s0_t[43]), .B0_f (key_s0_f[43]), .B1_t (key_s1_t[43]), .B1_f (key_s1_f[43]), .Z0_t (wk[43]), .Z0_f (new_AGEMA_signal_2191), .Z1_t (new_AGEMA_signal_2192), .Z1_f (new_AGEMA_signal_2193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U43 ( .A0_t (key_s0_t[106]), .A0_f (key_s0_f[106]), .A1_t (key_s1_t[106]), .A1_f (key_s1_f[106]), .B0_t (key_s0_t[42]), .B0_f (key_s0_f[42]), .B1_t (key_s1_t[42]), .B1_f (key_s1_f[42]), .Z0_t (wk[42]), .Z0_f (new_AGEMA_signal_2200), .Z1_t (new_AGEMA_signal_2201), .Z1_f (new_AGEMA_signal_2202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U42 ( .A0_t (key_s0_t[105]), .A0_f (key_s0_f[105]), .A1_t (key_s1_t[105]), .A1_f (key_s1_f[105]), .B0_t (key_s0_t[41]), .B0_f (key_s0_f[41]), .B1_t (key_s1_t[41]), .B1_f (key_s1_f[41]), .Z0_t (wk[41]), .Z0_f (new_AGEMA_signal_2209), .Z1_t (new_AGEMA_signal_2210), .Z1_f (new_AGEMA_signal_2211) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U41 ( .A0_t (key_s0_t[104]), .A0_f (key_s0_f[104]), .A1_t (key_s1_t[104]), .A1_f (key_s1_f[104]), .B0_t (key_s0_t[40]), .B0_f (key_s0_f[40]), .B1_t (key_s1_t[40]), .B1_f (key_s1_f[40]), .Z0_t (wk[40]), .Z0_f (new_AGEMA_signal_2218), .Z1_t (new_AGEMA_signal_2219), .Z1_f (new_AGEMA_signal_2220) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U40 ( .A0_t (key_s0_t[103]), .A0_f (key_s0_f[103]), .A1_t (key_s1_t[103]), .A1_f (key_s1_f[103]), .B0_t (key_s0_t[39]), .B0_f (key_s0_f[39]), .B1_t (key_s1_t[39]), .B1_f (key_s1_f[39]), .Z0_t (wk[39]), .Z0_f (new_AGEMA_signal_2227), .Z1_t (new_AGEMA_signal_2228), .Z1_f (new_AGEMA_signal_2229) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U39 ( .A0_t (key_s0_t[102]), .A0_f (key_s0_f[102]), .A1_t (key_s1_t[102]), .A1_f (key_s1_f[102]), .B0_t (key_s0_t[38]), .B0_f (key_s0_f[38]), .B1_t (key_s1_t[38]), .B1_f (key_s1_f[38]), .Z0_t (wk[38]), .Z0_f (new_AGEMA_signal_2236), .Z1_t (new_AGEMA_signal_2237), .Z1_f (new_AGEMA_signal_2238) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U38 ( .A0_t (key_s0_t[101]), .A0_f (key_s0_f[101]), .A1_t (key_s1_t[101]), .A1_f (key_s1_f[101]), .B0_t (key_s0_t[37]), .B0_f (key_s0_f[37]), .B1_t (key_s1_t[37]), .B1_f (key_s1_f[37]), .Z0_t (wk[37]), .Z0_f (new_AGEMA_signal_2245), .Z1_t (new_AGEMA_signal_2246), .Z1_f (new_AGEMA_signal_2247) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U37 ( .A0_t (key_s0_t[100]), .A0_f (key_s0_f[100]), .A1_t (key_s1_t[100]), .A1_f (key_s1_f[100]), .B0_t (key_s0_t[36]), .B0_f (key_s0_f[36]), .B1_t (key_s1_t[36]), .B1_f (key_s1_f[36]), .Z0_t (wk[36]), .Z0_f (new_AGEMA_signal_2254), .Z1_t (new_AGEMA_signal_2255), .Z1_f (new_AGEMA_signal_2256) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U36 ( .A0_t (key_s0_t[99]), .A0_f (key_s0_f[99]), .A1_t (key_s1_t[99]), .A1_f (key_s1_f[99]), .B0_t (key_s0_t[35]), .B0_f (key_s0_f[35]), .B1_t (key_s1_t[35]), .B1_f (key_s1_f[35]), .Z0_t (wk[35]), .Z0_f (new_AGEMA_signal_2263), .Z1_t (new_AGEMA_signal_2264), .Z1_f (new_AGEMA_signal_2265) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U35 ( .A0_t (key_s0_t[98]), .A0_f (key_s0_f[98]), .A1_t (key_s1_t[98]), .A1_f (key_s1_f[98]), .B0_t (key_s0_t[34]), .B0_f (key_s0_f[34]), .B1_t (key_s1_t[34]), .B1_f (key_s1_f[34]), .Z0_t (wk[34]), .Z0_f (new_AGEMA_signal_2272), .Z1_t (new_AGEMA_signal_2273), .Z1_f (new_AGEMA_signal_2274) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U34 ( .A0_t (key_s0_t[97]), .A0_f (key_s0_f[97]), .A1_t (key_s1_t[97]), .A1_f (key_s1_f[97]), .B0_t (key_s0_t[33]), .B0_f (key_s0_f[33]), .B1_t (key_s1_t[33]), .B1_f (key_s1_f[33]), .Z0_t (wk[33]), .Z0_f (new_AGEMA_signal_2281), .Z1_t (new_AGEMA_signal_2282), .Z1_f (new_AGEMA_signal_2283) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U33 ( .A0_t (key_s0_t[96]), .A0_f (key_s0_f[96]), .A1_t (key_s1_t[96]), .A1_f (key_s1_f[96]), .B0_t (key_s0_t[32]), .B0_f (key_s0_f[32]), .B1_t (key_s1_t[32]), .B1_f (key_s1_f[32]), .Z0_t (wk[32]), .Z0_f (new_AGEMA_signal_2290), .Z1_t (new_AGEMA_signal_2291), .Z1_f (new_AGEMA_signal_2292) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U32 ( .A0_t (key_s0_t[95]), .A0_f (key_s0_f[95]), .A1_t (key_s1_t[95]), .A1_f (key_s1_f[95]), .B0_t (key_s0_t[31]), .B0_f (key_s0_f[31]), .B1_t (key_s1_t[31]), .B1_f (key_s1_f[31]), .Z0_t (wk[31]), .Z0_f (new_AGEMA_signal_2299), .Z1_t (new_AGEMA_signal_2300), .Z1_f (new_AGEMA_signal_2301) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U31 ( .A0_t (key_s0_t[94]), .A0_f (key_s0_f[94]), .A1_t (key_s1_t[94]), .A1_f (key_s1_f[94]), .B0_t (key_s0_t[30]), .B0_f (key_s0_f[30]), .B1_t (key_s1_t[30]), .B1_f (key_s1_f[30]), .Z0_t (wk[30]), .Z0_f (new_AGEMA_signal_2308), .Z1_t (new_AGEMA_signal_2309), .Z1_f (new_AGEMA_signal_2310) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U30 ( .A0_t (key_s0_t[93]), .A0_f (key_s0_f[93]), .A1_t (key_s1_t[93]), .A1_f (key_s1_f[93]), .B0_t (key_s0_t[29]), .B0_f (key_s0_f[29]), .B1_t (key_s1_t[29]), .B1_f (key_s1_f[29]), .Z0_t (wk[29]), .Z0_f (new_AGEMA_signal_2317), .Z1_t (new_AGEMA_signal_2318), .Z1_f (new_AGEMA_signal_2319) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U29 ( .A0_t (key_s0_t[92]), .A0_f (key_s0_f[92]), .A1_t (key_s1_t[92]), .A1_f (key_s1_f[92]), .B0_t (key_s0_t[28]), .B0_f (key_s0_f[28]), .B1_t (key_s1_t[28]), .B1_f (key_s1_f[28]), .Z0_t (wk[28]), .Z0_f (new_AGEMA_signal_2326), .Z1_t (new_AGEMA_signal_2327), .Z1_f (new_AGEMA_signal_2328) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U28 ( .A0_t (key_s0_t[91]), .A0_f (key_s0_f[91]), .A1_t (key_s1_t[91]), .A1_f (key_s1_f[91]), .B0_t (key_s0_t[27]), .B0_f (key_s0_f[27]), .B1_t (key_s1_t[27]), .B1_f (key_s1_f[27]), .Z0_t (wk[27]), .Z0_f (new_AGEMA_signal_2335), .Z1_t (new_AGEMA_signal_2336), .Z1_f (new_AGEMA_signal_2337) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U27 ( .A0_t (key_s0_t[90]), .A0_f (key_s0_f[90]), .A1_t (key_s1_t[90]), .A1_f (key_s1_f[90]), .B0_t (key_s0_t[26]), .B0_f (key_s0_f[26]), .B1_t (key_s1_t[26]), .B1_f (key_s1_f[26]), .Z0_t (wk[26]), .Z0_f (new_AGEMA_signal_2344), .Z1_t (new_AGEMA_signal_2345), .Z1_f (new_AGEMA_signal_2346) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U26 ( .A0_t (key_s0_t[89]), .A0_f (key_s0_f[89]), .A1_t (key_s1_t[89]), .A1_f (key_s1_f[89]), .B0_t (key_s0_t[25]), .B0_f (key_s0_f[25]), .B1_t (key_s1_t[25]), .B1_f (key_s1_f[25]), .Z0_t (wk[25]), .Z0_f (new_AGEMA_signal_2353), .Z1_t (new_AGEMA_signal_2354), .Z1_f (new_AGEMA_signal_2355) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U25 ( .A0_t (key_s0_t[88]), .A0_f (key_s0_f[88]), .A1_t (key_s1_t[88]), .A1_f (key_s1_f[88]), .B0_t (key_s0_t[24]), .B0_f (key_s0_f[24]), .B1_t (key_s1_t[24]), .B1_f (key_s1_f[24]), .Z0_t (wk[24]), .Z0_f (new_AGEMA_signal_2362), .Z1_t (new_AGEMA_signal_2363), .Z1_f (new_AGEMA_signal_2364) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U24 ( .A0_t (key_s0_t[87]), .A0_f (key_s0_f[87]), .A1_t (key_s1_t[87]), .A1_f (key_s1_f[87]), .B0_t (key_s0_t[23]), .B0_f (key_s0_f[23]), .B1_t (key_s1_t[23]), .B1_f (key_s1_f[23]), .Z0_t (wk[23]), .Z0_f (new_AGEMA_signal_2371), .Z1_t (new_AGEMA_signal_2372), .Z1_f (new_AGEMA_signal_2373) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U23 ( .A0_t (key_s0_t[86]), .A0_f (key_s0_f[86]), .A1_t (key_s1_t[86]), .A1_f (key_s1_f[86]), .B0_t (key_s0_t[22]), .B0_f (key_s0_f[22]), .B1_t (key_s1_t[22]), .B1_f (key_s1_f[22]), .Z0_t (wk[22]), .Z0_f (new_AGEMA_signal_2380), .Z1_t (new_AGEMA_signal_2381), .Z1_f (new_AGEMA_signal_2382) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U22 ( .A0_t (key_s0_t[85]), .A0_f (key_s0_f[85]), .A1_t (key_s1_t[85]), .A1_f (key_s1_f[85]), .B0_t (key_s0_t[21]), .B0_f (key_s0_f[21]), .B1_t (key_s1_t[21]), .B1_f (key_s1_f[21]), .Z0_t (wk[21]), .Z0_f (new_AGEMA_signal_2389), .Z1_t (new_AGEMA_signal_2390), .Z1_f (new_AGEMA_signal_2391) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U21 ( .A0_t (key_s0_t[84]), .A0_f (key_s0_f[84]), .A1_t (key_s1_t[84]), .A1_f (key_s1_f[84]), .B0_t (key_s0_t[20]), .B0_f (key_s0_f[20]), .B1_t (key_s1_t[20]), .B1_f (key_s1_f[20]), .Z0_t (wk[20]), .Z0_f (new_AGEMA_signal_2398), .Z1_t (new_AGEMA_signal_2399), .Z1_f (new_AGEMA_signal_2400) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U20 ( .A0_t (key_s0_t[83]), .A0_f (key_s0_f[83]), .A1_t (key_s1_t[83]), .A1_f (key_s1_f[83]), .B0_t (key_s0_t[19]), .B0_f (key_s0_f[19]), .B1_t (key_s1_t[19]), .B1_f (key_s1_f[19]), .Z0_t (wk[19]), .Z0_f (new_AGEMA_signal_2407), .Z1_t (new_AGEMA_signal_2408), .Z1_f (new_AGEMA_signal_2409) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U19 ( .A0_t (key_s0_t[82]), .A0_f (key_s0_f[82]), .A1_t (key_s1_t[82]), .A1_f (key_s1_f[82]), .B0_t (key_s0_t[18]), .B0_f (key_s0_f[18]), .B1_t (key_s1_t[18]), .B1_f (key_s1_f[18]), .Z0_t (wk[18]), .Z0_f (new_AGEMA_signal_2416), .Z1_t (new_AGEMA_signal_2417), .Z1_f (new_AGEMA_signal_2418) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U18 ( .A0_t (key_s0_t[81]), .A0_f (key_s0_f[81]), .A1_t (key_s1_t[81]), .A1_f (key_s1_f[81]), .B0_t (key_s0_t[17]), .B0_f (key_s0_f[17]), .B1_t (key_s1_t[17]), .B1_f (key_s1_f[17]), .Z0_t (wk[17]), .Z0_f (new_AGEMA_signal_2425), .Z1_t (new_AGEMA_signal_2426), .Z1_f (new_AGEMA_signal_2427) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U17 ( .A0_t (key_s0_t[80]), .A0_f (key_s0_f[80]), .A1_t (key_s1_t[80]), .A1_f (key_s1_f[80]), .B0_t (key_s0_t[16]), .B0_f (key_s0_f[16]), .B1_t (key_s1_t[16]), .B1_f (key_s1_f[16]), .Z0_t (wk[16]), .Z0_f (new_AGEMA_signal_2434), .Z1_t (new_AGEMA_signal_2435), .Z1_f (new_AGEMA_signal_2436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U16 ( .A0_t (key_s0_t[79]), .A0_f (key_s0_f[79]), .A1_t (key_s1_t[79]), .A1_f (key_s1_f[79]), .B0_t (key_s0_t[15]), .B0_f (key_s0_f[15]), .B1_t (key_s1_t[15]), .B1_f (key_s1_f[15]), .Z0_t (wk[15]), .Z0_f (new_AGEMA_signal_2443), .Z1_t (new_AGEMA_signal_2444), .Z1_f (new_AGEMA_signal_2445) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U15 ( .A0_t (key_s0_t[78]), .A0_f (key_s0_f[78]), .A1_t (key_s1_t[78]), .A1_f (key_s1_f[78]), .B0_t (key_s0_t[14]), .B0_f (key_s0_f[14]), .B1_t (key_s1_t[14]), .B1_f (key_s1_f[14]), .Z0_t (wk[14]), .Z0_f (new_AGEMA_signal_2452), .Z1_t (new_AGEMA_signal_2453), .Z1_f (new_AGEMA_signal_2454) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U14 ( .A0_t (key_s0_t[77]), .A0_f (key_s0_f[77]), .A1_t (key_s1_t[77]), .A1_f (key_s1_f[77]), .B0_t (key_s0_t[13]), .B0_f (key_s0_f[13]), .B1_t (key_s1_t[13]), .B1_f (key_s1_f[13]), .Z0_t (wk[13]), .Z0_f (new_AGEMA_signal_2461), .Z1_t (new_AGEMA_signal_2462), .Z1_f (new_AGEMA_signal_2463) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U13 ( .A0_t (key_s0_t[76]), .A0_f (key_s0_f[76]), .A1_t (key_s1_t[76]), .A1_f (key_s1_f[76]), .B0_t (key_s0_t[12]), .B0_f (key_s0_f[12]), .B1_t (key_s1_t[12]), .B1_f (key_s1_f[12]), .Z0_t (wk[12]), .Z0_f (new_AGEMA_signal_2470), .Z1_t (new_AGEMA_signal_2471), .Z1_f (new_AGEMA_signal_2472) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U12 ( .A0_t (key_s0_t[75]), .A0_f (key_s0_f[75]), .A1_t (key_s1_t[75]), .A1_f (key_s1_f[75]), .B0_t (key_s0_t[11]), .B0_f (key_s0_f[11]), .B1_t (key_s1_t[11]), .B1_f (key_s1_f[11]), .Z0_t (wk[11]), .Z0_f (new_AGEMA_signal_2479), .Z1_t (new_AGEMA_signal_2480), .Z1_f (new_AGEMA_signal_2481) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U11 ( .A0_t (key_s0_t[74]), .A0_f (key_s0_f[74]), .A1_t (key_s1_t[74]), .A1_f (key_s1_f[74]), .B0_t (key_s0_t[10]), .B0_f (key_s0_f[10]), .B1_t (key_s1_t[10]), .B1_f (key_s1_f[10]), .Z0_t (wk[10]), .Z0_f (new_AGEMA_signal_2488), .Z1_t (new_AGEMA_signal_2489), .Z1_f (new_AGEMA_signal_2490) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U10 ( .A0_t (key_s0_t[73]), .A0_f (key_s0_f[73]), .A1_t (key_s1_t[73]), .A1_f (key_s1_f[73]), .B0_t (key_s0_t[9]), .B0_f (key_s0_f[9]), .B1_t (key_s1_t[9]), .B1_f (key_s1_f[9]), .Z0_t (wk[9]), .Z0_f (new_AGEMA_signal_2497), .Z1_t (new_AGEMA_signal_2498), .Z1_f (new_AGEMA_signal_2499) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U9 ( .A0_t (key_s0_t[72]), .A0_f (key_s0_f[72]), .A1_t (key_s1_t[72]), .A1_f (key_s1_f[72]), .B0_t (key_s0_t[8]), .B0_f (key_s0_f[8]), .B1_t (key_s1_t[8]), .B1_f (key_s1_f[8]), .Z0_t (wk[8]), .Z0_f (new_AGEMA_signal_2506), .Z1_t (new_AGEMA_signal_2507), .Z1_f (new_AGEMA_signal_2508) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U8 ( .A0_t (key_s0_t[71]), .A0_f (key_s0_f[71]), .A1_t (key_s1_t[71]), .A1_f (key_s1_f[71]), .B0_t (key_s0_t[7]), .B0_f (key_s0_f[7]), .B1_t (key_s1_t[7]), .B1_f (key_s1_f[7]), .Z0_t (wk[7]), .Z0_f (new_AGEMA_signal_2515), .Z1_t (new_AGEMA_signal_2516), .Z1_f (new_AGEMA_signal_2517) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U7 ( .A0_t (key_s0_t[70]), .A0_f (key_s0_f[70]), .A1_t (key_s1_t[70]), .A1_f (key_s1_f[70]), .B0_t (key_s0_t[6]), .B0_f (key_s0_f[6]), .B1_t (key_s1_t[6]), .B1_f (key_s1_f[6]), .Z0_t (wk[6]), .Z0_f (new_AGEMA_signal_2524), .Z1_t (new_AGEMA_signal_2525), .Z1_f (new_AGEMA_signal_2526) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U6 ( .A0_t (key_s0_t[69]), .A0_f (key_s0_f[69]), .A1_t (key_s1_t[69]), .A1_f (key_s1_f[69]), .B0_t (key_s0_t[5]), .B0_f (key_s0_f[5]), .B1_t (key_s1_t[5]), .B1_f (key_s1_f[5]), .Z0_t (wk[5]), .Z0_f (new_AGEMA_signal_2533), .Z1_t (new_AGEMA_signal_2534), .Z1_f (new_AGEMA_signal_2535) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U5 ( .A0_t (key_s0_t[68]), .A0_f (key_s0_f[68]), .A1_t (key_s1_t[68]), .A1_f (key_s1_f[68]), .B0_t (key_s0_t[4]), .B0_f (key_s0_f[4]), .B1_t (key_s1_t[4]), .B1_f (key_s1_f[4]), .Z0_t (wk[4]), .Z0_f (new_AGEMA_signal_2542), .Z1_t (new_AGEMA_signal_2543), .Z1_f (new_AGEMA_signal_2544) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U4 ( .A0_t (key_s0_t[67]), .A0_f (key_s0_f[67]), .A1_t (key_s1_t[67]), .A1_f (key_s1_f[67]), .B0_t (key_s0_t[3]), .B0_f (key_s0_f[3]), .B1_t (key_s1_t[3]), .B1_f (key_s1_f[3]), .Z0_t (wk[3]), .Z0_f (new_AGEMA_signal_2551), .Z1_t (new_AGEMA_signal_2552), .Z1_f (new_AGEMA_signal_2553) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U3 ( .A0_t (key_s0_t[66]), .A0_f (key_s0_f[66]), .A1_t (key_s1_t[66]), .A1_f (key_s1_f[66]), .B0_t (key_s0_t[2]), .B0_f (key_s0_f[2]), .B1_t (key_s1_t[2]), .B1_f (key_s1_f[2]), .Z0_t (wk[2]), .Z0_f (new_AGEMA_signal_2560), .Z1_t (new_AGEMA_signal_2561), .Z1_f (new_AGEMA_signal_2562) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U2 ( .A0_t (key_s0_t[65]), .A0_f (key_s0_f[65]), .A1_t (key_s1_t[65]), .A1_f (key_s1_f[65]), .B0_t (key_s0_t[1]), .B0_f (key_s0_f[1]), .B1_t (key_s1_t[1]), .B1_f (key_s1_f[1]), .Z0_t (wk[1]), .Z0_f (new_AGEMA_signal_2569), .Z1_t (new_AGEMA_signal_2570), .Z1_f (new_AGEMA_signal_2571) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U1 ( .A0_t (key_s0_t[64]), .A0_f (key_s0_f[64]), .A1_t (key_s1_t[64]), .A1_f (key_s1_f[64]), .B0_t (key_s0_t[0]), .B0_f (key_s0_f[0]), .B1_t (key_s1_t[0]), .B1_f (key_s1_f[0]), .Z0_t (wk[0]), .Z0_f (new_AGEMA_signal_2578), .Z1_t (new_AGEMA_signal_2579), .Z1_f (new_AGEMA_signal_2580) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_U3 ( .A0_t (controller_n2), .A0_f (new_AGEMA_signal_2586), .B0_t (controller_n1), .B0_f (new_AGEMA_signal_2583), .Z0_t (done_t), .Z0_f (done_f) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) controller_U2 ( .A0_t (round_Signal[1]), .A0_f (new_AGEMA_signal_2581), .B0_t (round_Signal[0]), .B0_f (new_AGEMA_signal_2582), .Z0_t (controller_n1), .Z0_f (new_AGEMA_signal_2583) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) controller_U1 ( .A0_t (round_Signal[3]), .A0_f (new_AGEMA_signal_2584), .B0_t (round_Signal[2]), .B0_f (new_AGEMA_signal_2585), .Z0_t (controller_n2), .Z0_f (new_AGEMA_signal_2586) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U10 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (controller_roundCounter_n15), .B0_f (new_AGEMA_signal_3226), .Z0_t (controller_roundCounter_n5), .Z0_f (new_AGEMA_signal_4056) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U8 ( .A0_t (round_Signal[1]), .A0_f (new_AGEMA_signal_2581), .B0_t (controller_roundCounter_n6), .B0_f (new_AGEMA_signal_2588), .Z0_t (controller_roundCounter_n15), .Z0_f (new_AGEMA_signal_3226) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U7 ( .A0_t (reset_t), .A0_f (reset_f), .B0_t (round_Signal[0]), .B0_f (new_AGEMA_signal_2582), .Z0_t (controller_roundCounter_n6), .Z0_f (new_AGEMA_signal_2588) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U6 ( .A0_t (controller_roundCounter_n14), .A0_f (new_AGEMA_signal_3227), .B0_t (controller_roundCounter_n13), .B0_f (new_AGEMA_signal_2589), .Z0_t (controller_roundCounter_n4), .Z0_f (new_AGEMA_signal_4057) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U5 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (reset_t), .B0_f (reset_f), .Z0_t (controller_roundCounter_n13), .Z0_f (new_AGEMA_signal_2589) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U3 ( .A0_t (controller_roundCounter_N7), .A0_f (new_AGEMA_signal_2591), .B0_t (controller_roundCounter_n8), .B0_f (new_AGEMA_signal_2590), .Z0_t (controller_roundCounter_n14), .Z0_f (new_AGEMA_signal_3227) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U2 ( .A0_t (reset_t), .A0_f (reset_f), .B0_t (round_Signal[1]), .B0_f (new_AGEMA_signal_2581), .Z0_t (controller_roundCounter_n8), .Z0_f (new_AGEMA_signal_2590) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U1 ( .A0_t (reset_t), .A0_f (reset_f), .B0_t (round_Signal[0]), .B0_f (new_AGEMA_signal_2582), .Z0_t (controller_roundCounter_N7), .Z0_f (new_AGEMA_signal_2591) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) controller_roundCounter_U9_XOR1_U1 ( .A0_t (controller_roundCounter_n5), .A0_f (new_AGEMA_signal_4056), .B0_t (controller_roundCounter_n4), .B0_f (new_AGEMA_signal_4057), .Z0_t (controller_roundCounter_U9_X), .Z0_f (new_AGEMA_signal_4472) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U9_AND1_U1 ( .A0_t (round_Signal[3]), .A0_f (new_AGEMA_signal_2584), .B0_t (controller_roundCounter_U9_X), .B0_f (new_AGEMA_signal_4472), .Z0_t (controller_roundCounter_U9_Y), .Z0_f (new_AGEMA_signal_4778) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) controller_roundCounter_U9_XOR2_U1 ( .A0_t (controller_roundCounter_U9_Y), .A0_f (new_AGEMA_signal_4778), .B0_t (controller_roundCounter_n5), .B0_f (new_AGEMA_signal_4056), .Z0_t (round_Signal[3]), .Z0_f (new_AGEMA_signal_2584) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) controller_roundCounter_U11_XOR1_U1 ( .A0_t (controller_roundCounter_n6), .A0_f (new_AGEMA_signal_2588), .B0_t (controller_roundCounter_N7), .B0_f (new_AGEMA_signal_2591), .Z0_t (controller_roundCounter_U11_X), .Z0_f (new_AGEMA_signal_3228) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U11_AND1_U1 ( .A0_t (round_Signal[1]), .A0_f (new_AGEMA_signal_2581), .B0_t (controller_roundCounter_U11_X), .B0_f (new_AGEMA_signal_3228), .Z0_t (controller_roundCounter_U11_Y), .Z0_f (new_AGEMA_signal_4058) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) controller_roundCounter_U11_XOR2_U1 ( .A0_t (controller_roundCounter_U11_Y), .A0_f (new_AGEMA_signal_4058), .B0_t (controller_roundCounter_n6), .B0_f (new_AGEMA_signal_2588), .Z0_t (round_Signal[1]), .Z0_f (new_AGEMA_signal_2581) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) controller_roundCounter_U15_XOR1_U1 ( .A0_t (controller_roundCounter_n14), .A0_f (new_AGEMA_signal_3227), .B0_t (controller_roundCounter_n15), .B0_f (new_AGEMA_signal_3226), .Z0_t (controller_roundCounter_U15_X), .Z0_f (new_AGEMA_signal_4059) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U15_AND1_U1 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (controller_roundCounter_U15_X), .B0_f (new_AGEMA_signal_4059), .Z0_t (controller_roundCounter_U15_Y), .Z0_f (new_AGEMA_signal_4473) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) controller_roundCounter_U15_XOR2_U1 ( .A0_t (controller_roundCounter_U15_Y), .A0_f (new_AGEMA_signal_4473), .B0_t (controller_roundCounter_n14), .B0_f (new_AGEMA_signal_3227), .Z0_t (round_Signal[2]), .Z0_f (new_AGEMA_signal_2585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U128 ( .A0_t (wk[63]), .A0_f (new_AGEMA_signal_2011), .A1_t (new_AGEMA_signal_2012), .A1_f (new_AGEMA_signal_2013), .B0_t (DataIn_s0_t[63]), .B0_f (DataIn_s0_f[63]), .B1_t (DataIn_s1_t[63]), .B1_f (DataIn_s1_f[63]), .Z0_t (Midori_add_Result_Start[63]), .Z0_f (new_AGEMA_signal_3232), .Z1_t (new_AGEMA_signal_3233), .Z1_f (new_AGEMA_signal_3234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U127 ( .A0_t (wk[62]), .A0_f (new_AGEMA_signal_2020), .A1_t (new_AGEMA_signal_2021), .A1_f (new_AGEMA_signal_2022), .B0_t (DataIn_s0_t[62]), .B0_f (DataIn_s0_f[62]), .B1_t (DataIn_s1_t[62]), .B1_f (DataIn_s1_f[62]), .Z0_t (Midori_add_Result_Start[62]), .Z0_f (new_AGEMA_signal_3238), .Z1_t (new_AGEMA_signal_3239), .Z1_f (new_AGEMA_signal_3240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U126 ( .A0_t (wk[61]), .A0_f (new_AGEMA_signal_2029), .A1_t (new_AGEMA_signal_2030), .A1_f (new_AGEMA_signal_2031), .B0_t (DataIn_s0_t[61]), .B0_f (DataIn_s0_f[61]), .B1_t (DataIn_s1_t[61]), .B1_f (DataIn_s1_f[61]), .Z0_t (Midori_add_Result_Start[61]), .Z0_f (new_AGEMA_signal_3244), .Z1_t (new_AGEMA_signal_3245), .Z1_f (new_AGEMA_signal_3246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U125 ( .A0_t (wk[60]), .A0_f (new_AGEMA_signal_2038), .A1_t (new_AGEMA_signal_2039), .A1_f (new_AGEMA_signal_2040), .B0_t (DataIn_s0_t[60]), .B0_f (DataIn_s0_f[60]), .B1_t (DataIn_s1_t[60]), .B1_f (DataIn_s1_f[60]), .Z0_t (Midori_add_Result_Start[60]), .Z0_f (new_AGEMA_signal_3250), .Z1_t (new_AGEMA_signal_3251), .Z1_f (new_AGEMA_signal_3252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U124 ( .A0_t (wk[59]), .A0_f (new_AGEMA_signal_2047), .A1_t (new_AGEMA_signal_2048), .A1_f (new_AGEMA_signal_2049), .B0_t (DataIn_s0_t[59]), .B0_f (DataIn_s0_f[59]), .B1_t (DataIn_s1_t[59]), .B1_f (DataIn_s1_f[59]), .Z0_t (Midori_add_Result_Start[59]), .Z0_f (new_AGEMA_signal_3256), .Z1_t (new_AGEMA_signal_3257), .Z1_f (new_AGEMA_signal_3258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U123 ( .A0_t (wk[58]), .A0_f (new_AGEMA_signal_2056), .A1_t (new_AGEMA_signal_2057), .A1_f (new_AGEMA_signal_2058), .B0_t (DataIn_s0_t[58]), .B0_f (DataIn_s0_f[58]), .B1_t (DataIn_s1_t[58]), .B1_f (DataIn_s1_f[58]), .Z0_t (Midori_add_Result_Start[58]), .Z0_f (new_AGEMA_signal_3262), .Z1_t (new_AGEMA_signal_3263), .Z1_f (new_AGEMA_signal_3264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U122 ( .A0_t (wk[57]), .A0_f (new_AGEMA_signal_2065), .A1_t (new_AGEMA_signal_2066), .A1_f (new_AGEMA_signal_2067), .B0_t (DataIn_s0_t[57]), .B0_f (DataIn_s0_f[57]), .B1_t (DataIn_s1_t[57]), .B1_f (DataIn_s1_f[57]), .Z0_t (Midori_add_Result_Start[57]), .Z0_f (new_AGEMA_signal_3268), .Z1_t (new_AGEMA_signal_3269), .Z1_f (new_AGEMA_signal_3270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U121 ( .A0_t (wk[56]), .A0_f (new_AGEMA_signal_2074), .A1_t (new_AGEMA_signal_2075), .A1_f (new_AGEMA_signal_2076), .B0_t (DataIn_s0_t[56]), .B0_f (DataIn_s0_f[56]), .B1_t (DataIn_s1_t[56]), .B1_f (DataIn_s1_f[56]), .Z0_t (Midori_add_Result_Start[56]), .Z0_f (new_AGEMA_signal_3274), .Z1_t (new_AGEMA_signal_3275), .Z1_f (new_AGEMA_signal_3276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U120 ( .A0_t (wk[55]), .A0_f (new_AGEMA_signal_2083), .A1_t (new_AGEMA_signal_2084), .A1_f (new_AGEMA_signal_2085), .B0_t (DataIn_s0_t[55]), .B0_f (DataIn_s0_f[55]), .B1_t (DataIn_s1_t[55]), .B1_f (DataIn_s1_f[55]), .Z0_t (Midori_add_Result_Start[55]), .Z0_f (new_AGEMA_signal_3280), .Z1_t (new_AGEMA_signal_3281), .Z1_f (new_AGEMA_signal_3282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U119 ( .A0_t (wk[54]), .A0_f (new_AGEMA_signal_2092), .A1_t (new_AGEMA_signal_2093), .A1_f (new_AGEMA_signal_2094), .B0_t (DataIn_s0_t[54]), .B0_f (DataIn_s0_f[54]), .B1_t (DataIn_s1_t[54]), .B1_f (DataIn_s1_f[54]), .Z0_t (Midori_add_Result_Start[54]), .Z0_f (new_AGEMA_signal_3286), .Z1_t (new_AGEMA_signal_3287), .Z1_f (new_AGEMA_signal_3288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U118 ( .A0_t (wk[53]), .A0_f (new_AGEMA_signal_2101), .A1_t (new_AGEMA_signal_2102), .A1_f (new_AGEMA_signal_2103), .B0_t (DataIn_s0_t[53]), .B0_f (DataIn_s0_f[53]), .B1_t (DataIn_s1_t[53]), .B1_f (DataIn_s1_f[53]), .Z0_t (Midori_add_Result_Start[53]), .Z0_f (new_AGEMA_signal_3292), .Z1_t (new_AGEMA_signal_3293), .Z1_f (new_AGEMA_signal_3294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U117 ( .A0_t (wk[52]), .A0_f (new_AGEMA_signal_2110), .A1_t (new_AGEMA_signal_2111), .A1_f (new_AGEMA_signal_2112), .B0_t (DataIn_s0_t[52]), .B0_f (DataIn_s0_f[52]), .B1_t (DataIn_s1_t[52]), .B1_f (DataIn_s1_f[52]), .Z0_t (Midori_add_Result_Start[52]), .Z0_f (new_AGEMA_signal_3298), .Z1_t (new_AGEMA_signal_3299), .Z1_f (new_AGEMA_signal_3300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U116 ( .A0_t (wk[51]), .A0_f (new_AGEMA_signal_2119), .A1_t (new_AGEMA_signal_2120), .A1_f (new_AGEMA_signal_2121), .B0_t (DataIn_s0_t[51]), .B0_f (DataIn_s0_f[51]), .B1_t (DataIn_s1_t[51]), .B1_f (DataIn_s1_f[51]), .Z0_t (Midori_add_Result_Start[51]), .Z0_f (new_AGEMA_signal_3304), .Z1_t (new_AGEMA_signal_3305), .Z1_f (new_AGEMA_signal_3306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U115 ( .A0_t (wk[50]), .A0_f (new_AGEMA_signal_2128), .A1_t (new_AGEMA_signal_2129), .A1_f (new_AGEMA_signal_2130), .B0_t (DataIn_s0_t[50]), .B0_f (DataIn_s0_f[50]), .B1_t (DataIn_s1_t[50]), .B1_f (DataIn_s1_f[50]), .Z0_t (Midori_add_Result_Start[50]), .Z0_f (new_AGEMA_signal_3310), .Z1_t (new_AGEMA_signal_3311), .Z1_f (new_AGEMA_signal_3312) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U114 ( .A0_t (wk[49]), .A0_f (new_AGEMA_signal_2137), .A1_t (new_AGEMA_signal_2138), .A1_f (new_AGEMA_signal_2139), .B0_t (DataIn_s0_t[49]), .B0_f (DataIn_s0_f[49]), .B1_t (DataIn_s1_t[49]), .B1_f (DataIn_s1_f[49]), .Z0_t (Midori_add_Result_Start[49]), .Z0_f (new_AGEMA_signal_3316), .Z1_t (new_AGEMA_signal_3317), .Z1_f (new_AGEMA_signal_3318) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U113 ( .A0_t (wk[48]), .A0_f (new_AGEMA_signal_2146), .A1_t (new_AGEMA_signal_2147), .A1_f (new_AGEMA_signal_2148), .B0_t (DataIn_s0_t[48]), .B0_f (DataIn_s0_f[48]), .B1_t (DataIn_s1_t[48]), .B1_f (DataIn_s1_f[48]), .Z0_t (Midori_add_Result_Start[48]), .Z0_f (new_AGEMA_signal_3322), .Z1_t (new_AGEMA_signal_3323), .Z1_f (new_AGEMA_signal_3324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U112 ( .A0_t (wk[47]), .A0_f (new_AGEMA_signal_2155), .A1_t (new_AGEMA_signal_2156), .A1_f (new_AGEMA_signal_2157), .B0_t (DataIn_s0_t[47]), .B0_f (DataIn_s0_f[47]), .B1_t (DataIn_s1_t[47]), .B1_f (DataIn_s1_f[47]), .Z0_t (Midori_add_Result_Start[47]), .Z0_f (new_AGEMA_signal_3328), .Z1_t (new_AGEMA_signal_3329), .Z1_f (new_AGEMA_signal_3330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U111 ( .A0_t (wk[46]), .A0_f (new_AGEMA_signal_2164), .A1_t (new_AGEMA_signal_2165), .A1_f (new_AGEMA_signal_2166), .B0_t (DataIn_s0_t[46]), .B0_f (DataIn_s0_f[46]), .B1_t (DataIn_s1_t[46]), .B1_f (DataIn_s1_f[46]), .Z0_t (Midori_add_Result_Start[46]), .Z0_f (new_AGEMA_signal_3334), .Z1_t (new_AGEMA_signal_3335), .Z1_f (new_AGEMA_signal_3336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U110 ( .A0_t (wk[45]), .A0_f (new_AGEMA_signal_2173), .A1_t (new_AGEMA_signal_2174), .A1_f (new_AGEMA_signal_2175), .B0_t (DataIn_s0_t[45]), .B0_f (DataIn_s0_f[45]), .B1_t (DataIn_s1_t[45]), .B1_f (DataIn_s1_f[45]), .Z0_t (Midori_add_Result_Start[45]), .Z0_f (new_AGEMA_signal_3340), .Z1_t (new_AGEMA_signal_3341), .Z1_f (new_AGEMA_signal_3342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U109 ( .A0_t (wk[44]), .A0_f (new_AGEMA_signal_2182), .A1_t (new_AGEMA_signal_2183), .A1_f (new_AGEMA_signal_2184), .B0_t (DataIn_s0_t[44]), .B0_f (DataIn_s0_f[44]), .B1_t (DataIn_s1_t[44]), .B1_f (DataIn_s1_f[44]), .Z0_t (Midori_add_Result_Start[44]), .Z0_f (new_AGEMA_signal_3346), .Z1_t (new_AGEMA_signal_3347), .Z1_f (new_AGEMA_signal_3348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U108 ( .A0_t (wk[43]), .A0_f (new_AGEMA_signal_2191), .A1_t (new_AGEMA_signal_2192), .A1_f (new_AGEMA_signal_2193), .B0_t (DataIn_s0_t[43]), .B0_f (DataIn_s0_f[43]), .B1_t (DataIn_s1_t[43]), .B1_f (DataIn_s1_f[43]), .Z0_t (Midori_add_Result_Start[43]), .Z0_f (new_AGEMA_signal_3352), .Z1_t (new_AGEMA_signal_3353), .Z1_f (new_AGEMA_signal_3354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U107 ( .A0_t (wk[42]), .A0_f (new_AGEMA_signal_2200), .A1_t (new_AGEMA_signal_2201), .A1_f (new_AGEMA_signal_2202), .B0_t (DataIn_s0_t[42]), .B0_f (DataIn_s0_f[42]), .B1_t (DataIn_s1_t[42]), .B1_f (DataIn_s1_f[42]), .Z0_t (Midori_add_Result_Start[42]), .Z0_f (new_AGEMA_signal_3358), .Z1_t (new_AGEMA_signal_3359), .Z1_f (new_AGEMA_signal_3360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U106 ( .A0_t (wk[41]), .A0_f (new_AGEMA_signal_2209), .A1_t (new_AGEMA_signal_2210), .A1_f (new_AGEMA_signal_2211), .B0_t (DataIn_s0_t[41]), .B0_f (DataIn_s0_f[41]), .B1_t (DataIn_s1_t[41]), .B1_f (DataIn_s1_f[41]), .Z0_t (Midori_add_Result_Start[41]), .Z0_f (new_AGEMA_signal_3364), .Z1_t (new_AGEMA_signal_3365), .Z1_f (new_AGEMA_signal_3366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U105 ( .A0_t (wk[40]), .A0_f (new_AGEMA_signal_2218), .A1_t (new_AGEMA_signal_2219), .A1_f (new_AGEMA_signal_2220), .B0_t (DataIn_s0_t[40]), .B0_f (DataIn_s0_f[40]), .B1_t (DataIn_s1_t[40]), .B1_f (DataIn_s1_f[40]), .Z0_t (Midori_add_Result_Start[40]), .Z0_f (new_AGEMA_signal_3370), .Z1_t (new_AGEMA_signal_3371), .Z1_f (new_AGEMA_signal_3372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U104 ( .A0_t (wk[39]), .A0_f (new_AGEMA_signal_2227), .A1_t (new_AGEMA_signal_2228), .A1_f (new_AGEMA_signal_2229), .B0_t (DataIn_s0_t[39]), .B0_f (DataIn_s0_f[39]), .B1_t (DataIn_s1_t[39]), .B1_f (DataIn_s1_f[39]), .Z0_t (Midori_add_Result_Start[39]), .Z0_f (new_AGEMA_signal_3376), .Z1_t (new_AGEMA_signal_3377), .Z1_f (new_AGEMA_signal_3378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U103 ( .A0_t (wk[38]), .A0_f (new_AGEMA_signal_2236), .A1_t (new_AGEMA_signal_2237), .A1_f (new_AGEMA_signal_2238), .B0_t (DataIn_s0_t[38]), .B0_f (DataIn_s0_f[38]), .B1_t (DataIn_s1_t[38]), .B1_f (DataIn_s1_f[38]), .Z0_t (Midori_add_Result_Start[38]), .Z0_f (new_AGEMA_signal_3382), .Z1_t (new_AGEMA_signal_3383), .Z1_f (new_AGEMA_signal_3384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U102 ( .A0_t (wk[37]), .A0_f (new_AGEMA_signal_2245), .A1_t (new_AGEMA_signal_2246), .A1_f (new_AGEMA_signal_2247), .B0_t (DataIn_s0_t[37]), .B0_f (DataIn_s0_f[37]), .B1_t (DataIn_s1_t[37]), .B1_f (DataIn_s1_f[37]), .Z0_t (Midori_add_Result_Start[37]), .Z0_f (new_AGEMA_signal_3388), .Z1_t (new_AGEMA_signal_3389), .Z1_f (new_AGEMA_signal_3390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U101 ( .A0_t (wk[36]), .A0_f (new_AGEMA_signal_2254), .A1_t (new_AGEMA_signal_2255), .A1_f (new_AGEMA_signal_2256), .B0_t (DataIn_s0_t[36]), .B0_f (DataIn_s0_f[36]), .B1_t (DataIn_s1_t[36]), .B1_f (DataIn_s1_f[36]), .Z0_t (Midori_add_Result_Start[36]), .Z0_f (new_AGEMA_signal_3394), .Z1_t (new_AGEMA_signal_3395), .Z1_f (new_AGEMA_signal_3396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U100 ( .A0_t (wk[35]), .A0_f (new_AGEMA_signal_2263), .A1_t (new_AGEMA_signal_2264), .A1_f (new_AGEMA_signal_2265), .B0_t (DataIn_s0_t[35]), .B0_f (DataIn_s0_f[35]), .B1_t (DataIn_s1_t[35]), .B1_f (DataIn_s1_f[35]), .Z0_t (Midori_add_Result_Start[35]), .Z0_f (new_AGEMA_signal_3400), .Z1_t (new_AGEMA_signal_3401), .Z1_f (new_AGEMA_signal_3402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U99 ( .A0_t (wk[34]), .A0_f (new_AGEMA_signal_2272), .A1_t (new_AGEMA_signal_2273), .A1_f (new_AGEMA_signal_2274), .B0_t (DataIn_s0_t[34]), .B0_f (DataIn_s0_f[34]), .B1_t (DataIn_s1_t[34]), .B1_f (DataIn_s1_f[34]), .Z0_t (Midori_add_Result_Start[34]), .Z0_f (new_AGEMA_signal_3406), .Z1_t (new_AGEMA_signal_3407), .Z1_f (new_AGEMA_signal_3408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U98 ( .A0_t (wk[33]), .A0_f (new_AGEMA_signal_2281), .A1_t (new_AGEMA_signal_2282), .A1_f (new_AGEMA_signal_2283), .B0_t (DataIn_s0_t[33]), .B0_f (DataIn_s0_f[33]), .B1_t (DataIn_s1_t[33]), .B1_f (DataIn_s1_f[33]), .Z0_t (Midori_add_Result_Start[33]), .Z0_f (new_AGEMA_signal_3412), .Z1_t (new_AGEMA_signal_3413), .Z1_f (new_AGEMA_signal_3414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U97 ( .A0_t (wk[32]), .A0_f (new_AGEMA_signal_2290), .A1_t (new_AGEMA_signal_2291), .A1_f (new_AGEMA_signal_2292), .B0_t (DataIn_s0_t[32]), .B0_f (DataIn_s0_f[32]), .B1_t (DataIn_s1_t[32]), .B1_f (DataIn_s1_f[32]), .Z0_t (Midori_add_Result_Start[32]), .Z0_f (new_AGEMA_signal_3418), .Z1_t (new_AGEMA_signal_3419), .Z1_f (new_AGEMA_signal_3420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U96 ( .A0_t (wk[31]), .A0_f (new_AGEMA_signal_2299), .A1_t (new_AGEMA_signal_2300), .A1_f (new_AGEMA_signal_2301), .B0_t (DataIn_s0_t[31]), .B0_f (DataIn_s0_f[31]), .B1_t (DataIn_s1_t[31]), .B1_f (DataIn_s1_f[31]), .Z0_t (Midori_add_Result_Start[31]), .Z0_f (new_AGEMA_signal_3424), .Z1_t (new_AGEMA_signal_3425), .Z1_f (new_AGEMA_signal_3426) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U95 ( .A0_t (wk[30]), .A0_f (new_AGEMA_signal_2308), .A1_t (new_AGEMA_signal_2309), .A1_f (new_AGEMA_signal_2310), .B0_t (DataIn_s0_t[30]), .B0_f (DataIn_s0_f[30]), .B1_t (DataIn_s1_t[30]), .B1_f (DataIn_s1_f[30]), .Z0_t (Midori_add_Result_Start[30]), .Z0_f (new_AGEMA_signal_3430), .Z1_t (new_AGEMA_signal_3431), .Z1_f (new_AGEMA_signal_3432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U94 ( .A0_t (wk[29]), .A0_f (new_AGEMA_signal_2317), .A1_t (new_AGEMA_signal_2318), .A1_f (new_AGEMA_signal_2319), .B0_t (DataIn_s0_t[29]), .B0_f (DataIn_s0_f[29]), .B1_t (DataIn_s1_t[29]), .B1_f (DataIn_s1_f[29]), .Z0_t (Midori_add_Result_Start[29]), .Z0_f (new_AGEMA_signal_3436), .Z1_t (new_AGEMA_signal_3437), .Z1_f (new_AGEMA_signal_3438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U93 ( .A0_t (wk[28]), .A0_f (new_AGEMA_signal_2326), .A1_t (new_AGEMA_signal_2327), .A1_f (new_AGEMA_signal_2328), .B0_t (DataIn_s0_t[28]), .B0_f (DataIn_s0_f[28]), .B1_t (DataIn_s1_t[28]), .B1_f (DataIn_s1_f[28]), .Z0_t (Midori_add_Result_Start[28]), .Z0_f (new_AGEMA_signal_3442), .Z1_t (new_AGEMA_signal_3443), .Z1_f (new_AGEMA_signal_3444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U92 ( .A0_t (wk[27]), .A0_f (new_AGEMA_signal_2335), .A1_t (new_AGEMA_signal_2336), .A1_f (new_AGEMA_signal_2337), .B0_t (DataIn_s0_t[27]), .B0_f (DataIn_s0_f[27]), .B1_t (DataIn_s1_t[27]), .B1_f (DataIn_s1_f[27]), .Z0_t (Midori_add_Result_Start[27]), .Z0_f (new_AGEMA_signal_3448), .Z1_t (new_AGEMA_signal_3449), .Z1_f (new_AGEMA_signal_3450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U91 ( .A0_t (wk[26]), .A0_f (new_AGEMA_signal_2344), .A1_t (new_AGEMA_signal_2345), .A1_f (new_AGEMA_signal_2346), .B0_t (DataIn_s0_t[26]), .B0_f (DataIn_s0_f[26]), .B1_t (DataIn_s1_t[26]), .B1_f (DataIn_s1_f[26]), .Z0_t (Midori_add_Result_Start[26]), .Z0_f (new_AGEMA_signal_3454), .Z1_t (new_AGEMA_signal_3455), .Z1_f (new_AGEMA_signal_3456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U90 ( .A0_t (wk[25]), .A0_f (new_AGEMA_signal_2353), .A1_t (new_AGEMA_signal_2354), .A1_f (new_AGEMA_signal_2355), .B0_t (DataIn_s0_t[25]), .B0_f (DataIn_s0_f[25]), .B1_t (DataIn_s1_t[25]), .B1_f (DataIn_s1_f[25]), .Z0_t (Midori_add_Result_Start[25]), .Z0_f (new_AGEMA_signal_3460), .Z1_t (new_AGEMA_signal_3461), .Z1_f (new_AGEMA_signal_3462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U89 ( .A0_t (wk[24]), .A0_f (new_AGEMA_signal_2362), .A1_t (new_AGEMA_signal_2363), .A1_f (new_AGEMA_signal_2364), .B0_t (DataIn_s0_t[24]), .B0_f (DataIn_s0_f[24]), .B1_t (DataIn_s1_t[24]), .B1_f (DataIn_s1_f[24]), .Z0_t (Midori_add_Result_Start[24]), .Z0_f (new_AGEMA_signal_3466), .Z1_t (new_AGEMA_signal_3467), .Z1_f (new_AGEMA_signal_3468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U88 ( .A0_t (wk[23]), .A0_f (new_AGEMA_signal_2371), .A1_t (new_AGEMA_signal_2372), .A1_f (new_AGEMA_signal_2373), .B0_t (DataIn_s0_t[23]), .B0_f (DataIn_s0_f[23]), .B1_t (DataIn_s1_t[23]), .B1_f (DataIn_s1_f[23]), .Z0_t (Midori_add_Result_Start[23]), .Z0_f (new_AGEMA_signal_3472), .Z1_t (new_AGEMA_signal_3473), .Z1_f (new_AGEMA_signal_3474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U87 ( .A0_t (wk[22]), .A0_f (new_AGEMA_signal_2380), .A1_t (new_AGEMA_signal_2381), .A1_f (new_AGEMA_signal_2382), .B0_t (DataIn_s0_t[22]), .B0_f (DataIn_s0_f[22]), .B1_t (DataIn_s1_t[22]), .B1_f (DataIn_s1_f[22]), .Z0_t (Midori_add_Result_Start[22]), .Z0_f (new_AGEMA_signal_3478), .Z1_t (new_AGEMA_signal_3479), .Z1_f (new_AGEMA_signal_3480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U86 ( .A0_t (wk[21]), .A0_f (new_AGEMA_signal_2389), .A1_t (new_AGEMA_signal_2390), .A1_f (new_AGEMA_signal_2391), .B0_t (DataIn_s0_t[21]), .B0_f (DataIn_s0_f[21]), .B1_t (DataIn_s1_t[21]), .B1_f (DataIn_s1_f[21]), .Z0_t (Midori_add_Result_Start[21]), .Z0_f (new_AGEMA_signal_3484), .Z1_t (new_AGEMA_signal_3485), .Z1_f (new_AGEMA_signal_3486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U85 ( .A0_t (wk[20]), .A0_f (new_AGEMA_signal_2398), .A1_t (new_AGEMA_signal_2399), .A1_f (new_AGEMA_signal_2400), .B0_t (DataIn_s0_t[20]), .B0_f (DataIn_s0_f[20]), .B1_t (DataIn_s1_t[20]), .B1_f (DataIn_s1_f[20]), .Z0_t (Midori_add_Result_Start[20]), .Z0_f (new_AGEMA_signal_3490), .Z1_t (new_AGEMA_signal_3491), .Z1_f (new_AGEMA_signal_3492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U84 ( .A0_t (wk[19]), .A0_f (new_AGEMA_signal_2407), .A1_t (new_AGEMA_signal_2408), .A1_f (new_AGEMA_signal_2409), .B0_t (DataIn_s0_t[19]), .B0_f (DataIn_s0_f[19]), .B1_t (DataIn_s1_t[19]), .B1_f (DataIn_s1_f[19]), .Z0_t (Midori_add_Result_Start[19]), .Z0_f (new_AGEMA_signal_3496), .Z1_t (new_AGEMA_signal_3497), .Z1_f (new_AGEMA_signal_3498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U83 ( .A0_t (wk[18]), .A0_f (new_AGEMA_signal_2416), .A1_t (new_AGEMA_signal_2417), .A1_f (new_AGEMA_signal_2418), .B0_t (DataIn_s0_t[18]), .B0_f (DataIn_s0_f[18]), .B1_t (DataIn_s1_t[18]), .B1_f (DataIn_s1_f[18]), .Z0_t (Midori_add_Result_Start[18]), .Z0_f (new_AGEMA_signal_3502), .Z1_t (new_AGEMA_signal_3503), .Z1_f (new_AGEMA_signal_3504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U82 ( .A0_t (wk[17]), .A0_f (new_AGEMA_signal_2425), .A1_t (new_AGEMA_signal_2426), .A1_f (new_AGEMA_signal_2427), .B0_t (DataIn_s0_t[17]), .B0_f (DataIn_s0_f[17]), .B1_t (DataIn_s1_t[17]), .B1_f (DataIn_s1_f[17]), .Z0_t (Midori_add_Result_Start[17]), .Z0_f (new_AGEMA_signal_3508), .Z1_t (new_AGEMA_signal_3509), .Z1_f (new_AGEMA_signal_3510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U81 ( .A0_t (wk[16]), .A0_f (new_AGEMA_signal_2434), .A1_t (new_AGEMA_signal_2435), .A1_f (new_AGEMA_signal_2436), .B0_t (DataIn_s0_t[16]), .B0_f (DataIn_s0_f[16]), .B1_t (DataIn_s1_t[16]), .B1_f (DataIn_s1_f[16]), .Z0_t (Midori_add_Result_Start[16]), .Z0_f (new_AGEMA_signal_3514), .Z1_t (new_AGEMA_signal_3515), .Z1_f (new_AGEMA_signal_3516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U80 ( .A0_t (wk[15]), .A0_f (new_AGEMA_signal_2443), .A1_t (new_AGEMA_signal_2444), .A1_f (new_AGEMA_signal_2445), .B0_t (DataIn_s0_t[15]), .B0_f (DataIn_s0_f[15]), .B1_t (DataIn_s1_t[15]), .B1_f (DataIn_s1_f[15]), .Z0_t (Midori_add_Result_Start[15]), .Z0_f (new_AGEMA_signal_3520), .Z1_t (new_AGEMA_signal_3521), .Z1_f (new_AGEMA_signal_3522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U79 ( .A0_t (wk[14]), .A0_f (new_AGEMA_signal_2452), .A1_t (new_AGEMA_signal_2453), .A1_f (new_AGEMA_signal_2454), .B0_t (DataIn_s0_t[14]), .B0_f (DataIn_s0_f[14]), .B1_t (DataIn_s1_t[14]), .B1_f (DataIn_s1_f[14]), .Z0_t (Midori_add_Result_Start[14]), .Z0_f (new_AGEMA_signal_3526), .Z1_t (new_AGEMA_signal_3527), .Z1_f (new_AGEMA_signal_3528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U78 ( .A0_t (wk[13]), .A0_f (new_AGEMA_signal_2461), .A1_t (new_AGEMA_signal_2462), .A1_f (new_AGEMA_signal_2463), .B0_t (DataIn_s0_t[13]), .B0_f (DataIn_s0_f[13]), .B1_t (DataIn_s1_t[13]), .B1_f (DataIn_s1_f[13]), .Z0_t (Midori_add_Result_Start[13]), .Z0_f (new_AGEMA_signal_3532), .Z1_t (new_AGEMA_signal_3533), .Z1_f (new_AGEMA_signal_3534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U77 ( .A0_t (wk[12]), .A0_f (new_AGEMA_signal_2470), .A1_t (new_AGEMA_signal_2471), .A1_f (new_AGEMA_signal_2472), .B0_t (DataIn_s0_t[12]), .B0_f (DataIn_s0_f[12]), .B1_t (DataIn_s1_t[12]), .B1_f (DataIn_s1_f[12]), .Z0_t (Midori_add_Result_Start[12]), .Z0_f (new_AGEMA_signal_3538), .Z1_t (new_AGEMA_signal_3539), .Z1_f (new_AGEMA_signal_3540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U76 ( .A0_t (wk[11]), .A0_f (new_AGEMA_signal_2479), .A1_t (new_AGEMA_signal_2480), .A1_f (new_AGEMA_signal_2481), .B0_t (DataIn_s0_t[11]), .B0_f (DataIn_s0_f[11]), .B1_t (DataIn_s1_t[11]), .B1_f (DataIn_s1_f[11]), .Z0_t (Midori_add_Result_Start[11]), .Z0_f (new_AGEMA_signal_3544), .Z1_t (new_AGEMA_signal_3545), .Z1_f (new_AGEMA_signal_3546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U75 ( .A0_t (wk[10]), .A0_f (new_AGEMA_signal_2488), .A1_t (new_AGEMA_signal_2489), .A1_f (new_AGEMA_signal_2490), .B0_t (DataIn_s0_t[10]), .B0_f (DataIn_s0_f[10]), .B1_t (DataIn_s1_t[10]), .B1_f (DataIn_s1_f[10]), .Z0_t (Midori_add_Result_Start[10]), .Z0_f (new_AGEMA_signal_3550), .Z1_t (new_AGEMA_signal_3551), .Z1_f (new_AGEMA_signal_3552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U74 ( .A0_t (wk[9]), .A0_f (new_AGEMA_signal_2497), .A1_t (new_AGEMA_signal_2498), .A1_f (new_AGEMA_signal_2499), .B0_t (DataIn_s0_t[9]), .B0_f (DataIn_s0_f[9]), .B1_t (DataIn_s1_t[9]), .B1_f (DataIn_s1_f[9]), .Z0_t (Midori_add_Result_Start[9]), .Z0_f (new_AGEMA_signal_3556), .Z1_t (new_AGEMA_signal_3557), .Z1_f (new_AGEMA_signal_3558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U73 ( .A0_t (wk[8]), .A0_f (new_AGEMA_signal_2506), .A1_t (new_AGEMA_signal_2507), .A1_f (new_AGEMA_signal_2508), .B0_t (DataIn_s0_t[8]), .B0_f (DataIn_s0_f[8]), .B1_t (DataIn_s1_t[8]), .B1_f (DataIn_s1_f[8]), .Z0_t (Midori_add_Result_Start[8]), .Z0_f (new_AGEMA_signal_3562), .Z1_t (new_AGEMA_signal_3563), .Z1_f (new_AGEMA_signal_3564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U72 ( .A0_t (wk[7]), .A0_f (new_AGEMA_signal_2515), .A1_t (new_AGEMA_signal_2516), .A1_f (new_AGEMA_signal_2517), .B0_t (DataIn_s0_t[7]), .B0_f (DataIn_s0_f[7]), .B1_t (DataIn_s1_t[7]), .B1_f (DataIn_s1_f[7]), .Z0_t (Midori_add_Result_Start[7]), .Z0_f (new_AGEMA_signal_3568), .Z1_t (new_AGEMA_signal_3569), .Z1_f (new_AGEMA_signal_3570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U71 ( .A0_t (wk[6]), .A0_f (new_AGEMA_signal_2524), .A1_t (new_AGEMA_signal_2525), .A1_f (new_AGEMA_signal_2526), .B0_t (DataIn_s0_t[6]), .B0_f (DataIn_s0_f[6]), .B1_t (DataIn_s1_t[6]), .B1_f (DataIn_s1_f[6]), .Z0_t (Midori_add_Result_Start[6]), .Z0_f (new_AGEMA_signal_3574), .Z1_t (new_AGEMA_signal_3575), .Z1_f (new_AGEMA_signal_3576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U70 ( .A0_t (wk[5]), .A0_f (new_AGEMA_signal_2533), .A1_t (new_AGEMA_signal_2534), .A1_f (new_AGEMA_signal_2535), .B0_t (DataIn_s0_t[5]), .B0_f (DataIn_s0_f[5]), .B1_t (DataIn_s1_t[5]), .B1_f (DataIn_s1_f[5]), .Z0_t (Midori_add_Result_Start[5]), .Z0_f (new_AGEMA_signal_3580), .Z1_t (new_AGEMA_signal_3581), .Z1_f (new_AGEMA_signal_3582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U69 ( .A0_t (wk[4]), .A0_f (new_AGEMA_signal_2542), .A1_t (new_AGEMA_signal_2543), .A1_f (new_AGEMA_signal_2544), .B0_t (DataIn_s0_t[4]), .B0_f (DataIn_s0_f[4]), .B1_t (DataIn_s1_t[4]), .B1_f (DataIn_s1_f[4]), .Z0_t (Midori_add_Result_Start[4]), .Z0_f (new_AGEMA_signal_3586), .Z1_t (new_AGEMA_signal_3587), .Z1_f (new_AGEMA_signal_3588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U68 ( .A0_t (wk[3]), .A0_f (new_AGEMA_signal_2551), .A1_t (new_AGEMA_signal_2552), .A1_f (new_AGEMA_signal_2553), .B0_t (DataIn_s0_t[3]), .B0_f (DataIn_s0_f[3]), .B1_t (DataIn_s1_t[3]), .B1_f (DataIn_s1_f[3]), .Z0_t (Midori_add_Result_Start[3]), .Z0_f (new_AGEMA_signal_3592), .Z1_t (new_AGEMA_signal_3593), .Z1_f (new_AGEMA_signal_3594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U67 ( .A0_t (wk[2]), .A0_f (new_AGEMA_signal_2560), .A1_t (new_AGEMA_signal_2561), .A1_f (new_AGEMA_signal_2562), .B0_t (DataIn_s0_t[2]), .B0_f (DataIn_s0_f[2]), .B1_t (DataIn_s1_t[2]), .B1_f (DataIn_s1_f[2]), .Z0_t (Midori_add_Result_Start[2]), .Z0_f (new_AGEMA_signal_3598), .Z1_t (new_AGEMA_signal_3599), .Z1_f (new_AGEMA_signal_3600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U66 ( .A0_t (wk[1]), .A0_f (new_AGEMA_signal_2569), .A1_t (new_AGEMA_signal_2570), .A1_f (new_AGEMA_signal_2571), .B0_t (DataIn_s0_t[1]), .B0_f (DataIn_s0_f[1]), .B1_t (DataIn_s1_t[1]), .B1_f (DataIn_s1_f[1]), .Z0_t (Midori_add_Result_Start[1]), .Z0_f (new_AGEMA_signal_3604), .Z1_t (new_AGEMA_signal_3605), .Z1_f (new_AGEMA_signal_3606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U65 ( .A0_t (wk[0]), .A0_f (new_AGEMA_signal_2578), .A1_t (new_AGEMA_signal_2579), .A1_f (new_AGEMA_signal_2580), .B0_t (DataIn_s0_t[0]), .B0_f (DataIn_s0_f[0]), .B1_t (DataIn_s1_t[0]), .B1_f (DataIn_s1_f[0]), .Z0_t (Midori_add_Result_Start[0]), .Z0_f (new_AGEMA_signal_3610), .Z1_t (new_AGEMA_signal_3611), .Z1_f (new_AGEMA_signal_3612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U64 ( .A0_t (wk[56]), .A0_f (new_AGEMA_signal_2074), .A1_t (new_AGEMA_signal_2075), .A1_f (new_AGEMA_signal_2076), .B0_t (Midori_rounds_SR_Result[32]), .B0_f (new_AGEMA_signal_4769), .B1_t (new_AGEMA_signal_4770), .B1_f (new_AGEMA_signal_4771), .Z0_t (DataOut_s0_t[56]), .Z0_f (DataOut_s0_f[56]), .Z1_t (DataOut_s1_t[56]), .Z1_f (DataOut_s1_f[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U63 ( .A0_t (wk[52]), .A0_f (new_AGEMA_signal_2110), .A1_t (new_AGEMA_signal_2111), .A1_f (new_AGEMA_signal_2112), .B0_t (Midori_rounds_SR_Result[4]), .B0_f (new_AGEMA_signal_4763), .B1_t (new_AGEMA_signal_4764), .B1_f (new_AGEMA_signal_4765), .Z0_t (DataOut_s0_t[52]), .Z0_f (DataOut_s0_f[52]), .Z1_t (DataOut_s1_t[52]), .Z1_f (DataOut_s1_f[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U62 ( .A0_t (wk[36]), .A0_f (new_AGEMA_signal_2254), .A1_t (new_AGEMA_signal_2255), .A1_f (new_AGEMA_signal_2256), .B0_t (Midori_rounds_SR_Result[16]), .B0_f (new_AGEMA_signal_4739), .B1_t (new_AGEMA_signal_4740), .B1_f (new_AGEMA_signal_4741), .Z0_t (DataOut_s0_t[36]), .Z0_f (DataOut_s0_f[36]), .Z1_t (DataOut_s1_t[36]), .Z1_f (DataOut_s1_f[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U61 ( .A0_t (wk[32]), .A0_f (new_AGEMA_signal_2290), .A1_t (new_AGEMA_signal_2291), .A1_f (new_AGEMA_signal_2292), .B0_t (Midori_rounds_SR_Result[12]), .B0_f (new_AGEMA_signal_4733), .B1_t (new_AGEMA_signal_4734), .B1_f (new_AGEMA_signal_4735), .Z0_t (DataOut_s0_t[32]), .Z0_f (DataOut_s0_f[32]), .Z1_t (DataOut_s1_t[32]), .Z1_f (DataOut_s1_f[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U60 ( .A0_t (wk[28]), .A0_f (new_AGEMA_signal_2326), .A1_t (new_AGEMA_signal_2327), .A1_f (new_AGEMA_signal_2328), .B0_t (Midori_rounds_SR_Result[0]), .B0_f (new_AGEMA_signal_4727), .B1_t (new_AGEMA_signal_4728), .B1_f (new_AGEMA_signal_4729), .Z0_t (DataOut_s0_t[28]), .Z0_f (DataOut_s0_f[28]), .Z1_t (DataOut_s1_t[28]), .Z1_f (DataOut_s1_f[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U59 ( .A0_t (wk[0]), .A0_f (new_AGEMA_signal_2578), .A1_t (new_AGEMA_signal_2579), .A1_f (new_AGEMA_signal_2580), .B0_t (Midori_rounds_SR_Result[48]), .B0_f (new_AGEMA_signal_4685), .B1_t (new_AGEMA_signal_4686), .B1_f (new_AGEMA_signal_4687), .Z0_t (DataOut_s0_t[0]), .Z0_f (DataOut_s0_f[0]), .Z1_t (DataOut_s1_t[0]), .Z1_f (DataOut_s1_f[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U58 ( .A0_t (wk[59]), .A0_f (new_AGEMA_signal_2047), .A1_t (new_AGEMA_signal_2048), .A1_f (new_AGEMA_signal_2049), .B0_t (Midori_rounds_SR_Result[35]), .B0_f (new_AGEMA_signal_4448), .B1_t (new_AGEMA_signal_4449), .B1_f (new_AGEMA_signal_4450), .Z0_t (DataOut_s0_t[59]), .Z0_f (DataOut_s0_f[59]), .Z1_t (DataOut_s1_t[59]), .Z1_f (DataOut_s1_f[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U57 ( .A0_t (wk[55]), .A0_f (new_AGEMA_signal_2083), .A1_t (new_AGEMA_signal_2084), .A1_f (new_AGEMA_signal_2085), .B0_t (Midori_rounds_SR_Result[7]), .B0_f (new_AGEMA_signal_4436), .B1_t (new_AGEMA_signal_4437), .B1_f (new_AGEMA_signal_4438), .Z0_t (DataOut_s0_t[55]), .Z0_f (DataOut_s0_f[55]), .Z1_t (DataOut_s1_t[55]), .Z1_f (DataOut_s1_f[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U56 ( .A0_t (wk[39]), .A0_f (new_AGEMA_signal_2227), .A1_t (new_AGEMA_signal_2228), .A1_f (new_AGEMA_signal_2229), .B0_t (Midori_rounds_SR_Result[19]), .B0_f (new_AGEMA_signal_4388), .B1_t (new_AGEMA_signal_4389), .B1_f (new_AGEMA_signal_4390), .Z0_t (DataOut_s0_t[39]), .Z0_f (DataOut_s0_f[39]), .Z1_t (DataOut_s1_t[39]), .Z1_f (DataOut_s1_f[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U55 ( .A0_t (wk[35]), .A0_f (new_AGEMA_signal_2263), .A1_t (new_AGEMA_signal_2264), .A1_f (new_AGEMA_signal_2265), .B0_t (Midori_rounds_SR_Result[15]), .B0_f (new_AGEMA_signal_4376), .B1_t (new_AGEMA_signal_4377), .B1_f (new_AGEMA_signal_4378), .Z0_t (DataOut_s0_t[35]), .Z0_f (DataOut_s0_f[35]), .Z1_t (DataOut_s1_t[35]), .Z1_f (DataOut_s1_f[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U54 ( .A0_t (wk[31]), .A0_f (new_AGEMA_signal_2299), .A1_t (new_AGEMA_signal_2300), .A1_f (new_AGEMA_signal_2301), .B0_t (Midori_rounds_SR_Result[3]), .B0_f (new_AGEMA_signal_4364), .B1_t (new_AGEMA_signal_4365), .B1_f (new_AGEMA_signal_4366), .Z0_t (DataOut_s0_t[31]), .Z0_f (DataOut_s0_f[31]), .Z1_t (DataOut_s1_t[31]), .Z1_f (DataOut_s1_f[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U53 ( .A0_t (wk[3]), .A0_f (new_AGEMA_signal_2551), .A1_t (new_AGEMA_signal_2552), .A1_f (new_AGEMA_signal_2553), .B0_t (Midori_rounds_SR_Result[51]), .B0_f (new_AGEMA_signal_4280), .B1_t (new_AGEMA_signal_4281), .B1_f (new_AGEMA_signal_4282), .Z0_t (DataOut_s0_t[3]), .Z0_f (DataOut_s0_f[3]), .Z1_t (DataOut_s1_t[3]), .Z1_f (DataOut_s1_f[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U52 ( .A0_t (wk[63]), .A0_f (new_AGEMA_signal_2011), .A1_t (new_AGEMA_signal_2012), .A1_f (new_AGEMA_signal_2013), .B0_t (Midori_rounds_SR_Result[63]), .B0_f (new_AGEMA_signal_4466), .B1_t (new_AGEMA_signal_4467), .B1_f (new_AGEMA_signal_4468), .Z0_t (DataOut_s0_t[63]), .Z0_f (DataOut_s0_f[63]), .Z1_t (DataOut_s1_t[63]), .Z1_f (DataOut_s1_f[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U51 ( .A0_t (wk[62]), .A0_f (new_AGEMA_signal_2020), .A1_t (new_AGEMA_signal_2021), .A1_f (new_AGEMA_signal_2022), .B0_t (Midori_rounds_SR_Result[62]), .B0_f (new_AGEMA_signal_4775), .B1_t (new_AGEMA_signal_4776), .B1_f (new_AGEMA_signal_4777), .Z0_t (DataOut_s0_t[62]), .Z0_f (DataOut_s0_f[62]), .Z1_t (DataOut_s1_t[62]), .Z1_f (DataOut_s1_f[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U50 ( .A0_t (wk[61]), .A0_f (new_AGEMA_signal_2029), .A1_t (new_AGEMA_signal_2030), .A1_f (new_AGEMA_signal_2031), .B0_t (Midori_rounds_SR_Result[61]), .B0_f (new_AGEMA_signal_4469), .B1_t (new_AGEMA_signal_4470), .B1_f (new_AGEMA_signal_4471), .Z0_t (DataOut_s0_t[61]), .Z0_f (DataOut_s0_f[61]), .Z1_t (DataOut_s1_t[61]), .Z1_f (DataOut_s1_f[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U49 ( .A0_t (wk[58]), .A0_f (new_AGEMA_signal_2056), .A1_t (new_AGEMA_signal_2057), .A1_f (new_AGEMA_signal_2058), .B0_t (Midori_rounds_SR_Result[34]), .B0_f (new_AGEMA_signal_4766), .B1_t (new_AGEMA_signal_4767), .B1_f (new_AGEMA_signal_4768), .Z0_t (DataOut_s0_t[58]), .Z0_f (DataOut_s0_f[58]), .Z1_t (DataOut_s1_t[58]), .Z1_f (DataOut_s1_f[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U48 ( .A0_t (wk[57]), .A0_f (new_AGEMA_signal_2065), .A1_t (new_AGEMA_signal_2066), .A1_f (new_AGEMA_signal_2067), .B0_t (Midori_rounds_SR_Result[33]), .B0_f (new_AGEMA_signal_4451), .B1_t (new_AGEMA_signal_4452), .B1_f (new_AGEMA_signal_4453), .Z0_t (DataOut_s0_t[57]), .Z0_f (DataOut_s0_f[57]), .Z1_t (DataOut_s1_t[57]), .Z1_f (DataOut_s1_f[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U47 ( .A0_t (wk[54]), .A0_f (new_AGEMA_signal_2092), .A1_t (new_AGEMA_signal_2093), .A1_f (new_AGEMA_signal_2094), .B0_t (Midori_rounds_SR_Result[6]), .B0_f (new_AGEMA_signal_4760), .B1_t (new_AGEMA_signal_4761), .B1_f (new_AGEMA_signal_4762), .Z0_t (DataOut_s0_t[54]), .Z0_f (DataOut_s0_f[54]), .Z1_t (DataOut_s1_t[54]), .Z1_f (DataOut_s1_f[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U46 ( .A0_t (wk[53]), .A0_f (new_AGEMA_signal_2101), .A1_t (new_AGEMA_signal_2102), .A1_f (new_AGEMA_signal_2103), .B0_t (Midori_rounds_SR_Result[5]), .B0_f (new_AGEMA_signal_4439), .B1_t (new_AGEMA_signal_4440), .B1_f (new_AGEMA_signal_4441), .Z0_t (DataOut_s0_t[53]), .Z0_f (DataOut_s0_f[53]), .Z1_t (DataOut_s1_t[53]), .Z1_f (DataOut_s1_f[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U45 ( .A0_t (wk[51]), .A0_f (new_AGEMA_signal_2119), .A1_t (new_AGEMA_signal_2120), .A1_f (new_AGEMA_signal_2121), .B0_t (Midori_rounds_SR_Result[27]), .B0_f (new_AGEMA_signal_4430), .B1_t (new_AGEMA_signal_4431), .B1_f (new_AGEMA_signal_4432), .Z0_t (DataOut_s0_t[51]), .Z0_f (DataOut_s0_f[51]), .Z1_t (DataOut_s1_t[51]), .Z1_f (DataOut_s1_f[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U44 ( .A0_t (wk[50]), .A0_f (new_AGEMA_signal_2128), .A1_t (new_AGEMA_signal_2129), .A1_f (new_AGEMA_signal_2130), .B0_t (Midori_rounds_SR_Result[26]), .B0_f (new_AGEMA_signal_4757), .B1_t (new_AGEMA_signal_4758), .B1_f (new_AGEMA_signal_4759), .Z0_t (DataOut_s0_t[50]), .Z0_f (DataOut_s0_f[50]), .Z1_t (DataOut_s1_t[50]), .Z1_f (DataOut_s1_f[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U43 ( .A0_t (wk[49]), .A0_f (new_AGEMA_signal_2137), .A1_t (new_AGEMA_signal_2138), .A1_f (new_AGEMA_signal_2139), .B0_t (Midori_rounds_SR_Result[25]), .B0_f (new_AGEMA_signal_4433), .B1_t (new_AGEMA_signal_4434), .B1_f (new_AGEMA_signal_4435), .Z0_t (DataOut_s0_t[49]), .Z0_f (DataOut_s0_f[49]), .Z1_t (DataOut_s1_t[49]), .Z1_f (DataOut_s1_f[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U42 ( .A0_t (wk[47]), .A0_f (new_AGEMA_signal_2155), .A1_t (new_AGEMA_signal_2156), .A1_f (new_AGEMA_signal_2157), .B0_t (Midori_rounds_SR_Result[43]), .B0_f (new_AGEMA_signal_4418), .B1_t (new_AGEMA_signal_4419), .B1_f (new_AGEMA_signal_4420), .Z0_t (DataOut_s0_t[47]), .Z0_f (DataOut_s0_f[47]), .Z1_t (DataOut_s1_t[47]), .Z1_f (DataOut_s1_f[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U41 ( .A0_t (wk[46]), .A0_f (new_AGEMA_signal_2164), .A1_t (new_AGEMA_signal_2165), .A1_f (new_AGEMA_signal_2166), .B0_t (Midori_rounds_SR_Result[42]), .B0_f (new_AGEMA_signal_4751), .B1_t (new_AGEMA_signal_4752), .B1_f (new_AGEMA_signal_4753), .Z0_t (DataOut_s0_t[46]), .Z0_f (DataOut_s0_f[46]), .Z1_t (DataOut_s1_t[46]), .Z1_f (DataOut_s1_f[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U40 ( .A0_t (wk[45]), .A0_f (new_AGEMA_signal_2173), .A1_t (new_AGEMA_signal_2174), .A1_f (new_AGEMA_signal_2175), .B0_t (Midori_rounds_SR_Result[41]), .B0_f (new_AGEMA_signal_4421), .B1_t (new_AGEMA_signal_4422), .B1_f (new_AGEMA_signal_4423), .Z0_t (DataOut_s0_t[45]), .Z0_f (DataOut_s0_f[45]), .Z1_t (DataOut_s1_t[45]), .Z1_f (DataOut_s1_f[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U39 ( .A0_t (wk[43]), .A0_f (new_AGEMA_signal_2191), .A1_t (new_AGEMA_signal_2192), .A1_f (new_AGEMA_signal_2193), .B0_t (Midori_rounds_SR_Result[55]), .B0_f (new_AGEMA_signal_4406), .B1_t (new_AGEMA_signal_4407), .B1_f (new_AGEMA_signal_4408), .Z0_t (DataOut_s0_t[43]), .Z0_f (DataOut_s0_f[43]), .Z1_t (DataOut_s1_t[43]), .Z1_f (DataOut_s1_f[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U38 ( .A0_t (wk[41]), .A0_f (new_AGEMA_signal_2209), .A1_t (new_AGEMA_signal_2210), .A1_f (new_AGEMA_signal_2211), .B0_t (Midori_rounds_SR_Result[53]), .B0_f (new_AGEMA_signal_4409), .B1_t (new_AGEMA_signal_4410), .B1_f (new_AGEMA_signal_4411), .Z0_t (DataOut_s0_t[41]), .Z0_f (DataOut_s0_f[41]), .Z1_t (DataOut_s1_t[41]), .Z1_f (DataOut_s1_f[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U37 ( .A0_t (wk[38]), .A0_f (new_AGEMA_signal_2236), .A1_t (new_AGEMA_signal_2237), .A1_f (new_AGEMA_signal_2238), .B0_t (Midori_rounds_SR_Result[18]), .B0_f (new_AGEMA_signal_4736), .B1_t (new_AGEMA_signal_4737), .B1_f (new_AGEMA_signal_4738), .Z0_t (DataOut_s0_t[38]), .Z0_f (DataOut_s0_f[38]), .Z1_t (DataOut_s1_t[38]), .Z1_f (DataOut_s1_f[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U36 ( .A0_t (wk[6]), .A0_f (new_AGEMA_signal_2524), .A1_t (new_AGEMA_signal_2525), .A1_f (new_AGEMA_signal_2526), .B0_t (Midori_rounds_SR_Result[46]), .B0_f (new_AGEMA_signal_4691), .B1_t (new_AGEMA_signal_4692), .B1_f (new_AGEMA_signal_4693), .Z0_t (DataOut_s0_t[6]), .Z0_f (DataOut_s0_f[6]), .Z1_t (DataOut_s1_t[6]), .Z1_f (DataOut_s1_f[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U35 ( .A0_t (wk[5]), .A0_f (new_AGEMA_signal_2533), .A1_t (new_AGEMA_signal_2534), .A1_f (new_AGEMA_signal_2535), .B0_t (Midori_rounds_SR_Result[45]), .B0_f (new_AGEMA_signal_4301), .B1_t (new_AGEMA_signal_4302), .B1_f (new_AGEMA_signal_4303), .Z0_t (DataOut_s0_t[5]), .Z0_f (DataOut_s0_f[5]), .Z1_t (DataOut_s1_t[5]), .Z1_f (DataOut_s1_f[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U34 ( .A0_t (wk[2]), .A0_f (new_AGEMA_signal_2560), .A1_t (new_AGEMA_signal_2561), .A1_f (new_AGEMA_signal_2562), .B0_t (Midori_rounds_SR_Result[50]), .B0_f (new_AGEMA_signal_4682), .B1_t (new_AGEMA_signal_4683), .B1_f (new_AGEMA_signal_4684), .Z0_t (DataOut_s0_t[2]), .Z0_f (DataOut_s0_f[2]), .Z1_t (DataOut_s1_t[2]), .Z1_f (DataOut_s1_f[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U33 ( .A0_t (wk[1]), .A0_f (new_AGEMA_signal_2569), .A1_t (new_AGEMA_signal_2570), .A1_f (new_AGEMA_signal_2571), .B0_t (Midori_rounds_SR_Result[49]), .B0_f (new_AGEMA_signal_4283), .B1_t (new_AGEMA_signal_4284), .B1_f (new_AGEMA_signal_4285), .Z0_t (DataOut_s0_t[1]), .Z0_f (DataOut_s0_f[1]), .Z1_t (DataOut_s1_t[1]), .Z1_f (DataOut_s1_f[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U32 ( .A0_t (wk[60]), .A0_f (new_AGEMA_signal_2038), .A1_t (new_AGEMA_signal_2039), .A1_f (new_AGEMA_signal_2040), .B0_t (Midori_rounds_SR_Result[60]), .B0_f (new_AGEMA_signal_4772), .B1_t (new_AGEMA_signal_4773), .B1_f (new_AGEMA_signal_4774), .Z0_t (DataOut_s0_t[60]), .Z0_f (DataOut_s0_f[60]), .Z1_t (DataOut_s1_t[60]), .Z1_f (DataOut_s1_f[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U31 ( .A0_t (wk[48]), .A0_f (new_AGEMA_signal_2146), .A1_t (new_AGEMA_signal_2147), .A1_f (new_AGEMA_signal_2148), .B0_t (Midori_rounds_SR_Result[24]), .B0_f (new_AGEMA_signal_4754), .B1_t (new_AGEMA_signal_4755), .B1_f (new_AGEMA_signal_4756), .Z0_t (DataOut_s0_t[48]), .Z0_f (DataOut_s0_f[48]), .Z1_t (DataOut_s1_t[48]), .Z1_f (DataOut_s1_f[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U30 ( .A0_t (wk[44]), .A0_f (new_AGEMA_signal_2182), .A1_t (new_AGEMA_signal_2183), .A1_f (new_AGEMA_signal_2184), .B0_t (Midori_rounds_SR_Result[40]), .B0_f (new_AGEMA_signal_4748), .B1_t (new_AGEMA_signal_4749), .B1_f (new_AGEMA_signal_4750), .Z0_t (DataOut_s0_t[44]), .Z0_f (DataOut_s0_f[44]), .Z1_t (DataOut_s1_t[44]), .Z1_f (DataOut_s1_f[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U29 ( .A0_t (wk[42]), .A0_f (new_AGEMA_signal_2200), .A1_t (new_AGEMA_signal_2201), .A1_f (new_AGEMA_signal_2202), .B0_t (Midori_rounds_SR_Result[54]), .B0_f (new_AGEMA_signal_4745), .B1_t (new_AGEMA_signal_4746), .B1_f (new_AGEMA_signal_4747), .Z0_t (DataOut_s0_t[42]), .Z0_f (DataOut_s0_f[42]), .Z1_t (DataOut_s1_t[42]), .Z1_f (DataOut_s1_f[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U28 ( .A0_t (wk[37]), .A0_f (new_AGEMA_signal_2245), .A1_t (new_AGEMA_signal_2246), .A1_f (new_AGEMA_signal_2247), .B0_t (Midori_rounds_SR_Result[17]), .B0_f (new_AGEMA_signal_4391), .B1_t (new_AGEMA_signal_4392), .B1_f (new_AGEMA_signal_4393), .Z0_t (DataOut_s0_t[37]), .Z0_f (DataOut_s0_f[37]), .Z1_t (DataOut_s1_t[37]), .Z1_f (DataOut_s1_f[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U27 ( .A0_t (wk[34]), .A0_f (new_AGEMA_signal_2272), .A1_t (new_AGEMA_signal_2273), .A1_f (new_AGEMA_signal_2274), .B0_t (Midori_rounds_SR_Result[14]), .B0_f (new_AGEMA_signal_4730), .B1_t (new_AGEMA_signal_4731), .B1_f (new_AGEMA_signal_4732), .Z0_t (DataOut_s0_t[34]), .Z0_f (DataOut_s0_f[34]), .Z1_t (DataOut_s1_t[34]), .Z1_f (DataOut_s1_f[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U26 ( .A0_t (wk[33]), .A0_f (new_AGEMA_signal_2281), .A1_t (new_AGEMA_signal_2282), .A1_f (new_AGEMA_signal_2283), .B0_t (Midori_rounds_SR_Result[13]), .B0_f (new_AGEMA_signal_4379), .B1_t (new_AGEMA_signal_4380), .B1_f (new_AGEMA_signal_4381), .Z0_t (DataOut_s0_t[33]), .Z0_f (DataOut_s0_f[33]), .Z1_t (DataOut_s1_t[33]), .Z1_f (DataOut_s1_f[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U25 ( .A0_t (wk[30]), .A0_f (new_AGEMA_signal_2308), .A1_t (new_AGEMA_signal_2309), .A1_f (new_AGEMA_signal_2310), .B0_t (Midori_rounds_SR_Result[2]), .B0_f (new_AGEMA_signal_4724), .B1_t (new_AGEMA_signal_4725), .B1_f (new_AGEMA_signal_4726), .Z0_t (DataOut_s0_t[30]), .Z0_f (DataOut_s0_f[30]), .Z1_t (DataOut_s1_t[30]), .Z1_f (DataOut_s1_f[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U24 ( .A0_t (wk[29]), .A0_f (new_AGEMA_signal_2317), .A1_t (new_AGEMA_signal_2318), .A1_f (new_AGEMA_signal_2319), .B0_t (Midori_rounds_SR_Result[1]), .B0_f (new_AGEMA_signal_4367), .B1_t (new_AGEMA_signal_4368), .B1_f (new_AGEMA_signal_4369), .Z0_t (DataOut_s0_t[29]), .Z0_f (DataOut_s0_f[29]), .Z1_t (DataOut_s1_t[29]), .Z1_f (DataOut_s1_f[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U23 ( .A0_t (wk[27]), .A0_f (new_AGEMA_signal_2335), .A1_t (new_AGEMA_signal_2336), .A1_f (new_AGEMA_signal_2337), .B0_t (Midori_rounds_SR_Result[31]), .B0_f (new_AGEMA_signal_4358), .B1_t (new_AGEMA_signal_4359), .B1_f (new_AGEMA_signal_4360), .Z0_t (DataOut_s0_t[27]), .Z0_f (DataOut_s0_f[27]), .Z1_t (DataOut_s1_t[27]), .Z1_f (DataOut_s1_f[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U22 ( .A0_t (wk[26]), .A0_f (new_AGEMA_signal_2344), .A1_t (new_AGEMA_signal_2345), .A1_f (new_AGEMA_signal_2346), .B0_t (Midori_rounds_SR_Result[30]), .B0_f (new_AGEMA_signal_4721), .B1_t (new_AGEMA_signal_4722), .B1_f (new_AGEMA_signal_4723), .Z0_t (DataOut_s0_t[26]), .Z0_f (DataOut_s0_f[26]), .Z1_t (DataOut_s1_t[26]), .Z1_f (DataOut_s1_f[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U21 ( .A0_t (wk[25]), .A0_f (new_AGEMA_signal_2353), .A1_t (new_AGEMA_signal_2354), .A1_f (new_AGEMA_signal_2355), .B0_t (Midori_rounds_SR_Result[29]), .B0_f (new_AGEMA_signal_4361), .B1_t (new_AGEMA_signal_4362), .B1_f (new_AGEMA_signal_4363), .Z0_t (DataOut_s0_t[25]), .Z0_f (DataOut_s0_f[25]), .Z1_t (DataOut_s1_t[25]), .Z1_f (DataOut_s1_f[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U20 ( .A0_t (wk[23]), .A0_f (new_AGEMA_signal_2371), .A1_t (new_AGEMA_signal_2372), .A1_f (new_AGEMA_signal_2373), .B0_t (Midori_rounds_SR_Result[59]), .B0_f (new_AGEMA_signal_4346), .B1_t (new_AGEMA_signal_4347), .B1_f (new_AGEMA_signal_4348), .Z0_t (DataOut_s0_t[23]), .Z0_f (DataOut_s0_f[23]), .Z1_t (DataOut_s1_t[23]), .Z1_f (DataOut_s1_f[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U19 ( .A0_t (wk[22]), .A0_f (new_AGEMA_signal_2380), .A1_t (new_AGEMA_signal_2381), .A1_f (new_AGEMA_signal_2382), .B0_t (Midori_rounds_SR_Result[58]), .B0_f (new_AGEMA_signal_4715), .B1_t (new_AGEMA_signal_4716), .B1_f (new_AGEMA_signal_4717), .Z0_t (DataOut_s0_t[22]), .Z0_f (DataOut_s0_f[22]), .Z1_t (DataOut_s1_t[22]), .Z1_f (DataOut_s1_f[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U18 ( .A0_t (wk[21]), .A0_f (new_AGEMA_signal_2389), .A1_t (new_AGEMA_signal_2390), .A1_f (new_AGEMA_signal_2391), .B0_t (Midori_rounds_SR_Result[57]), .B0_f (new_AGEMA_signal_4349), .B1_t (new_AGEMA_signal_4350), .B1_f (new_AGEMA_signal_4351), .Z0_t (DataOut_s0_t[21]), .Z0_f (DataOut_s0_f[21]), .Z1_t (DataOut_s1_t[21]), .Z1_f (DataOut_s1_f[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U17 ( .A0_t (wk[19]), .A0_f (new_AGEMA_signal_2407), .A1_t (new_AGEMA_signal_2408), .A1_f (new_AGEMA_signal_2409), .B0_t (Midori_rounds_SR_Result[39]), .B0_f (new_AGEMA_signal_4334), .B1_t (new_AGEMA_signal_4335), .B1_f (new_AGEMA_signal_4336), .Z0_t (DataOut_s0_t[19]), .Z0_f (DataOut_s0_f[19]), .Z1_t (DataOut_s1_t[19]), .Z1_f (DataOut_s1_f[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U16 ( .A0_t (wk[18]), .A0_f (new_AGEMA_signal_2416), .A1_t (new_AGEMA_signal_2417), .A1_f (new_AGEMA_signal_2418), .B0_t (Midori_rounds_SR_Result[38]), .B0_f (new_AGEMA_signal_4709), .B1_t (new_AGEMA_signal_4710), .B1_f (new_AGEMA_signal_4711), .Z0_t (DataOut_s0_t[18]), .Z0_f (DataOut_s0_f[18]), .Z1_t (DataOut_s1_t[18]), .Z1_f (DataOut_s1_f[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U15 ( .A0_t (wk[17]), .A0_f (new_AGEMA_signal_2425), .A1_t (new_AGEMA_signal_2426), .A1_f (new_AGEMA_signal_2427), .B0_t (Midori_rounds_SR_Result[37]), .B0_f (new_AGEMA_signal_4337), .B1_t (new_AGEMA_signal_4338), .B1_f (new_AGEMA_signal_4339), .Z0_t (DataOut_s0_t[17]), .Z0_f (DataOut_s0_f[17]), .Z1_t (DataOut_s1_t[17]), .Z1_f (DataOut_s1_f[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U14 ( .A0_t (wk[15]), .A0_f (new_AGEMA_signal_2443), .A1_t (new_AGEMA_signal_2444), .A1_f (new_AGEMA_signal_2445), .B0_t (Midori_rounds_SR_Result[23]), .B0_f (new_AGEMA_signal_4322), .B1_t (new_AGEMA_signal_4323), .B1_f (new_AGEMA_signal_4324), .Z0_t (DataOut_s0_t[15]), .Z0_f (DataOut_s0_f[15]), .Z1_t (DataOut_s1_t[15]), .Z1_f (DataOut_s1_f[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U13 ( .A0_t (wk[14]), .A0_f (new_AGEMA_signal_2452), .A1_t (new_AGEMA_signal_2453), .A1_f (new_AGEMA_signal_2454), .B0_t (Midori_rounds_SR_Result[22]), .B0_f (new_AGEMA_signal_4703), .B1_t (new_AGEMA_signal_4704), .B1_f (new_AGEMA_signal_4705), .Z0_t (DataOut_s0_t[14]), .Z0_f (DataOut_s0_f[14]), .Z1_t (DataOut_s1_t[14]), .Z1_f (DataOut_s1_f[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U12 ( .A0_t (wk[13]), .A0_f (new_AGEMA_signal_2461), .A1_t (new_AGEMA_signal_2462), .A1_f (new_AGEMA_signal_2463), .B0_t (Midori_rounds_SR_Result[21]), .B0_f (new_AGEMA_signal_4325), .B1_t (new_AGEMA_signal_4326), .B1_f (new_AGEMA_signal_4327), .Z0_t (DataOut_s0_t[13]), .Z0_f (DataOut_s0_f[13]), .Z1_t (DataOut_s1_t[13]), .Z1_f (DataOut_s1_f[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U11 ( .A0_t (wk[11]), .A0_f (new_AGEMA_signal_2479), .A1_t (new_AGEMA_signal_2480), .A1_f (new_AGEMA_signal_2481), .B0_t (Midori_rounds_SR_Result[11]), .B0_f (new_AGEMA_signal_4310), .B1_t (new_AGEMA_signal_4311), .B1_f (new_AGEMA_signal_4312), .Z0_t (DataOut_s0_t[11]), .Z0_f (DataOut_s0_f[11]), .Z1_t (DataOut_s1_t[11]), .Z1_f (DataOut_s1_f[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U10 ( .A0_t (wk[10]), .A0_f (new_AGEMA_signal_2488), .A1_t (new_AGEMA_signal_2489), .A1_f (new_AGEMA_signal_2490), .B0_t (Midori_rounds_SR_Result[10]), .B0_f (new_AGEMA_signal_4697), .B1_t (new_AGEMA_signal_4698), .B1_f (new_AGEMA_signal_4699), .Z0_t (DataOut_s0_t[10]), .Z0_f (DataOut_s0_f[10]), .Z1_t (DataOut_s1_t[10]), .Z1_f (DataOut_s1_f[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U9 ( .A0_t (wk[9]), .A0_f (new_AGEMA_signal_2497), .A1_t (new_AGEMA_signal_2498), .A1_f (new_AGEMA_signal_2499), .B0_t (Midori_rounds_SR_Result[9]), .B0_f (new_AGEMA_signal_4313), .B1_t (new_AGEMA_signal_4314), .B1_f (new_AGEMA_signal_4315), .Z0_t (DataOut_s0_t[9]), .Z0_f (DataOut_s0_f[9]), .Z1_t (DataOut_s1_t[9]), .Z1_f (DataOut_s1_f[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U8 ( .A0_t (wk[7]), .A0_f (new_AGEMA_signal_2515), .A1_t (new_AGEMA_signal_2516), .A1_f (new_AGEMA_signal_2517), .B0_t (Midori_rounds_SR_Result[47]), .B0_f (new_AGEMA_signal_4298), .B1_t (new_AGEMA_signal_4299), .B1_f (new_AGEMA_signal_4300), .Z0_t (DataOut_s0_t[7]), .Z0_f (DataOut_s0_f[7]), .Z1_t (DataOut_s1_t[7]), .Z1_f (DataOut_s1_f[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U7 ( .A0_t (wk[40]), .A0_f (new_AGEMA_signal_2218), .A1_t (new_AGEMA_signal_2219), .A1_f (new_AGEMA_signal_2220), .B0_t (Midori_rounds_SR_Result[52]), .B0_f (new_AGEMA_signal_4742), .B1_t (new_AGEMA_signal_4743), .B1_f (new_AGEMA_signal_4744), .Z0_t (DataOut_s0_t[40]), .Z0_f (DataOut_s0_f[40]), .Z1_t (DataOut_s1_t[40]), .Z1_f (DataOut_s1_f[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U6 ( .A0_t (wk[24]), .A0_f (new_AGEMA_signal_2362), .A1_t (new_AGEMA_signal_2363), .A1_f (new_AGEMA_signal_2364), .B0_t (Midori_rounds_SR_Result[28]), .B0_f (new_AGEMA_signal_4718), .B1_t (new_AGEMA_signal_4719), .B1_f (new_AGEMA_signal_4720), .Z0_t (DataOut_s0_t[24]), .Z0_f (DataOut_s0_f[24]), .Z1_t (DataOut_s1_t[24]), .Z1_f (DataOut_s1_f[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U5 ( .A0_t (wk[20]), .A0_f (new_AGEMA_signal_2398), .A1_t (new_AGEMA_signal_2399), .A1_f (new_AGEMA_signal_2400), .B0_t (Midori_rounds_SR_Result[56]), .B0_f (new_AGEMA_signal_4712), .B1_t (new_AGEMA_signal_4713), .B1_f (new_AGEMA_signal_4714), .Z0_t (DataOut_s0_t[20]), .Z0_f (DataOut_s0_f[20]), .Z1_t (DataOut_s1_t[20]), .Z1_f (DataOut_s1_f[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U4 ( .A0_t (wk[16]), .A0_f (new_AGEMA_signal_2434), .A1_t (new_AGEMA_signal_2435), .A1_f (new_AGEMA_signal_2436), .B0_t (Midori_rounds_SR_Result[36]), .B0_f (new_AGEMA_signal_4706), .B1_t (new_AGEMA_signal_4707), .B1_f (new_AGEMA_signal_4708), .Z0_t (DataOut_s0_t[16]), .Z0_f (DataOut_s0_f[16]), .Z1_t (DataOut_s1_t[16]), .Z1_f (DataOut_s1_f[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U3 ( .A0_t (wk[12]), .A0_f (new_AGEMA_signal_2470), .A1_t (new_AGEMA_signal_2471), .A1_f (new_AGEMA_signal_2472), .B0_t (Midori_rounds_SR_Result[20]), .B0_f (new_AGEMA_signal_4700), .B1_t (new_AGEMA_signal_4701), .B1_f (new_AGEMA_signal_4702), .Z0_t (DataOut_s0_t[12]), .Z0_f (DataOut_s0_f[12]), .Z1_t (DataOut_s1_t[12]), .Z1_f (DataOut_s1_f[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U2 ( .A0_t (wk[8]), .A0_f (new_AGEMA_signal_2506), .A1_t (new_AGEMA_signal_2507), .A1_f (new_AGEMA_signal_2508), .B0_t (Midori_rounds_SR_Result[8]), .B0_f (new_AGEMA_signal_4694), .B1_t (new_AGEMA_signal_4695), .B1_f (new_AGEMA_signal_4696), .Z0_t (DataOut_s0_t[8]), .Z0_f (DataOut_s0_f[8]), .Z1_t (DataOut_s1_t[8]), .Z1_f (DataOut_s1_f[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U1 ( .A0_t (wk[4]), .A0_f (new_AGEMA_signal_2542), .A1_t (new_AGEMA_signal_2543), .A1_f (new_AGEMA_signal_2544), .B0_t (Midori_rounds_SR_Result[44]), .B0_f (new_AGEMA_signal_4688), .B1_t (new_AGEMA_signal_4689), .B1_f (new_AGEMA_signal_4690), .Z0_t (DataOut_s0_t[4]), .Z0_f (DataOut_s0_f[4]), .Z1_t (DataOut_s1_t[4]), .Z1_f (DataOut_s1_f[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U144 ( .A0_t (Midori_rounds_SR_Result[60]), .A0_f (new_AGEMA_signal_4772), .A1_t (new_AGEMA_signal_4773), .A1_f (new_AGEMA_signal_4774), .B0_t (Midori_rounds_n16), .B0_f (new_AGEMA_signal_5458), .B1_t (new_AGEMA_signal_5459), .B1_f (new_AGEMA_signal_5460), .Z0_t (Midori_rounds_sub_ResultXORkey[60]), .Z0_f (new_AGEMA_signal_5604), .Z1_t (new_AGEMA_signal_5605), .Z1_f (new_AGEMA_signal_5606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U143 ( .A0_t (Midori_rounds_SR_Inv_Result[60]), .A0_f (new_AGEMA_signal_6797), .A1_t (new_AGEMA_signal_6798), .A1_f (new_AGEMA_signal_6799), .B0_t (Midori_rounds_n16), .B0_f (new_AGEMA_signal_5458), .B1_t (new_AGEMA_signal_5459), .B1_f (new_AGEMA_signal_5460), .Z0_t (Midori_rounds_mul_ResultXORkey[60]), .Z0_f (new_AGEMA_signal_6821), .Z1_t (new_AGEMA_signal_6822), .Z1_f (new_AGEMA_signal_6823) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U142 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[15]), .A1_f (new_AGEMA_signal_5353), .B0_t (Midori_rounds_SelectedKey[60]), .B0_f (new_AGEMA_signal_4268), .B1_t (new_AGEMA_signal_4269), .B1_f (new_AGEMA_signal_4270), .Z0_t (Midori_rounds_n16), .Z0_f (new_AGEMA_signal_5458), .Z1_t (new_AGEMA_signal_5459), .Z1_f (new_AGEMA_signal_5460) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U141 ( .A0_t (Midori_rounds_SR_Result[44]), .A0_f (new_AGEMA_signal_4688), .A1_t (new_AGEMA_signal_4689), .A1_f (new_AGEMA_signal_4690), .B0_t (Midori_rounds_n15), .B0_f (new_AGEMA_signal_5978), .B1_t (new_AGEMA_signal_5979), .B1_f (new_AGEMA_signal_5980), .Z0_t (Midori_rounds_sub_ResultXORkey[4]), .Z0_f (new_AGEMA_signal_6167), .Z1_t (new_AGEMA_signal_6168), .Z1_f (new_AGEMA_signal_6169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U140 ( .A0_t (Midori_rounds_SR_Inv_Result[52]), .A0_f (new_AGEMA_signal_6779), .A1_t (new_AGEMA_signal_6780), .A1_f (new_AGEMA_signal_6781), .B0_t (Midori_rounds_n15), .B0_f (new_AGEMA_signal_5978), .B1_t (new_AGEMA_signal_5979), .B1_f (new_AGEMA_signal_5980), .Z0_t (Midori_rounds_mul_ResultXORkey[4]), .Z0_f (new_AGEMA_signal_6782), .Z1_t (new_AGEMA_signal_6783), .Z1_f (new_AGEMA_signal_6784) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U139 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[1]), .A1_f (new_AGEMA_signal_5863), .B0_t (Midori_rounds_SelectedKey[4]), .B0_f (new_AGEMA_signal_4100), .B1_t (new_AGEMA_signal_4101), .B1_f (new_AGEMA_signal_4102), .Z0_t (Midori_rounds_n15), .Z0_f (new_AGEMA_signal_5978), .Z1_t (new_AGEMA_signal_5979), .Z1_f (new_AGEMA_signal_5980) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U138 ( .A0_t (Midori_rounds_SR_Result[32]), .A0_f (new_AGEMA_signal_4769), .A1_t (new_AGEMA_signal_4770), .A1_f (new_AGEMA_signal_4771), .B0_t (Midori_rounds_n14), .B0_f (new_AGEMA_signal_5461), .B1_t (new_AGEMA_signal_5462), .B1_f (new_AGEMA_signal_5463), .Z0_t (Midori_rounds_sub_ResultXORkey[56]), .Z0_f (new_AGEMA_signal_5607), .Z1_t (new_AGEMA_signal_5608), .Z1_f (new_AGEMA_signal_5609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U137 ( .A0_t (Midori_rounds_SR_Inv_Result[20]), .A0_f (new_AGEMA_signal_6800), .A1_t (new_AGEMA_signal_6801), .A1_f (new_AGEMA_signal_6802), .B0_t (Midori_rounds_n14), .B0_f (new_AGEMA_signal_5461), .B1_t (new_AGEMA_signal_5462), .B1_f (new_AGEMA_signal_5463), .Z0_t (Midori_rounds_mul_ResultXORkey[56]), .Z0_f (new_AGEMA_signal_6824), .Z1_t (new_AGEMA_signal_6825), .Z1_f (new_AGEMA_signal_6826) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U136 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[14]), .A1_f (new_AGEMA_signal_5354), .B0_t (Midori_rounds_SelectedKey[56]), .B0_f (new_AGEMA_signal_4256), .B1_t (new_AGEMA_signal_4257), .B1_f (new_AGEMA_signal_4258), .Z0_t (Midori_rounds_n14), .Z0_f (new_AGEMA_signal_5461), .Z1_t (new_AGEMA_signal_5462), .Z1_f (new_AGEMA_signal_5463) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U135 ( .A0_t (Midori_rounds_SR_Result[4]), .A0_f (new_AGEMA_signal_4763), .A1_t (new_AGEMA_signal_4764), .A1_f (new_AGEMA_signal_4765), .B0_t (Midori_rounds_n13), .B0_f (new_AGEMA_signal_5610), .B1_t (new_AGEMA_signal_5611), .B1_f (new_AGEMA_signal_5612), .Z0_t (Midori_rounds_sub_ResultXORkey[52]), .Z0_f (new_AGEMA_signal_5788), .Z1_t (new_AGEMA_signal_5789), .Z1_f (new_AGEMA_signal_5790) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U134 ( .A0_t (Midori_rounds_SR_Inv_Result[40]), .A0_f (new_AGEMA_signal_6761), .A1_t (new_AGEMA_signal_6762), .A1_f (new_AGEMA_signal_6763), .B0_t (Midori_rounds_n13), .B0_f (new_AGEMA_signal_5610), .B1_t (new_AGEMA_signal_5611), .B1_f (new_AGEMA_signal_5612), .Z0_t (Midori_rounds_mul_ResultXORkey[52]), .Z0_f (new_AGEMA_signal_6785), .Z1_t (new_AGEMA_signal_6786), .Z1_f (new_AGEMA_signal_6787) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U133 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[13]), .A1_f (new_AGEMA_signal_5477), .B0_t (Midori_rounds_SelectedKey[52]), .B0_f (new_AGEMA_signal_4244), .B1_t (new_AGEMA_signal_4245), .B1_f (new_AGEMA_signal_4246), .Z0_t (Midori_rounds_n13), .Z0_f (new_AGEMA_signal_5610), .Z1_t (new_AGEMA_signal_5611), .Z1_f (new_AGEMA_signal_5612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U132 ( .A0_t (Midori_rounds_SR_Result[20]), .A0_f (new_AGEMA_signal_4700), .A1_t (new_AGEMA_signal_4701), .A1_f (new_AGEMA_signal_4702), .B0_t (Midori_rounds_n12), .B0_f (new_AGEMA_signal_5613), .B1_t (new_AGEMA_signal_5614), .B1_f (new_AGEMA_signal_5615), .Z0_t (Midori_rounds_sub_ResultXORkey[12]), .Z0_f (new_AGEMA_signal_5791), .Z1_t (new_AGEMA_signal_5792), .Z1_f (new_AGEMA_signal_5793) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U131 ( .A0_t (Midori_rounds_SR_Inv_Result[32]), .A0_f (new_AGEMA_signal_6842), .A1_t (new_AGEMA_signal_6843), .A1_f (new_AGEMA_signal_6844), .B0_t (Midori_rounds_n12), .B0_f (new_AGEMA_signal_5613), .B1_t (new_AGEMA_signal_5614), .B1_f (new_AGEMA_signal_5615), .Z0_t (Midori_rounds_mul_ResultXORkey[12]), .Z0_f (new_AGEMA_signal_6866), .Z1_t (new_AGEMA_signal_6867), .Z1_f (new_AGEMA_signal_6868) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U130 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[3]), .A1_f (new_AGEMA_signal_5473), .B0_t (Midori_rounds_SelectedKey[12]), .B0_f (new_AGEMA_signal_4124), .B1_t (new_AGEMA_signal_4125), .B1_f (new_AGEMA_signal_4126), .Z0_t (Midori_rounds_n12), .Z0_f (new_AGEMA_signal_5613), .Z1_t (new_AGEMA_signal_5614), .Z1_f (new_AGEMA_signal_5615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U129 ( .A0_t (Midori_rounds_SR_Result[16]), .A0_f (new_AGEMA_signal_4739), .A1_t (new_AGEMA_signal_4740), .A1_f (new_AGEMA_signal_4741), .B0_t (Midori_rounds_n11), .B0_f (new_AGEMA_signal_5616), .B1_t (new_AGEMA_signal_5617), .B1_f (new_AGEMA_signal_5618), .Z0_t (Midori_rounds_sub_ResultXORkey[36]), .Z0_f (new_AGEMA_signal_5794), .Z1_t (new_AGEMA_signal_5795), .Z1_f (new_AGEMA_signal_5796) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U128 ( .A0_t (Midori_rounds_SR_Inv_Result[16]), .A0_f (new_AGEMA_signal_6767), .A1_t (new_AGEMA_signal_6768), .A1_f (new_AGEMA_signal_6769), .B0_t (Midori_rounds_n11), .B0_f (new_AGEMA_signal_5616), .B1_t (new_AGEMA_signal_5617), .B1_f (new_AGEMA_signal_5618), .Z0_t (Midori_rounds_mul_ResultXORkey[36]), .Z0_f (new_AGEMA_signal_6788), .Z1_t (new_AGEMA_signal_6789), .Z1_f (new_AGEMA_signal_6790) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U127 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[9]), .A1_f (new_AGEMA_signal_5474), .B0_t (Midori_rounds_SelectedKey[36]), .B0_f (new_AGEMA_signal_4196), .B1_t (new_AGEMA_signal_4197), .B1_f (new_AGEMA_signal_4198), .Z0_t (Midori_rounds_n11), .Z0_f (new_AGEMA_signal_5616), .Z1_t (new_AGEMA_signal_5617), .Z1_f (new_AGEMA_signal_5618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U126 ( .A0_t (Midori_rounds_SR_Result[24]), .A0_f (new_AGEMA_signal_4754), .A1_t (new_AGEMA_signal_4755), .A1_f (new_AGEMA_signal_4756), .B0_t (Midori_rounds_n10), .B0_f (new_AGEMA_signal_5797), .B1_t (new_AGEMA_signal_5798), .B1_f (new_AGEMA_signal_5799), .Z0_t (Midori_rounds_sub_ResultXORkey[48]), .Z0_f (new_AGEMA_signal_5981), .Z1_t (new_AGEMA_signal_5982), .Z1_f (new_AGEMA_signal_5983) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U125 ( .A0_t (Midori_rounds_SR_Inv_Result[0]), .A0_f (new_AGEMA_signal_6689), .A1_t (new_AGEMA_signal_6690), .A1_f (new_AGEMA_signal_6691), .B0_t (Midori_rounds_n10), .B0_f (new_AGEMA_signal_5797), .B1_t (new_AGEMA_signal_5798), .B1_f (new_AGEMA_signal_5799), .Z0_t (Midori_rounds_mul_ResultXORkey[48]), .Z0_f (new_AGEMA_signal_6701), .Z1_t (new_AGEMA_signal_6702), .Z1_f (new_AGEMA_signal_6703) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U124 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[12]), .A1_f (new_AGEMA_signal_5730), .B0_t (Midori_rounds_SelectedKey[48]), .B0_f (new_AGEMA_signal_4232), .B1_t (new_AGEMA_signal_4233), .B1_f (new_AGEMA_signal_4234), .Z0_t (Midori_rounds_n10), .Z0_f (new_AGEMA_signal_5797), .Z1_t (new_AGEMA_signal_5798), .Z1_f (new_AGEMA_signal_5799) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U123 ( .A0_t (Midori_rounds_SR_Result[12]), .A0_f (new_AGEMA_signal_4733), .A1_t (new_AGEMA_signal_4734), .A1_f (new_AGEMA_signal_4735), .B0_t (Midori_rounds_n9), .B0_f (new_AGEMA_signal_5800), .B1_t (new_AGEMA_signal_5801), .B1_f (new_AGEMA_signal_5802), .Z0_t (Midori_rounds_sub_ResultXORkey[32]), .Z0_f (new_AGEMA_signal_5984), .Z1_t (new_AGEMA_signal_5985), .Z1_f (new_AGEMA_signal_5986) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U122 ( .A0_t (Midori_rounds_SR_Inv_Result[56]), .A0_f (new_AGEMA_signal_6692), .A1_t (new_AGEMA_signal_6693), .A1_f (new_AGEMA_signal_6694), .B0_t (Midori_rounds_n9), .B0_f (new_AGEMA_signal_5800), .B1_t (new_AGEMA_signal_5801), .B1_f (new_AGEMA_signal_5802), .Z0_t (Midori_rounds_mul_ResultXORkey[32]), .Z0_f (new_AGEMA_signal_6704), .Z1_t (new_AGEMA_signal_6705), .Z1_f (new_AGEMA_signal_6706) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U121 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[8]), .A1_f (new_AGEMA_signal_5733), .B0_t (Midori_rounds_SelectedKey[32]), .B0_f (new_AGEMA_signal_4184), .B1_t (new_AGEMA_signal_4185), .B1_f (new_AGEMA_signal_4186), .Z0_t (Midori_rounds_n9), .Z0_f (new_AGEMA_signal_5800), .Z1_t (new_AGEMA_signal_5801), .Z1_f (new_AGEMA_signal_5802) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U120 ( .A0_t (Midori_rounds_SR_Result[0]), .A0_f (new_AGEMA_signal_4727), .A1_t (new_AGEMA_signal_4728), .A1_f (new_AGEMA_signal_4729), .B0_t (Midori_rounds_n8), .B0_f (new_AGEMA_signal_5619), .B1_t (new_AGEMA_signal_5620), .B1_f (new_AGEMA_signal_5621), .Z0_t (Midori_rounds_sub_ResultXORkey[28]), .Z0_f (new_AGEMA_signal_5803), .Z1_t (new_AGEMA_signal_5804), .Z1_f (new_AGEMA_signal_5805) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U119 ( .A0_t (Midori_rounds_SR_Inv_Result[24]), .A0_f (new_AGEMA_signal_6809), .A1_t (new_AGEMA_signal_6810), .A1_f (new_AGEMA_signal_6811), .B0_t (Midori_rounds_n8), .B0_f (new_AGEMA_signal_5619), .B1_t (new_AGEMA_signal_5620), .B1_f (new_AGEMA_signal_5621), .Z0_t (Midori_rounds_mul_ResultXORkey[28]), .Z0_f (new_AGEMA_signal_6827), .Z1_t (new_AGEMA_signal_6828), .Z1_f (new_AGEMA_signal_6829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U118 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[7]), .A1_f (new_AGEMA_signal_5475), .B0_t (Midori_rounds_SelectedKey[28]), .B0_f (new_AGEMA_signal_4172), .B1_t (new_AGEMA_signal_4173), .B1_f (new_AGEMA_signal_4174), .Z0_t (Midori_rounds_n8), .Z0_f (new_AGEMA_signal_5619), .Z1_t (new_AGEMA_signal_5620), .Z1_f (new_AGEMA_signal_5621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U117 ( .A0_t (Midori_rounds_SR_Result[40]), .A0_f (new_AGEMA_signal_4748), .A1_t (new_AGEMA_signal_4749), .A1_f (new_AGEMA_signal_4750), .B0_t (Midori_rounds_n7), .B0_f (new_AGEMA_signal_5188), .B1_t (new_AGEMA_signal_5189), .B1_f (new_AGEMA_signal_5190), .Z0_t (Midori_rounds_sub_ResultXORkey[44]), .Z0_f (new_AGEMA_signal_5345), .Z1_t (new_AGEMA_signal_5346), .Z1_f (new_AGEMA_signal_5347) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U116 ( .A0_t (Midori_rounds_SR_Inv_Result[4]), .A0_f (new_AGEMA_signal_6803), .A1_t (new_AGEMA_signal_6804), .A1_f (new_AGEMA_signal_6805), .B0_t (Midori_rounds_n7), .B0_f (new_AGEMA_signal_5188), .B1_t (new_AGEMA_signal_5189), .B1_f (new_AGEMA_signal_5190), .Z0_t (Midori_rounds_mul_ResultXORkey[44]), .Z0_f (new_AGEMA_signal_6830), .Z1_t (new_AGEMA_signal_6831), .Z1_f (new_AGEMA_signal_6832) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U115 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[11]), .A1_f (new_AGEMA_signal_5033), .B0_t (Midori_rounds_SelectedKey[44]), .B0_f (new_AGEMA_signal_4220), .B1_t (new_AGEMA_signal_4221), .B1_f (new_AGEMA_signal_4222), .Z0_t (Midori_rounds_n7), .Z0_f (new_AGEMA_signal_5188), .Z1_t (new_AGEMA_signal_5189), .Z1_f (new_AGEMA_signal_5190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U114 ( .A0_t (Midori_rounds_SR_Result[28]), .A0_f (new_AGEMA_signal_4718), .A1_t (new_AGEMA_signal_4719), .A1_f (new_AGEMA_signal_4720), .B0_t (Midori_rounds_n6), .B0_f (new_AGEMA_signal_5348), .B1_t (new_AGEMA_signal_5349), .B1_f (new_AGEMA_signal_5350), .Z0_t (Midori_rounds_sub_ResultXORkey[24]), .Z0_f (new_AGEMA_signal_5464), .Z1_t (new_AGEMA_signal_5465), .Z1_f (new_AGEMA_signal_5466) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U113 ( .A0_t (Midori_rounds_SR_Inv_Result[48]), .A0_f (new_AGEMA_signal_6812), .A1_t (new_AGEMA_signal_6813), .A1_f (new_AGEMA_signal_6814), .B0_t (Midori_rounds_n6), .B0_f (new_AGEMA_signal_5348), .B1_t (new_AGEMA_signal_5349), .B1_f (new_AGEMA_signal_5350), .Z0_t (Midori_rounds_mul_ResultXORkey[24]), .Z0_f (new_AGEMA_signal_6833), .Z1_t (new_AGEMA_signal_6834), .Z1_f (new_AGEMA_signal_6835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U112 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[6]), .A1_f (new_AGEMA_signal_5196), .B0_t (Midori_rounds_SelectedKey[24]), .B0_f (new_AGEMA_signal_4160), .B1_t (new_AGEMA_signal_4161), .B1_f (new_AGEMA_signal_4162), .Z0_t (Midori_rounds_n6), .Z0_f (new_AGEMA_signal_5348), .Z1_t (new_AGEMA_signal_5349), .Z1_f (new_AGEMA_signal_5350) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U111 ( .A0_t (Midori_rounds_SR_Result[8]), .A0_f (new_AGEMA_signal_4694), .A1_t (new_AGEMA_signal_4695), .A1_f (new_AGEMA_signal_4696), .B0_t (Midori_rounds_n5), .B0_f (new_AGEMA_signal_5622), .B1_t (new_AGEMA_signal_5623), .B1_f (new_AGEMA_signal_5624), .Z0_t (Midori_rounds_sub_ResultXORkey[8]), .Z0_f (new_AGEMA_signal_5806), .Z1_t (new_AGEMA_signal_5807), .Z1_f (new_AGEMA_signal_5808) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U110 ( .A0_t (Midori_rounds_SR_Inv_Result[8]), .A0_f (new_AGEMA_signal_6845), .A1_t (new_AGEMA_signal_6846), .A1_f (new_AGEMA_signal_6847), .B0_t (Midori_rounds_n5), .B0_f (new_AGEMA_signal_5622), .B1_t (new_AGEMA_signal_5623), .B1_f (new_AGEMA_signal_5624), .Z0_t (Midori_rounds_mul_ResultXORkey[8]), .Z0_f (new_AGEMA_signal_6869), .Z1_t (new_AGEMA_signal_6870), .Z1_f (new_AGEMA_signal_6871) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U109 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[2]), .A1_f (new_AGEMA_signal_5478), .B0_t (Midori_rounds_SelectedKey[8]), .B0_f (new_AGEMA_signal_4112), .B1_t (new_AGEMA_signal_4113), .B1_f (new_AGEMA_signal_4114), .Z0_t (Midori_rounds_n5), .Z0_f (new_AGEMA_signal_5622), .Z1_t (new_AGEMA_signal_5623), .Z1_f (new_AGEMA_signal_5624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U108 ( .A0_t (Midori_rounds_SR_Result[48]), .A0_f (new_AGEMA_signal_4685), .A1_t (new_AGEMA_signal_4686), .A1_f (new_AGEMA_signal_4687), .B0_t (Midori_rounds_n4), .B0_f (new_AGEMA_signal_5625), .B1_t (new_AGEMA_signal_5626), .B1_f (new_AGEMA_signal_5627), .Z0_t (Midori_rounds_sub_ResultXORkey[0]), .Z0_f (new_AGEMA_signal_5809), .Z1_t (new_AGEMA_signal_5810), .Z1_f (new_AGEMA_signal_5811) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U107 ( .A0_t (Midori_rounds_SR_Inv_Result[28]), .A0_f (new_AGEMA_signal_6818), .A1_t (new_AGEMA_signal_6819), .A1_f (new_AGEMA_signal_6820), .B0_t (Midori_rounds_n4), .B0_f (new_AGEMA_signal_5625), .B1_t (new_AGEMA_signal_5626), .B1_f (new_AGEMA_signal_5627), .Z0_t (Midori_rounds_mul_ResultXORkey[0]), .Z0_f (new_AGEMA_signal_6836), .Z1_t (new_AGEMA_signal_6837), .Z1_f (new_AGEMA_signal_6838) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U106 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[0]), .A1_f (new_AGEMA_signal_5479), .B0_t (Midori_rounds_SelectedKey[0]), .B0_f (new_AGEMA_signal_4088), .B1_t (new_AGEMA_signal_4089), .B1_f (new_AGEMA_signal_4090), .Z0_t (Midori_rounds_n4), .Z0_f (new_AGEMA_signal_5625), .Z1_t (new_AGEMA_signal_5626), .Z1_f (new_AGEMA_signal_5627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U105 ( .A0_t (Midori_rounds_SR_Result[52]), .A0_f (new_AGEMA_signal_4742), .A1_t (new_AGEMA_signal_4743), .A1_f (new_AGEMA_signal_4744), .B0_t (Midori_rounds_n3), .B0_f (new_AGEMA_signal_5467), .B1_t (new_AGEMA_signal_5468), .B1_f (new_AGEMA_signal_5469), .Z0_t (Midori_rounds_sub_ResultXORkey[40]), .Z0_f (new_AGEMA_signal_5628), .Z1_t (new_AGEMA_signal_5629), .Z1_f (new_AGEMA_signal_5630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U104 ( .A0_t (Midori_rounds_SR_Inv_Result[44]), .A0_f (new_AGEMA_signal_6806), .A1_t (new_AGEMA_signal_6807), .A1_f (new_AGEMA_signal_6808), .B0_t (Midori_rounds_n3), .B0_f (new_AGEMA_signal_5467), .B1_t (new_AGEMA_signal_5468), .B1_f (new_AGEMA_signal_5469), .Z0_t (Midori_rounds_mul_ResultXORkey[40]), .Z0_f (new_AGEMA_signal_6839), .Z1_t (new_AGEMA_signal_6840), .Z1_f (new_AGEMA_signal_6841) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U103 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[10]), .A1_f (new_AGEMA_signal_5355), .B0_t (Midori_rounds_SelectedKey[40]), .B0_f (new_AGEMA_signal_4208), .B1_t (new_AGEMA_signal_4209), .B1_f (new_AGEMA_signal_4210), .Z0_t (Midori_rounds_n3), .Z0_f (new_AGEMA_signal_5467), .Z1_t (new_AGEMA_signal_5468), .Z1_f (new_AGEMA_signal_5469) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U102 ( .A0_t (Midori_rounds_SR_Result[56]), .A0_f (new_AGEMA_signal_4712), .A1_t (new_AGEMA_signal_4713), .A1_f (new_AGEMA_signal_4714), .B0_t (Midori_rounds_n2), .B0_f (new_AGEMA_signal_5470), .B1_t (new_AGEMA_signal_5471), .B1_f (new_AGEMA_signal_5472), .Z0_t (Midori_rounds_sub_ResultXORkey[20]), .Z0_f (new_AGEMA_signal_5631), .Z1_t (new_AGEMA_signal_5632), .Z1_f (new_AGEMA_signal_5633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U101 ( .A0_t (Midori_rounds_SR_Inv_Result[12]), .A0_f (new_AGEMA_signal_6773), .A1_t (new_AGEMA_signal_6774), .A1_f (new_AGEMA_signal_6775), .B0_t (Midori_rounds_n2), .B0_f (new_AGEMA_signal_5470), .B1_t (new_AGEMA_signal_5471), .B1_f (new_AGEMA_signal_5472), .Z0_t (Midori_rounds_mul_ResultXORkey[20]), .Z0_f (new_AGEMA_signal_6791), .Z1_t (new_AGEMA_signal_6792), .Z1_f (new_AGEMA_signal_6793) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U100 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[5]), .A1_f (new_AGEMA_signal_5356), .B0_t (Midori_rounds_SelectedKey[20]), .B0_f (new_AGEMA_signal_4148), .B1_t (new_AGEMA_signal_4149), .B1_f (new_AGEMA_signal_4150), .Z0_t (Midori_rounds_n2), .Z0_f (new_AGEMA_signal_5470), .Z1_t (new_AGEMA_signal_5471), .Z1_f (new_AGEMA_signal_5472) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U99 ( .A0_t (Midori_rounds_SR_Result[36]), .A0_f (new_AGEMA_signal_4706), .A1_t (new_AGEMA_signal_4707), .A1_f (new_AGEMA_signal_4708), .B0_t (Midori_rounds_n1), .B0_f (new_AGEMA_signal_5812), .B1_t (new_AGEMA_signal_5813), .B1_f (new_AGEMA_signal_5814), .Z0_t (Midori_rounds_sub_ResultXORkey[16]), .Z0_f (new_AGEMA_signal_5987), .Z1_t (new_AGEMA_signal_5988), .Z1_f (new_AGEMA_signal_5989) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U98 ( .A0_t (Midori_rounds_SR_Inv_Result[36]), .A0_f (new_AGEMA_signal_6776), .A1_t (new_AGEMA_signal_6777), .A1_f (new_AGEMA_signal_6778), .B0_t (Midori_rounds_n1), .B0_f (new_AGEMA_signal_5812), .B1_t (new_AGEMA_signal_5813), .B1_f (new_AGEMA_signal_5814), .Z0_t (Midori_rounds_mul_ResultXORkey[16]), .Z0_f (new_AGEMA_signal_6794), .Z1_t (new_AGEMA_signal_6795), .Z1_f (new_AGEMA_signal_6796) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U97 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Midori_rounds_round_Constant[4]), .A1_f (new_AGEMA_signal_5732), .B0_t (Midori_rounds_SelectedKey[16]), .B0_f (new_AGEMA_signal_4136), .B1_t (new_AGEMA_signal_4137), .B1_f (new_AGEMA_signal_4138), .Z0_t (Midori_rounds_n1), .Z0_f (new_AGEMA_signal_5812), .Z1_t (new_AGEMA_signal_5813), .Z1_f (new_AGEMA_signal_5814) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U96 ( .A0_t (Midori_rounds_SelectedKey[51]), .A0_f (new_AGEMA_signal_4241), .A1_t (new_AGEMA_signal_4242), .A1_f (new_AGEMA_signal_4243), .B0_t (Midori_rounds_SR_Result[27]), .B0_f (new_AGEMA_signal_4430), .B1_t (new_AGEMA_signal_4431), .B1_f (new_AGEMA_signal_4432), .Z0_t (Midori_rounds_sub_ResultXORkey[51]), .Z0_f (new_AGEMA_signal_4570), .Z1_t (new_AGEMA_signal_4571), .Z1_f (new_AGEMA_signal_4572) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U95 ( .A0_t (Midori_rounds_SelectedKey[54]), .A0_f (new_AGEMA_signal_4250), .A1_t (new_AGEMA_signal_4251), .A1_f (new_AGEMA_signal_4252), .B0_t (Midori_rounds_SR_Result[6]), .B0_f (new_AGEMA_signal_4760), .B1_t (new_AGEMA_signal_4761), .B1_f (new_AGEMA_signal_4762), .Z0_t (Midori_rounds_sub_ResultXORkey[54]), .Z0_f (new_AGEMA_signal_4875), .Z1_t (new_AGEMA_signal_4876), .Z1_f (new_AGEMA_signal_4877) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U94 ( .A0_t (Midori_rounds_SelectedKey[49]), .A0_f (new_AGEMA_signal_4235), .A1_t (new_AGEMA_signal_4236), .A1_f (new_AGEMA_signal_4237), .B0_t (Midori_rounds_SR_Result[25]), .B0_f (new_AGEMA_signal_4433), .B1_t (new_AGEMA_signal_4434), .B1_f (new_AGEMA_signal_4435), .Z0_t (Midori_rounds_sub_ResultXORkey[49]), .Z0_f (new_AGEMA_signal_4573), .Z1_t (new_AGEMA_signal_4574), .Z1_f (new_AGEMA_signal_4575) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U93 ( .A0_t (Midori_rounds_SelectedKey[39]), .A0_f (new_AGEMA_signal_4205), .A1_t (new_AGEMA_signal_4206), .A1_f (new_AGEMA_signal_4207), .B0_t (Midori_rounds_SR_Result[19]), .B0_f (new_AGEMA_signal_4388), .B1_t (new_AGEMA_signal_4389), .B1_f (new_AGEMA_signal_4390), .Z0_t (Midori_rounds_sub_ResultXORkey[39]), .Z0_f (new_AGEMA_signal_4576), .Z1_t (new_AGEMA_signal_4577), .Z1_f (new_AGEMA_signal_4578) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U92 ( .A0_t (Midori_rounds_SelectedKey[37]), .A0_f (new_AGEMA_signal_4199), .A1_t (new_AGEMA_signal_4200), .A1_f (new_AGEMA_signal_4201), .B0_t (Midori_rounds_SR_Result[17]), .B0_f (new_AGEMA_signal_4391), .B1_t (new_AGEMA_signal_4392), .B1_f (new_AGEMA_signal_4393), .Z0_t (Midori_rounds_sub_ResultXORkey[37]), .Z0_f (new_AGEMA_signal_4579), .Z1_t (new_AGEMA_signal_4580), .Z1_f (new_AGEMA_signal_4581) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U91 ( .A0_t (Midori_rounds_SelectedKey[19]), .A0_f (new_AGEMA_signal_4145), .A1_t (new_AGEMA_signal_4146), .A1_f (new_AGEMA_signal_4147), .B0_t (Midori_rounds_SR_Result[39]), .B0_f (new_AGEMA_signal_4334), .B1_t (new_AGEMA_signal_4335), .B1_f (new_AGEMA_signal_4336), .Z0_t (Midori_rounds_sub_ResultXORkey[19]), .Z0_f (new_AGEMA_signal_4582), .Z1_t (new_AGEMA_signal_4583), .Z1_f (new_AGEMA_signal_4584) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U90 ( .A0_t (Midori_rounds_SelectedKey[17]), .A0_f (new_AGEMA_signal_4139), .A1_t (new_AGEMA_signal_4140), .A1_f (new_AGEMA_signal_4141), .B0_t (Midori_rounds_SR_Result[37]), .B0_f (new_AGEMA_signal_4337), .B1_t (new_AGEMA_signal_4338), .B1_f (new_AGEMA_signal_4339), .Z0_t (Midori_rounds_sub_ResultXORkey[17]), .Z0_f (new_AGEMA_signal_4585), .Z1_t (new_AGEMA_signal_4586), .Z1_f (new_AGEMA_signal_4587) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U89 ( .A0_t (Midori_rounds_SelectedKey[34]), .A0_f (new_AGEMA_signal_4190), .A1_t (new_AGEMA_signal_4191), .A1_f (new_AGEMA_signal_4192), .B0_t (Midori_rounds_SR_Result[14]), .B0_f (new_AGEMA_signal_4730), .B1_t (new_AGEMA_signal_4731), .B1_f (new_AGEMA_signal_4732), .Z0_t (Midori_rounds_sub_ResultXORkey[34]), .Z0_f (new_AGEMA_signal_4878), .Z1_t (new_AGEMA_signal_4879), .Z1_f (new_AGEMA_signal_4880) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U88 ( .A0_t (Midori_rounds_SelectedKey[18]), .A0_f (new_AGEMA_signal_4142), .A1_t (new_AGEMA_signal_4143), .A1_f (new_AGEMA_signal_4144), .B0_t (Midori_rounds_SR_Result[38]), .B0_f (new_AGEMA_signal_4709), .B1_t (new_AGEMA_signal_4710), .B1_f (new_AGEMA_signal_4711), .Z0_t (Midori_rounds_sub_ResultXORkey[18]), .Z0_f (new_AGEMA_signal_4881), .Z1_t (new_AGEMA_signal_4882), .Z1_f (new_AGEMA_signal_4883) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U87 ( .A0_t (Midori_rounds_SelectedKey[55]), .A0_f (new_AGEMA_signal_4253), .A1_t (new_AGEMA_signal_4254), .A1_f (new_AGEMA_signal_4255), .B0_t (Midori_rounds_SR_Result[7]), .B0_f (new_AGEMA_signal_4436), .B1_t (new_AGEMA_signal_4437), .B1_f (new_AGEMA_signal_4438), .Z0_t (Midori_rounds_sub_ResultXORkey[55]), .Z0_f (new_AGEMA_signal_4588), .Z1_t (new_AGEMA_signal_4589), .Z1_f (new_AGEMA_signal_4590) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U86 ( .A0_t (Midori_rounds_SelectedKey[50]), .A0_f (new_AGEMA_signal_4238), .A1_t (new_AGEMA_signal_4239), .A1_f (new_AGEMA_signal_4240), .B0_t (Midori_rounds_SR_Result[26]), .B0_f (new_AGEMA_signal_4757), .B1_t (new_AGEMA_signal_4758), .B1_f (new_AGEMA_signal_4759), .Z0_t (Midori_rounds_sub_ResultXORkey[50]), .Z0_f (new_AGEMA_signal_4884), .Z1_t (new_AGEMA_signal_4885), .Z1_f (new_AGEMA_signal_4886) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U85 ( .A0_t (Midori_rounds_SelectedKey[53]), .A0_f (new_AGEMA_signal_4247), .A1_t (new_AGEMA_signal_4248), .A1_f (new_AGEMA_signal_4249), .B0_t (Midori_rounds_SR_Result[5]), .B0_f (new_AGEMA_signal_4439), .B1_t (new_AGEMA_signal_4440), .B1_f (new_AGEMA_signal_4441), .Z0_t (Midori_rounds_sub_ResultXORkey[53]), .Z0_f (new_AGEMA_signal_4591), .Z1_t (new_AGEMA_signal_4592), .Z1_f (new_AGEMA_signal_4593) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U84 ( .A0_t (Midori_rounds_SelectedKey[35]), .A0_f (new_AGEMA_signal_4193), .A1_t (new_AGEMA_signal_4194), .A1_f (new_AGEMA_signal_4195), .B0_t (Midori_rounds_SR_Result[15]), .B0_f (new_AGEMA_signal_4376), .B1_t (new_AGEMA_signal_4377), .B1_f (new_AGEMA_signal_4378), .Z0_t (Midori_rounds_sub_ResultXORkey[35]), .Z0_f (new_AGEMA_signal_4594), .Z1_t (new_AGEMA_signal_4595), .Z1_f (new_AGEMA_signal_4596) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U83 ( .A0_t (Midori_rounds_SelectedKey[38]), .A0_f (new_AGEMA_signal_4202), .A1_t (new_AGEMA_signal_4203), .A1_f (new_AGEMA_signal_4204), .B0_t (Midori_rounds_SR_Result[18]), .B0_f (new_AGEMA_signal_4736), .B1_t (new_AGEMA_signal_4737), .B1_f (new_AGEMA_signal_4738), .Z0_t (Midori_rounds_sub_ResultXORkey[38]), .Z0_f (new_AGEMA_signal_4887), .Z1_t (new_AGEMA_signal_4888), .Z1_f (new_AGEMA_signal_4889) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U82 ( .A0_t (Midori_rounds_SelectedKey[33]), .A0_f (new_AGEMA_signal_4187), .A1_t (new_AGEMA_signal_4188), .A1_f (new_AGEMA_signal_4189), .B0_t (Midori_rounds_SR_Result[13]), .B0_f (new_AGEMA_signal_4379), .B1_t (new_AGEMA_signal_4380), .B1_f (new_AGEMA_signal_4381), .Z0_t (Midori_rounds_sub_ResultXORkey[33]), .Z0_f (new_AGEMA_signal_4597), .Z1_t (new_AGEMA_signal_4598), .Z1_f (new_AGEMA_signal_4599) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U81 ( .A0_t (Midori_rounds_SelectedKey[23]), .A0_f (new_AGEMA_signal_4157), .A1_t (new_AGEMA_signal_4158), .A1_f (new_AGEMA_signal_4159), .B0_t (Midori_rounds_SR_Result[59]), .B0_f (new_AGEMA_signal_4346), .B1_t (new_AGEMA_signal_4347), .B1_f (new_AGEMA_signal_4348), .Z0_t (Midori_rounds_sub_ResultXORkey[23]), .Z0_f (new_AGEMA_signal_4600), .Z1_t (new_AGEMA_signal_4601), .Z1_f (new_AGEMA_signal_4602) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U80 ( .A0_t (Midori_rounds_SelectedKey[22]), .A0_f (new_AGEMA_signal_4154), .A1_t (new_AGEMA_signal_4155), .A1_f (new_AGEMA_signal_4156), .B0_t (Midori_rounds_SR_Result[58]), .B0_f (new_AGEMA_signal_4715), .B1_t (new_AGEMA_signal_4716), .B1_f (new_AGEMA_signal_4717), .Z0_t (Midori_rounds_sub_ResultXORkey[22]), .Z0_f (new_AGEMA_signal_4890), .Z1_t (new_AGEMA_signal_4891), .Z1_f (new_AGEMA_signal_4892) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U79 ( .A0_t (Midori_rounds_SelectedKey[21]), .A0_f (new_AGEMA_signal_4151), .A1_t (new_AGEMA_signal_4152), .A1_f (new_AGEMA_signal_4153), .B0_t (Midori_rounds_SR_Result[57]), .B0_f (new_AGEMA_signal_4349), .B1_t (new_AGEMA_signal_4350), .B1_f (new_AGEMA_signal_4351), .Z0_t (Midori_rounds_sub_ResultXORkey[21]), .Z0_f (new_AGEMA_signal_4603), .Z1_t (new_AGEMA_signal_4604), .Z1_f (new_AGEMA_signal_4605) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U78 ( .A0_t (Midori_rounds_SelectedKey[7]), .A0_f (new_AGEMA_signal_4109), .A1_t (new_AGEMA_signal_4110), .A1_f (new_AGEMA_signal_4111), .B0_t (Midori_rounds_SR_Result[47]), .B0_f (new_AGEMA_signal_4298), .B1_t (new_AGEMA_signal_4299), .B1_f (new_AGEMA_signal_4300), .Z0_t (Midori_rounds_sub_ResultXORkey[7]), .Z0_f (new_AGEMA_signal_4606), .Z1_t (new_AGEMA_signal_4607), .Z1_f (new_AGEMA_signal_4608) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U77 ( .A0_t (Midori_rounds_SelectedKey[2]), .A0_f (new_AGEMA_signal_4094), .A1_t (new_AGEMA_signal_4095), .A1_f (new_AGEMA_signal_4096), .B0_t (Midori_rounds_SR_Result[50]), .B0_f (new_AGEMA_signal_4682), .B1_t (new_AGEMA_signal_4683), .B1_f (new_AGEMA_signal_4684), .Z0_t (Midori_rounds_sub_ResultXORkey[2]), .Z0_f (new_AGEMA_signal_4893), .Z1_t (new_AGEMA_signal_4894), .Z1_f (new_AGEMA_signal_4895) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U76 ( .A0_t (Midori_rounds_SelectedKey[5]), .A0_f (new_AGEMA_signal_4103), .A1_t (new_AGEMA_signal_4104), .A1_f (new_AGEMA_signal_4105), .B0_t (Midori_rounds_SR_Result[45]), .B0_f (new_AGEMA_signal_4301), .B1_t (new_AGEMA_signal_4302), .B1_f (new_AGEMA_signal_4303), .Z0_t (Midori_rounds_sub_ResultXORkey[5]), .Z0_f (new_AGEMA_signal_4609), .Z1_t (new_AGEMA_signal_4610), .Z1_f (new_AGEMA_signal_4611) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U75 ( .A0_t (Midori_rounds_SelectedKey[3]), .A0_f (new_AGEMA_signal_4097), .A1_t (new_AGEMA_signal_4098), .A1_f (new_AGEMA_signal_4099), .B0_t (Midori_rounds_SR_Result[51]), .B0_f (new_AGEMA_signal_4280), .B1_t (new_AGEMA_signal_4281), .B1_f (new_AGEMA_signal_4282), .Z0_t (Midori_rounds_sub_ResultXORkey[3]), .Z0_f (new_AGEMA_signal_4612), .Z1_t (new_AGEMA_signal_4613), .Z1_f (new_AGEMA_signal_4614) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U74 ( .A0_t (Midori_rounds_SelectedKey[6]), .A0_f (new_AGEMA_signal_4106), .A1_t (new_AGEMA_signal_4107), .A1_f (new_AGEMA_signal_4108), .B0_t (Midori_rounds_SR_Result[46]), .B0_f (new_AGEMA_signal_4691), .B1_t (new_AGEMA_signal_4692), .B1_f (new_AGEMA_signal_4693), .Z0_t (Midori_rounds_sub_ResultXORkey[6]), .Z0_f (new_AGEMA_signal_4896), .Z1_t (new_AGEMA_signal_4897), .Z1_f (new_AGEMA_signal_4898) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U73 ( .A0_t (Midori_rounds_SelectedKey[1]), .A0_f (new_AGEMA_signal_4091), .A1_t (new_AGEMA_signal_4092), .A1_f (new_AGEMA_signal_4093), .B0_t (Midori_rounds_SR_Result[49]), .B0_f (new_AGEMA_signal_4283), .B1_t (new_AGEMA_signal_4284), .B1_f (new_AGEMA_signal_4285), .Z0_t (Midori_rounds_sub_ResultXORkey[1]), .Z0_f (new_AGEMA_signal_4615), .Z1_t (new_AGEMA_signal_4616), .Z1_f (new_AGEMA_signal_4617) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U72 ( .A0_t (Midori_rounds_SelectedKey[63]), .A0_f (new_AGEMA_signal_4277), .A1_t (new_AGEMA_signal_4278), .A1_f (new_AGEMA_signal_4279), .B0_t (Midori_rounds_SR_Inv_Result[63]), .B0_f (new_AGEMA_signal_5484), .B1_t (new_AGEMA_signal_5485), .B1_f (new_AGEMA_signal_5486), .Z0_t (Midori_rounds_mul_ResultXORkey[63]), .Z0_f (new_AGEMA_signal_5634), .Z1_t (new_AGEMA_signal_5635), .Z1_f (new_AGEMA_signal_5636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U71 ( .A0_t (Midori_rounds_SelectedKey[62]), .A0_f (new_AGEMA_signal_4274), .A1_t (new_AGEMA_signal_4275), .A1_f (new_AGEMA_signal_4276), .B0_t (Midori_rounds_SR_Inv_Result[62]), .B0_f (new_AGEMA_signal_5740), .B1_t (new_AGEMA_signal_5741), .B1_f (new_AGEMA_signal_5742), .Z0_t (Midori_rounds_mul_ResultXORkey[62]), .Z0_f (new_AGEMA_signal_5815), .Z1_t (new_AGEMA_signal_5816), .Z1_f (new_AGEMA_signal_5817) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U70 ( .A0_t (Midori_rounds_SelectedKey[61]), .A0_f (new_AGEMA_signal_4271), .A1_t (new_AGEMA_signal_4272), .A1_f (new_AGEMA_signal_4273), .B0_t (Midori_rounds_SR_Inv_Result[61]), .B0_f (new_AGEMA_signal_5499), .B1_t (new_AGEMA_signal_5500), .B1_f (new_AGEMA_signal_5501), .Z0_t (Midori_rounds_mul_ResultXORkey[61]), .Z0_f (new_AGEMA_signal_5637), .Z1_t (new_AGEMA_signal_5638), .Z1_f (new_AGEMA_signal_5639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U69 ( .A0_t (Midori_rounds_SelectedKey[59]), .A0_f (new_AGEMA_signal_4265), .A1_t (new_AGEMA_signal_4266), .A1_f (new_AGEMA_signal_4267), .B0_t (Midori_rounds_SR_Inv_Result[23]), .B0_f (new_AGEMA_signal_5487), .B1_t (new_AGEMA_signal_5488), .B1_f (new_AGEMA_signal_5489), .Z0_t (Midori_rounds_mul_ResultXORkey[59]), .Z0_f (new_AGEMA_signal_5640), .Z1_t (new_AGEMA_signal_5641), .Z1_f (new_AGEMA_signal_5642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U68 ( .A0_t (Midori_rounds_SelectedKey[58]), .A0_f (new_AGEMA_signal_4262), .A1_t (new_AGEMA_signal_4263), .A1_f (new_AGEMA_signal_4264), .B0_t (Midori_rounds_SR_Inv_Result[22]), .B0_f (new_AGEMA_signal_5743), .B1_t (new_AGEMA_signal_5744), .B1_f (new_AGEMA_signal_5745), .Z0_t (Midori_rounds_mul_ResultXORkey[58]), .Z0_f (new_AGEMA_signal_5818), .Z1_t (new_AGEMA_signal_5819), .Z1_f (new_AGEMA_signal_5820) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U67 ( .A0_t (Midori_rounds_SelectedKey[57]), .A0_f (new_AGEMA_signal_4259), .A1_t (new_AGEMA_signal_4260), .A1_f (new_AGEMA_signal_4261), .B0_t (Midori_rounds_SR_Inv_Result[21]), .B0_f (new_AGEMA_signal_5502), .B1_t (new_AGEMA_signal_5503), .B1_f (new_AGEMA_signal_5504), .Z0_t (Midori_rounds_mul_ResultXORkey[57]), .Z0_f (new_AGEMA_signal_5643), .Z1_t (new_AGEMA_signal_5644), .Z1_f (new_AGEMA_signal_5645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U66 ( .A0_t (Midori_rounds_SelectedKey[55]), .A0_f (new_AGEMA_signal_4253), .A1_t (new_AGEMA_signal_4254), .A1_f (new_AGEMA_signal_4255), .B0_t (Midori_rounds_SR_Inv_Result[43]), .B0_f (new_AGEMA_signal_5493), .B1_t (new_AGEMA_signal_5494), .B1_f (new_AGEMA_signal_5495), .Z0_t (Midori_rounds_mul_ResultXORkey[55]), .Z0_f (new_AGEMA_signal_5646), .Z1_t (new_AGEMA_signal_5647), .Z1_f (new_AGEMA_signal_5648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U65 ( .A0_t (Midori_rounds_SelectedKey[54]), .A0_f (new_AGEMA_signal_4250), .A1_t (new_AGEMA_signal_4251), .A1_f (new_AGEMA_signal_4252), .B0_t (Midori_rounds_SR_Inv_Result[42]), .B0_f (new_AGEMA_signal_5746), .B1_t (new_AGEMA_signal_5747), .B1_f (new_AGEMA_signal_5748), .Z0_t (Midori_rounds_mul_ResultXORkey[54]), .Z0_f (new_AGEMA_signal_5821), .Z1_t (new_AGEMA_signal_5822), .Z1_f (new_AGEMA_signal_5823) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U64 ( .A0_t (Midori_rounds_SelectedKey[53]), .A0_f (new_AGEMA_signal_4247), .A1_t (new_AGEMA_signal_4248), .A1_f (new_AGEMA_signal_4249), .B0_t (Midori_rounds_SR_Inv_Result[41]), .B0_f (new_AGEMA_signal_5508), .B1_t (new_AGEMA_signal_5509), .B1_f (new_AGEMA_signal_5510), .Z0_t (Midori_rounds_mul_ResultXORkey[53]), .Z0_f (new_AGEMA_signal_5649), .Z1_t (new_AGEMA_signal_5650), .Z1_f (new_AGEMA_signal_5651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U63 ( .A0_t (Midori_rounds_SelectedKey[51]), .A0_f (new_AGEMA_signal_4241), .A1_t (new_AGEMA_signal_4242), .A1_f (new_AGEMA_signal_4243), .B0_t (Midori_rounds_SR_Inv_Result[3]), .B0_f (new_AGEMA_signal_5496), .B1_t (new_AGEMA_signal_5497), .B1_f (new_AGEMA_signal_5498), .Z0_t (Midori_rounds_mul_ResultXORkey[51]), .Z0_f (new_AGEMA_signal_5652), .Z1_t (new_AGEMA_signal_5653), .Z1_f (new_AGEMA_signal_5654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U62 ( .A0_t (Midori_rounds_SelectedKey[50]), .A0_f (new_AGEMA_signal_4238), .A1_t (new_AGEMA_signal_4239), .A1_f (new_AGEMA_signal_4240), .B0_t (Midori_rounds_SR_Inv_Result[2]), .B0_f (new_AGEMA_signal_5749), .B1_t (new_AGEMA_signal_5750), .B1_f (new_AGEMA_signal_5751), .Z0_t (Midori_rounds_mul_ResultXORkey[50]), .Z0_f (new_AGEMA_signal_5824), .Z1_t (new_AGEMA_signal_5825), .Z1_f (new_AGEMA_signal_5826) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U61 ( .A0_t (Midori_rounds_SelectedKey[49]), .A0_f (new_AGEMA_signal_4235), .A1_t (new_AGEMA_signal_4236), .A1_f (new_AGEMA_signal_4237), .B0_t (Midori_rounds_SR_Inv_Result[1]), .B0_f (new_AGEMA_signal_5511), .B1_t (new_AGEMA_signal_5512), .B1_f (new_AGEMA_signal_5513), .Z0_t (Midori_rounds_mul_ResultXORkey[49]), .Z0_f (new_AGEMA_signal_5655), .Z1_t (new_AGEMA_signal_5656), .Z1_f (new_AGEMA_signal_5657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U60 ( .A0_t (Midori_rounds_SelectedKey[47]), .A0_f (new_AGEMA_signal_4229), .A1_t (new_AGEMA_signal_4230), .A1_f (new_AGEMA_signal_4231), .B0_t (Midori_rounds_SR_Inv_Result[7]), .B0_f (new_AGEMA_signal_5514), .B1_t (new_AGEMA_signal_5515), .B1_f (new_AGEMA_signal_5516), .Z0_t (Midori_rounds_mul_ResultXORkey[47]), .Z0_f (new_AGEMA_signal_5658), .Z1_t (new_AGEMA_signal_5659), .Z1_f (new_AGEMA_signal_5660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U59 ( .A0_t (Midori_rounds_SelectedKey[46]), .A0_f (new_AGEMA_signal_4226), .A1_t (new_AGEMA_signal_4227), .A1_f (new_AGEMA_signal_4228), .B0_t (Midori_rounds_SR_Inv_Result[6]), .B0_f (new_AGEMA_signal_5752), .B1_t (new_AGEMA_signal_5753), .B1_f (new_AGEMA_signal_5754), .Z0_t (Midori_rounds_mul_ResultXORkey[46]), .Z0_f (new_AGEMA_signal_5827), .Z1_t (new_AGEMA_signal_5828), .Z1_f (new_AGEMA_signal_5829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U58 ( .A0_t (Midori_rounds_SelectedKey[45]), .A0_f (new_AGEMA_signal_4223), .A1_t (new_AGEMA_signal_4224), .A1_f (new_AGEMA_signal_4225), .B0_t (Midori_rounds_SR_Inv_Result[5]), .B0_f (new_AGEMA_signal_5529), .B1_t (new_AGEMA_signal_5530), .B1_f (new_AGEMA_signal_5531), .Z0_t (Midori_rounds_mul_ResultXORkey[45]), .Z0_f (new_AGEMA_signal_5661), .Z1_t (new_AGEMA_signal_5662), .Z1_f (new_AGEMA_signal_5663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U57 ( .A0_t (Midori_rounds_SelectedKey[43]), .A0_f (new_AGEMA_signal_4217), .A1_t (new_AGEMA_signal_4218), .A1_f (new_AGEMA_signal_4219), .B0_t (Midori_rounds_SR_Inv_Result[47]), .B0_f (new_AGEMA_signal_5517), .B1_t (new_AGEMA_signal_5518), .B1_f (new_AGEMA_signal_5519), .Z0_t (Midori_rounds_mul_ResultXORkey[43]), .Z0_f (new_AGEMA_signal_5664), .Z1_t (new_AGEMA_signal_5665), .Z1_f (new_AGEMA_signal_5666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U56 ( .A0_t (Midori_rounds_SelectedKey[42]), .A0_f (new_AGEMA_signal_4214), .A1_t (new_AGEMA_signal_4215), .A1_f (new_AGEMA_signal_4216), .B0_t (Midori_rounds_SR_Inv_Result[46]), .B0_f (new_AGEMA_signal_5755), .B1_t (new_AGEMA_signal_5756), .B1_f (new_AGEMA_signal_5757), .Z0_t (Midori_rounds_mul_ResultXORkey[42]), .Z0_f (new_AGEMA_signal_5830), .Z1_t (new_AGEMA_signal_5831), .Z1_f (new_AGEMA_signal_5832) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U55 ( .A0_t (Midori_rounds_SelectedKey[41]), .A0_f (new_AGEMA_signal_4211), .A1_t (new_AGEMA_signal_4212), .A1_f (new_AGEMA_signal_4213), .B0_t (Midori_rounds_SR_Inv_Result[45]), .B0_f (new_AGEMA_signal_5532), .B1_t (new_AGEMA_signal_5533), .B1_f (new_AGEMA_signal_5534), .Z0_t (Midori_rounds_mul_ResultXORkey[41]), .Z0_f (new_AGEMA_signal_5667), .Z1_t (new_AGEMA_signal_5668), .Z1_f (new_AGEMA_signal_5669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U54 ( .A0_t (Midori_rounds_SelectedKey[39]), .A0_f (new_AGEMA_signal_4205), .A1_t (new_AGEMA_signal_4206), .A1_f (new_AGEMA_signal_4207), .B0_t (Midori_rounds_SR_Inv_Result[19]), .B0_f (new_AGEMA_signal_5523), .B1_t (new_AGEMA_signal_5524), .B1_f (new_AGEMA_signal_5525), .Z0_t (Midori_rounds_mul_ResultXORkey[39]), .Z0_f (new_AGEMA_signal_5670), .Z1_t (new_AGEMA_signal_5671), .Z1_f (new_AGEMA_signal_5672) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U53 ( .A0_t (Midori_rounds_SelectedKey[38]), .A0_f (new_AGEMA_signal_4202), .A1_t (new_AGEMA_signal_4203), .A1_f (new_AGEMA_signal_4204), .B0_t (Midori_rounds_SR_Inv_Result[18]), .B0_f (new_AGEMA_signal_5758), .B1_t (new_AGEMA_signal_5759), .B1_f (new_AGEMA_signal_5760), .Z0_t (Midori_rounds_mul_ResultXORkey[38]), .Z0_f (new_AGEMA_signal_5833), .Z1_t (new_AGEMA_signal_5834), .Z1_f (new_AGEMA_signal_5835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U52 ( .A0_t (Midori_rounds_SelectedKey[37]), .A0_f (new_AGEMA_signal_4199), .A1_t (new_AGEMA_signal_4200), .A1_f (new_AGEMA_signal_4201), .B0_t (Midori_rounds_SR_Inv_Result[17]), .B0_f (new_AGEMA_signal_5538), .B1_t (new_AGEMA_signal_5539), .B1_f (new_AGEMA_signal_5540), .Z0_t (Midori_rounds_mul_ResultXORkey[37]), .Z0_f (new_AGEMA_signal_5673), .Z1_t (new_AGEMA_signal_5674), .Z1_f (new_AGEMA_signal_5675) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U51 ( .A0_t (Midori_rounds_SelectedKey[35]), .A0_f (new_AGEMA_signal_4193), .A1_t (new_AGEMA_signal_4194), .A1_f (new_AGEMA_signal_4195), .B0_t (Midori_rounds_SR_Inv_Result[59]), .B0_f (new_AGEMA_signal_5526), .B1_t (new_AGEMA_signal_5527), .B1_f (new_AGEMA_signal_5528), .Z0_t (Midori_rounds_mul_ResultXORkey[35]), .Z0_f (new_AGEMA_signal_5676), .Z1_t (new_AGEMA_signal_5677), .Z1_f (new_AGEMA_signal_5678) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U50 ( .A0_t (Midori_rounds_SelectedKey[34]), .A0_f (new_AGEMA_signal_4190), .A1_t (new_AGEMA_signal_4191), .A1_f (new_AGEMA_signal_4192), .B0_t (Midori_rounds_SR_Inv_Result[58]), .B0_f (new_AGEMA_signal_5761), .B1_t (new_AGEMA_signal_5762), .B1_f (new_AGEMA_signal_5763), .Z0_t (Midori_rounds_mul_ResultXORkey[34]), .Z0_f (new_AGEMA_signal_5836), .Z1_t (new_AGEMA_signal_5837), .Z1_f (new_AGEMA_signal_5838) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U49 ( .A0_t (Midori_rounds_SelectedKey[33]), .A0_f (new_AGEMA_signal_4187), .A1_t (new_AGEMA_signal_4188), .A1_f (new_AGEMA_signal_4189), .B0_t (Midori_rounds_SR_Inv_Result[57]), .B0_f (new_AGEMA_signal_5541), .B1_t (new_AGEMA_signal_5542), .B1_f (new_AGEMA_signal_5543), .Z0_t (Midori_rounds_mul_ResultXORkey[33]), .Z0_f (new_AGEMA_signal_5679), .Z1_t (new_AGEMA_signal_5680), .Z1_f (new_AGEMA_signal_5681) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U48 ( .A0_t (Midori_rounds_SelectedKey[31]), .A0_f (new_AGEMA_signal_4181), .A1_t (new_AGEMA_signal_4182), .A1_f (new_AGEMA_signal_4183), .B0_t (Midori_rounds_SR_Inv_Result[27]), .B0_f (new_AGEMA_signal_5544), .B1_t (new_AGEMA_signal_5545), .B1_f (new_AGEMA_signal_5546), .Z0_t (Midori_rounds_mul_ResultXORkey[31]), .Z0_f (new_AGEMA_signal_5682), .Z1_t (new_AGEMA_signal_5683), .Z1_f (new_AGEMA_signal_5684) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U47 ( .A0_t (Midori_rounds_SelectedKey[30]), .A0_f (new_AGEMA_signal_4178), .A1_t (new_AGEMA_signal_4179), .A1_f (new_AGEMA_signal_4180), .B0_t (Midori_rounds_SR_Inv_Result[26]), .B0_f (new_AGEMA_signal_5764), .B1_t (new_AGEMA_signal_5765), .B1_f (new_AGEMA_signal_5766), .Z0_t (Midori_rounds_mul_ResultXORkey[30]), .Z0_f (new_AGEMA_signal_5839), .Z1_t (new_AGEMA_signal_5840), .Z1_f (new_AGEMA_signal_5841) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U46 ( .A0_t (Midori_rounds_SelectedKey[29]), .A0_f (new_AGEMA_signal_4175), .A1_t (new_AGEMA_signal_4176), .A1_f (new_AGEMA_signal_4177), .B0_t (Midori_rounds_SR_Inv_Result[25]), .B0_f (new_AGEMA_signal_5559), .B1_t (new_AGEMA_signal_5560), .B1_f (new_AGEMA_signal_5561), .Z0_t (Midori_rounds_mul_ResultXORkey[29]), .Z0_f (new_AGEMA_signal_5685), .Z1_t (new_AGEMA_signal_5686), .Z1_f (new_AGEMA_signal_5687) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U45 ( .A0_t (Midori_rounds_SelectedKey[27]), .A0_f (new_AGEMA_signal_4169), .A1_t (new_AGEMA_signal_4170), .A1_f (new_AGEMA_signal_4171), .B0_t (Midori_rounds_SR_Inv_Result[51]), .B0_f (new_AGEMA_signal_5547), .B1_t (new_AGEMA_signal_5548), .B1_f (new_AGEMA_signal_5549), .Z0_t (Midori_rounds_mul_ResultXORkey[27]), .Z0_f (new_AGEMA_signal_5688), .Z1_t (new_AGEMA_signal_5689), .Z1_f (new_AGEMA_signal_5690) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U44 ( .A0_t (Midori_rounds_SelectedKey[26]), .A0_f (new_AGEMA_signal_4166), .A1_t (new_AGEMA_signal_4167), .A1_f (new_AGEMA_signal_4168), .B0_t (Midori_rounds_SR_Inv_Result[50]), .B0_f (new_AGEMA_signal_5767), .B1_t (new_AGEMA_signal_5768), .B1_f (new_AGEMA_signal_5769), .Z0_t (Midori_rounds_mul_ResultXORkey[26]), .Z0_f (new_AGEMA_signal_5842), .Z1_t (new_AGEMA_signal_5843), .Z1_f (new_AGEMA_signal_5844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U43 ( .A0_t (Midori_rounds_SelectedKey[25]), .A0_f (new_AGEMA_signal_4163), .A1_t (new_AGEMA_signal_4164), .A1_f (new_AGEMA_signal_4165), .B0_t (Midori_rounds_SR_Inv_Result[49]), .B0_f (new_AGEMA_signal_5562), .B1_t (new_AGEMA_signal_5563), .B1_f (new_AGEMA_signal_5564), .Z0_t (Midori_rounds_mul_ResultXORkey[25]), .Z0_f (new_AGEMA_signal_5691), .Z1_t (new_AGEMA_signal_5692), .Z1_f (new_AGEMA_signal_5693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U42 ( .A0_t (Midori_rounds_SelectedKey[23]), .A0_f (new_AGEMA_signal_4157), .A1_t (new_AGEMA_signal_4158), .A1_f (new_AGEMA_signal_4159), .B0_t (Midori_rounds_SR_Inv_Result[15]), .B0_f (new_AGEMA_signal_5553), .B1_t (new_AGEMA_signal_5554), .B1_f (new_AGEMA_signal_5555), .Z0_t (Midori_rounds_mul_ResultXORkey[23]), .Z0_f (new_AGEMA_signal_5694), .Z1_t (new_AGEMA_signal_5695), .Z1_f (new_AGEMA_signal_5696) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U41 ( .A0_t (Midori_rounds_SelectedKey[22]), .A0_f (new_AGEMA_signal_4154), .A1_t (new_AGEMA_signal_4155), .A1_f (new_AGEMA_signal_4156), .B0_t (Midori_rounds_SR_Inv_Result[14]), .B0_f (new_AGEMA_signal_5770), .B1_t (new_AGEMA_signal_5771), .B1_f (new_AGEMA_signal_5772), .Z0_t (Midori_rounds_mul_ResultXORkey[22]), .Z0_f (new_AGEMA_signal_5845), .Z1_t (new_AGEMA_signal_5846), .Z1_f (new_AGEMA_signal_5847) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U40 ( .A0_t (Midori_rounds_SelectedKey[21]), .A0_f (new_AGEMA_signal_4151), .A1_t (new_AGEMA_signal_4152), .A1_f (new_AGEMA_signal_4153), .B0_t (Midori_rounds_SR_Inv_Result[13]), .B0_f (new_AGEMA_signal_5568), .B1_t (new_AGEMA_signal_5569), .B1_f (new_AGEMA_signal_5570), .Z0_t (Midori_rounds_mul_ResultXORkey[21]), .Z0_f (new_AGEMA_signal_5697), .Z1_t (new_AGEMA_signal_5698), .Z1_f (new_AGEMA_signal_5699) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U39 ( .A0_t (Midori_rounds_SelectedKey[19]), .A0_f (new_AGEMA_signal_4145), .A1_t (new_AGEMA_signal_4146), .A1_f (new_AGEMA_signal_4147), .B0_t (Midori_rounds_SR_Inv_Result[39]), .B0_f (new_AGEMA_signal_5556), .B1_t (new_AGEMA_signal_5557), .B1_f (new_AGEMA_signal_5558), .Z0_t (Midori_rounds_mul_ResultXORkey[19]), .Z0_f (new_AGEMA_signal_5700), .Z1_t (new_AGEMA_signal_5701), .Z1_f (new_AGEMA_signal_5702) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U38 ( .A0_t (Midori_rounds_SelectedKey[18]), .A0_f (new_AGEMA_signal_4142), .A1_t (new_AGEMA_signal_4143), .A1_f (new_AGEMA_signal_4144), .B0_t (Midori_rounds_SR_Inv_Result[38]), .B0_f (new_AGEMA_signal_5773), .B1_t (new_AGEMA_signal_5774), .B1_f (new_AGEMA_signal_5775), .Z0_t (Midori_rounds_mul_ResultXORkey[18]), .Z0_f (new_AGEMA_signal_5848), .Z1_t (new_AGEMA_signal_5849), .Z1_f (new_AGEMA_signal_5850) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U37 ( .A0_t (Midori_rounds_SelectedKey[17]), .A0_f (new_AGEMA_signal_4139), .A1_t (new_AGEMA_signal_4140), .A1_f (new_AGEMA_signal_4141), .B0_t (Midori_rounds_SR_Inv_Result[37]), .B0_f (new_AGEMA_signal_5571), .B1_t (new_AGEMA_signal_5572), .B1_f (new_AGEMA_signal_5573), .Z0_t (Midori_rounds_mul_ResultXORkey[17]), .Z0_f (new_AGEMA_signal_5703), .Z1_t (new_AGEMA_signal_5704), .Z1_f (new_AGEMA_signal_5705) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U36 ( .A0_t (Midori_rounds_SelectedKey[15]), .A0_f (new_AGEMA_signal_4133), .A1_t (new_AGEMA_signal_4134), .A1_f (new_AGEMA_signal_4135), .B0_t (Midori_rounds_SR_Inv_Result[35]), .B0_f (new_AGEMA_signal_5574), .B1_t (new_AGEMA_signal_5575), .B1_f (new_AGEMA_signal_5576), .Z0_t (Midori_rounds_mul_ResultXORkey[15]), .Z0_f (new_AGEMA_signal_5706), .Z1_t (new_AGEMA_signal_5707), .Z1_f (new_AGEMA_signal_5708) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U35 ( .A0_t (Midori_rounds_SelectedKey[14]), .A0_f (new_AGEMA_signal_4130), .A1_t (new_AGEMA_signal_4131), .A1_f (new_AGEMA_signal_4132), .B0_t (Midori_rounds_SR_Inv_Result[34]), .B0_f (new_AGEMA_signal_5776), .B1_t (new_AGEMA_signal_5777), .B1_f (new_AGEMA_signal_5778), .Z0_t (Midori_rounds_mul_ResultXORkey[14]), .Z0_f (new_AGEMA_signal_5851), .Z1_t (new_AGEMA_signal_5852), .Z1_f (new_AGEMA_signal_5853) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U34 ( .A0_t (Midori_rounds_SelectedKey[13]), .A0_f (new_AGEMA_signal_4127), .A1_t (new_AGEMA_signal_4128), .A1_f (new_AGEMA_signal_4129), .B0_t (Midori_rounds_SR_Inv_Result[33]), .B0_f (new_AGEMA_signal_5589), .B1_t (new_AGEMA_signal_5590), .B1_f (new_AGEMA_signal_5591), .Z0_t (Midori_rounds_mul_ResultXORkey[13]), .Z0_f (new_AGEMA_signal_5709), .Z1_t (new_AGEMA_signal_5710), .Z1_f (new_AGEMA_signal_5711) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U33 ( .A0_t (Midori_rounds_SelectedKey[11]), .A0_f (new_AGEMA_signal_4121), .A1_t (new_AGEMA_signal_4122), .A1_f (new_AGEMA_signal_4123), .B0_t (Midori_rounds_SR_Inv_Result[11]), .B0_f (new_AGEMA_signal_5577), .B1_t (new_AGEMA_signal_5578), .B1_f (new_AGEMA_signal_5579), .Z0_t (Midori_rounds_mul_ResultXORkey[11]), .Z0_f (new_AGEMA_signal_5712), .Z1_t (new_AGEMA_signal_5713), .Z1_f (new_AGEMA_signal_5714) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U32 ( .A0_t (Midori_rounds_SelectedKey[10]), .A0_f (new_AGEMA_signal_4118), .A1_t (new_AGEMA_signal_4119), .A1_f (new_AGEMA_signal_4120), .B0_t (Midori_rounds_SR_Inv_Result[10]), .B0_f (new_AGEMA_signal_5779), .B1_t (new_AGEMA_signal_5780), .B1_f (new_AGEMA_signal_5781), .Z0_t (Midori_rounds_mul_ResultXORkey[10]), .Z0_f (new_AGEMA_signal_5854), .Z1_t (new_AGEMA_signal_5855), .Z1_f (new_AGEMA_signal_5856) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U31 ( .A0_t (Midori_rounds_SelectedKey[9]), .A0_f (new_AGEMA_signal_4115), .A1_t (new_AGEMA_signal_4116), .A1_f (new_AGEMA_signal_4117), .B0_t (Midori_rounds_SR_Inv_Result[9]), .B0_f (new_AGEMA_signal_5592), .B1_t (new_AGEMA_signal_5593), .B1_f (new_AGEMA_signal_5594), .Z0_t (Midori_rounds_mul_ResultXORkey[9]), .Z0_f (new_AGEMA_signal_5715), .Z1_t (new_AGEMA_signal_5716), .Z1_f (new_AGEMA_signal_5717) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U30 ( .A0_t (Midori_rounds_SelectedKey[7]), .A0_f (new_AGEMA_signal_4109), .A1_t (new_AGEMA_signal_4110), .A1_f (new_AGEMA_signal_4111), .B0_t (Midori_rounds_SR_Inv_Result[55]), .B0_f (new_AGEMA_signal_5583), .B1_t (new_AGEMA_signal_5584), .B1_f (new_AGEMA_signal_5585), .Z0_t (Midori_rounds_mul_ResultXORkey[7]), .Z0_f (new_AGEMA_signal_5718), .Z1_t (new_AGEMA_signal_5719), .Z1_f (new_AGEMA_signal_5720) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U29 ( .A0_t (Midori_rounds_SelectedKey[6]), .A0_f (new_AGEMA_signal_4106), .A1_t (new_AGEMA_signal_4107), .A1_f (new_AGEMA_signal_4108), .B0_t (Midori_rounds_SR_Inv_Result[54]), .B0_f (new_AGEMA_signal_5782), .B1_t (new_AGEMA_signal_5783), .B1_f (new_AGEMA_signal_5784), .Z0_t (Midori_rounds_mul_ResultXORkey[6]), .Z0_f (new_AGEMA_signal_5857), .Z1_t (new_AGEMA_signal_5858), .Z1_f (new_AGEMA_signal_5859) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U28 ( .A0_t (Midori_rounds_SelectedKey[5]), .A0_f (new_AGEMA_signal_4103), .A1_t (new_AGEMA_signal_4104), .A1_f (new_AGEMA_signal_4105), .B0_t (Midori_rounds_SR_Inv_Result[53]), .B0_f (new_AGEMA_signal_5598), .B1_t (new_AGEMA_signal_5599), .B1_f (new_AGEMA_signal_5600), .Z0_t (Midori_rounds_mul_ResultXORkey[5]), .Z0_f (new_AGEMA_signal_5721), .Z1_t (new_AGEMA_signal_5722), .Z1_f (new_AGEMA_signal_5723) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U27 ( .A0_t (Midori_rounds_SelectedKey[3]), .A0_f (new_AGEMA_signal_4097), .A1_t (new_AGEMA_signal_4098), .A1_f (new_AGEMA_signal_4099), .B0_t (Midori_rounds_SR_Inv_Result[31]), .B0_f (new_AGEMA_signal_5586), .B1_t (new_AGEMA_signal_5587), .B1_f (new_AGEMA_signal_5588), .Z0_t (Midori_rounds_mul_ResultXORkey[3]), .Z0_f (new_AGEMA_signal_5724), .Z1_t (new_AGEMA_signal_5725), .Z1_f (new_AGEMA_signal_5726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U26 ( .A0_t (Midori_rounds_SelectedKey[2]), .A0_f (new_AGEMA_signal_4094), .A1_t (new_AGEMA_signal_4095), .A1_f (new_AGEMA_signal_4096), .B0_t (Midori_rounds_SR_Inv_Result[30]), .B0_f (new_AGEMA_signal_5785), .B1_t (new_AGEMA_signal_5786), .B1_f (new_AGEMA_signal_5787), .Z0_t (Midori_rounds_mul_ResultXORkey[2]), .Z0_f (new_AGEMA_signal_5860), .Z1_t (new_AGEMA_signal_5861), .Z1_f (new_AGEMA_signal_5862) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U25 ( .A0_t (Midori_rounds_SelectedKey[1]), .A0_f (new_AGEMA_signal_4091), .A1_t (new_AGEMA_signal_4092), .A1_f (new_AGEMA_signal_4093), .B0_t (Midori_rounds_SR_Inv_Result[29]), .B0_f (new_AGEMA_signal_5601), .B1_t (new_AGEMA_signal_5602), .B1_f (new_AGEMA_signal_5603), .Z0_t (Midori_rounds_mul_ResultXORkey[1]), .Z0_f (new_AGEMA_signal_5727), .Z1_t (new_AGEMA_signal_5728), .Z1_f (new_AGEMA_signal_5729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U24 ( .A0_t (Midori_rounds_SelectedKey[43]), .A0_f (new_AGEMA_signal_4217), .A1_t (new_AGEMA_signal_4218), .A1_f (new_AGEMA_signal_4219), .B0_t (Midori_rounds_SR_Result[55]), .B0_f (new_AGEMA_signal_4406), .B1_t (new_AGEMA_signal_4407), .B1_f (new_AGEMA_signal_4408), .Z0_t (Midori_rounds_sub_ResultXORkey[43]), .Z0_f (new_AGEMA_signal_4618), .Z1_t (new_AGEMA_signal_4619), .Z1_f (new_AGEMA_signal_4620) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U23 ( .A0_t (Midori_rounds_SelectedKey[41]), .A0_f (new_AGEMA_signal_4211), .A1_t (new_AGEMA_signal_4212), .A1_f (new_AGEMA_signal_4213), .B0_t (Midori_rounds_SR_Result[53]), .B0_f (new_AGEMA_signal_4409), .B1_t (new_AGEMA_signal_4410), .B1_f (new_AGEMA_signal_4411), .Z0_t (Midori_rounds_sub_ResultXORkey[41]), .Z0_f (new_AGEMA_signal_4621), .Z1_t (new_AGEMA_signal_4622), .Z1_f (new_AGEMA_signal_4623) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U22 ( .A0_t (Midori_rounds_SelectedKey[31]), .A0_f (new_AGEMA_signal_4181), .A1_t (new_AGEMA_signal_4182), .A1_f (new_AGEMA_signal_4183), .B0_t (Midori_rounds_SR_Result[3]), .B0_f (new_AGEMA_signal_4364), .B1_t (new_AGEMA_signal_4365), .B1_f (new_AGEMA_signal_4366), .Z0_t (Midori_rounds_sub_ResultXORkey[31]), .Z0_f (new_AGEMA_signal_4624), .Z1_t (new_AGEMA_signal_4625), .Z1_f (new_AGEMA_signal_4626) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U21 ( .A0_t (Midori_rounds_SelectedKey[29]), .A0_f (new_AGEMA_signal_4175), .A1_t (new_AGEMA_signal_4176), .A1_f (new_AGEMA_signal_4177), .B0_t (Midori_rounds_SR_Result[1]), .B0_f (new_AGEMA_signal_4367), .B1_t (new_AGEMA_signal_4368), .B1_f (new_AGEMA_signal_4369), .Z0_t (Midori_rounds_sub_ResultXORkey[29]), .Z0_f (new_AGEMA_signal_4627), .Z1_t (new_AGEMA_signal_4628), .Z1_f (new_AGEMA_signal_4629) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U20 ( .A0_t (Midori_rounds_SelectedKey[63]), .A0_f (new_AGEMA_signal_4277), .A1_t (new_AGEMA_signal_4278), .A1_f (new_AGEMA_signal_4279), .B0_t (Midori_rounds_SR_Result[63]), .B0_f (new_AGEMA_signal_4466), .B1_t (new_AGEMA_signal_4467), .B1_f (new_AGEMA_signal_4468), .Z0_t (Midori_rounds_sub_ResultXORkey[63]), .Z0_f (new_AGEMA_signal_4630), .Z1_t (new_AGEMA_signal_4631), .Z1_f (new_AGEMA_signal_4632) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U19 ( .A0_t (Midori_rounds_SelectedKey[61]), .A0_f (new_AGEMA_signal_4271), .A1_t (new_AGEMA_signal_4272), .A1_f (new_AGEMA_signal_4273), .B0_t (Midori_rounds_SR_Result[61]), .B0_f (new_AGEMA_signal_4469), .B1_t (new_AGEMA_signal_4470), .B1_f (new_AGEMA_signal_4471), .Z0_t (Midori_rounds_sub_ResultXORkey[61]), .Z0_f (new_AGEMA_signal_4633), .Z1_t (new_AGEMA_signal_4634), .Z1_f (new_AGEMA_signal_4635) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U18 ( .A0_t (Midori_rounds_SelectedKey[26]), .A0_f (new_AGEMA_signal_4166), .A1_t (new_AGEMA_signal_4167), .A1_f (new_AGEMA_signal_4168), .B0_t (Midori_rounds_SR_Result[30]), .B0_f (new_AGEMA_signal_4721), .B1_t (new_AGEMA_signal_4722), .B1_f (new_AGEMA_signal_4723), .Z0_t (Midori_rounds_sub_ResultXORkey[26]), .Z0_f (new_AGEMA_signal_4899), .Z1_t (new_AGEMA_signal_4900), .Z1_f (new_AGEMA_signal_4901) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U17 ( .A0_t (Midori_rounds_SelectedKey[62]), .A0_f (new_AGEMA_signal_4274), .A1_t (new_AGEMA_signal_4275), .A1_f (new_AGEMA_signal_4276), .B0_t (Midori_rounds_SR_Result[62]), .B0_f (new_AGEMA_signal_4775), .B1_t (new_AGEMA_signal_4776), .B1_f (new_AGEMA_signal_4777), .Z0_t (Midori_rounds_sub_ResultXORkey[62]), .Z0_f (new_AGEMA_signal_4902), .Z1_t (new_AGEMA_signal_4903), .Z1_f (new_AGEMA_signal_4904) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U16 ( .A0_t (Midori_rounds_SelectedKey[42]), .A0_f (new_AGEMA_signal_4214), .A1_t (new_AGEMA_signal_4215), .A1_f (new_AGEMA_signal_4216), .B0_t (Midori_rounds_SR_Result[54]), .B0_f (new_AGEMA_signal_4745), .B1_t (new_AGEMA_signal_4746), .B1_f (new_AGEMA_signal_4747), .Z0_t (Midori_rounds_sub_ResultXORkey[42]), .Z0_f (new_AGEMA_signal_4905), .Z1_t (new_AGEMA_signal_4906), .Z1_f (new_AGEMA_signal_4907) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U15 ( .A0_t (Midori_rounds_SelectedKey[59]), .A0_f (new_AGEMA_signal_4265), .A1_t (new_AGEMA_signal_4266), .A1_f (new_AGEMA_signal_4267), .B0_t (Midori_rounds_SR_Result[35]), .B0_f (new_AGEMA_signal_4448), .B1_t (new_AGEMA_signal_4449), .B1_f (new_AGEMA_signal_4450), .Z0_t (Midori_rounds_sub_ResultXORkey[59]), .Z0_f (new_AGEMA_signal_4636), .Z1_t (new_AGEMA_signal_4637), .Z1_f (new_AGEMA_signal_4638) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U14 ( .A0_t (Midori_rounds_SelectedKey[58]), .A0_f (new_AGEMA_signal_4262), .A1_t (new_AGEMA_signal_4263), .A1_f (new_AGEMA_signal_4264), .B0_t (Midori_rounds_SR_Result[34]), .B0_f (new_AGEMA_signal_4766), .B1_t (new_AGEMA_signal_4767), .B1_f (new_AGEMA_signal_4768), .Z0_t (Midori_rounds_sub_ResultXORkey[58]), .Z0_f (new_AGEMA_signal_4908), .Z1_t (new_AGEMA_signal_4909), .Z1_f (new_AGEMA_signal_4910) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U13 ( .A0_t (Midori_rounds_SelectedKey[57]), .A0_f (new_AGEMA_signal_4259), .A1_t (new_AGEMA_signal_4260), .A1_f (new_AGEMA_signal_4261), .B0_t (Midori_rounds_SR_Result[33]), .B0_f (new_AGEMA_signal_4451), .B1_t (new_AGEMA_signal_4452), .B1_f (new_AGEMA_signal_4453), .Z0_t (Midori_rounds_sub_ResultXORkey[57]), .Z0_f (new_AGEMA_signal_4639), .Z1_t (new_AGEMA_signal_4640), .Z1_f (new_AGEMA_signal_4641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U12 ( .A0_t (Midori_rounds_SelectedKey[47]), .A0_f (new_AGEMA_signal_4229), .A1_t (new_AGEMA_signal_4230), .A1_f (new_AGEMA_signal_4231), .B0_t (Midori_rounds_SR_Result[43]), .B0_f (new_AGEMA_signal_4418), .B1_t (new_AGEMA_signal_4419), .B1_f (new_AGEMA_signal_4420), .Z0_t (Midori_rounds_sub_ResultXORkey[47]), .Z0_f (new_AGEMA_signal_4642), .Z1_t (new_AGEMA_signal_4643), .Z1_f (new_AGEMA_signal_4644) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U11 ( .A0_t (Midori_rounds_SelectedKey[46]), .A0_f (new_AGEMA_signal_4226), .A1_t (new_AGEMA_signal_4227), .A1_f (new_AGEMA_signal_4228), .B0_t (Midori_rounds_SR_Result[42]), .B0_f (new_AGEMA_signal_4751), .B1_t (new_AGEMA_signal_4752), .B1_f (new_AGEMA_signal_4753), .Z0_t (Midori_rounds_sub_ResultXORkey[46]), .Z0_f (new_AGEMA_signal_4911), .Z1_t (new_AGEMA_signal_4912), .Z1_f (new_AGEMA_signal_4913) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U10 ( .A0_t (Midori_rounds_SelectedKey[45]), .A0_f (new_AGEMA_signal_4223), .A1_t (new_AGEMA_signal_4224), .A1_f (new_AGEMA_signal_4225), .B0_t (Midori_rounds_SR_Result[41]), .B0_f (new_AGEMA_signal_4421), .B1_t (new_AGEMA_signal_4422), .B1_f (new_AGEMA_signal_4423), .Z0_t (Midori_rounds_sub_ResultXORkey[45]), .Z0_f (new_AGEMA_signal_4645), .Z1_t (new_AGEMA_signal_4646), .Z1_f (new_AGEMA_signal_4647) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U9 ( .A0_t (Midori_rounds_SelectedKey[27]), .A0_f (new_AGEMA_signal_4169), .A1_t (new_AGEMA_signal_4170), .A1_f (new_AGEMA_signal_4171), .B0_t (Midori_rounds_SR_Result[31]), .B0_f (new_AGEMA_signal_4358), .B1_t (new_AGEMA_signal_4359), .B1_f (new_AGEMA_signal_4360), .Z0_t (Midori_rounds_sub_ResultXORkey[27]), .Z0_f (new_AGEMA_signal_4648), .Z1_t (new_AGEMA_signal_4649), .Z1_f (new_AGEMA_signal_4650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U8 ( .A0_t (Midori_rounds_SelectedKey[30]), .A0_f (new_AGEMA_signal_4178), .A1_t (new_AGEMA_signal_4179), .A1_f (new_AGEMA_signal_4180), .B0_t (Midori_rounds_SR_Result[2]), .B0_f (new_AGEMA_signal_4724), .B1_t (new_AGEMA_signal_4725), .B1_f (new_AGEMA_signal_4726), .Z0_t (Midori_rounds_sub_ResultXORkey[30]), .Z0_f (new_AGEMA_signal_4914), .Z1_t (new_AGEMA_signal_4915), .Z1_f (new_AGEMA_signal_4916) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U7 ( .A0_t (Midori_rounds_SelectedKey[25]), .A0_f (new_AGEMA_signal_4163), .A1_t (new_AGEMA_signal_4164), .A1_f (new_AGEMA_signal_4165), .B0_t (Midori_rounds_SR_Result[29]), .B0_f (new_AGEMA_signal_4361), .B1_t (new_AGEMA_signal_4362), .B1_f (new_AGEMA_signal_4363), .Z0_t (Midori_rounds_sub_ResultXORkey[25]), .Z0_f (new_AGEMA_signal_4651), .Z1_t (new_AGEMA_signal_4652), .Z1_f (new_AGEMA_signal_4653) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U6 ( .A0_t (Midori_rounds_SelectedKey[11]), .A0_f (new_AGEMA_signal_4121), .A1_t (new_AGEMA_signal_4122), .A1_f (new_AGEMA_signal_4123), .B0_t (Midori_rounds_SR_Result[11]), .B0_f (new_AGEMA_signal_4310), .B1_t (new_AGEMA_signal_4311), .B1_f (new_AGEMA_signal_4312), .Z0_t (Midori_rounds_sub_ResultXORkey[11]), .Z0_f (new_AGEMA_signal_4654), .Z1_t (new_AGEMA_signal_4655), .Z1_f (new_AGEMA_signal_4656) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U5 ( .A0_t (Midori_rounds_SelectedKey[10]), .A0_f (new_AGEMA_signal_4118), .A1_t (new_AGEMA_signal_4119), .A1_f (new_AGEMA_signal_4120), .B0_t (Midori_rounds_SR_Result[10]), .B0_f (new_AGEMA_signal_4697), .B1_t (new_AGEMA_signal_4698), .B1_f (new_AGEMA_signal_4699), .Z0_t (Midori_rounds_sub_ResultXORkey[10]), .Z0_f (new_AGEMA_signal_4917), .Z1_t (new_AGEMA_signal_4918), .Z1_f (new_AGEMA_signal_4919) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U4 ( .A0_t (Midori_rounds_SelectedKey[9]), .A0_f (new_AGEMA_signal_4115), .A1_t (new_AGEMA_signal_4116), .A1_f (new_AGEMA_signal_4117), .B0_t (Midori_rounds_SR_Result[9]), .B0_f (new_AGEMA_signal_4313), .B1_t (new_AGEMA_signal_4314), .B1_f (new_AGEMA_signal_4315), .Z0_t (Midori_rounds_sub_ResultXORkey[9]), .Z0_f (new_AGEMA_signal_4657), .Z1_t (new_AGEMA_signal_4658), .Z1_f (new_AGEMA_signal_4659) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U3 ( .A0_t (Midori_rounds_SelectedKey[15]), .A0_f (new_AGEMA_signal_4133), .A1_t (new_AGEMA_signal_4134), .A1_f (new_AGEMA_signal_4135), .B0_t (Midori_rounds_SR_Result[23]), .B0_f (new_AGEMA_signal_4322), .B1_t (new_AGEMA_signal_4323), .B1_f (new_AGEMA_signal_4324), .Z0_t (Midori_rounds_sub_ResultXORkey[15]), .Z0_f (new_AGEMA_signal_4660), .Z1_t (new_AGEMA_signal_4661), .Z1_f (new_AGEMA_signal_4662) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U2 ( .A0_t (Midori_rounds_SelectedKey[14]), .A0_f (new_AGEMA_signal_4130), .A1_t (new_AGEMA_signal_4131), .A1_f (new_AGEMA_signal_4132), .B0_t (Midori_rounds_SR_Result[22]), .B0_f (new_AGEMA_signal_4703), .B1_t (new_AGEMA_signal_4704), .B1_f (new_AGEMA_signal_4705), .Z0_t (Midori_rounds_sub_ResultXORkey[14]), .Z0_f (new_AGEMA_signal_4920), .Z1_t (new_AGEMA_signal_4921), .Z1_f (new_AGEMA_signal_4922) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U1 ( .A0_t (Midori_rounds_SelectedKey[13]), .A0_f (new_AGEMA_signal_4127), .A1_t (new_AGEMA_signal_4128), .A1_f (new_AGEMA_signal_4129), .B0_t (Midori_rounds_SR_Result[21]), .B0_f (new_AGEMA_signal_4325), .B1_t (new_AGEMA_signal_4326), .B1_f (new_AGEMA_signal_4327), .Z0_t (Midori_rounds_sub_ResultXORkey[13]), .Z0_f (new_AGEMA_signal_4663), .Z1_t (new_AGEMA_signal_4664), .Z1_f (new_AGEMA_signal_4665) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U134 ( .A0_t (Midori_rounds_constant_MUX_n139), .A0_f (new_AGEMA_signal_5359), .B0_t (Midori_rounds_constant_MUX_n138), .B0_f (new_AGEMA_signal_5032), .Z0_t (Midori_rounds_round_Constant[3]), .Z0_f (new_AGEMA_signal_5473) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U133 ( .A0_t (Midori_rounds_constant_MUX_n137), .A0_f (new_AGEMA_signal_4671), .B0_t (Midori_rounds_constant_MUX_n136), .B0_f (new_AGEMA_signal_4928), .Z0_t (Midori_rounds_constant_MUX_n138), .Z0_f (new_AGEMA_signal_5032) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U132 ( .A0_t (Midori_rounds_constant_MUX_n103), .A0_f (new_AGEMA_signal_4679), .B0_t (Midori_rounds_constant_MUX_n134), .B0_f (new_AGEMA_signal_5351), .Z0_t (Midori_rounds_round_Constant[9]), .Z0_f (new_AGEMA_signal_5474) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U131 ( .A0_t (Midori_rounds_constant_MUX_n133), .A0_f (new_AGEMA_signal_5198), .B0_t (Midori_rounds_constant_MUX_n132), .B0_f (new_AGEMA_signal_5191), .Z0_t (Midori_rounds_constant_MUX_n134), .Z0_f (new_AGEMA_signal_5351) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U130 ( .A0_t (Midori_rounds_constant_MUX_n131), .A0_f (new_AGEMA_signal_4672), .B0_t (Midori_rounds_constant_MUX_n130), .B0_f (new_AGEMA_signal_5042), .Z0_t (Midori_rounds_constant_MUX_n132), .Z0_f (new_AGEMA_signal_5191) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U129 ( .A0_t (Midori_rounds_constant_MUX_n129), .A0_f (new_AGEMA_signal_4923), .B0_t (Midori_rounds_constant_MUX_n128), .B0_f (new_AGEMA_signal_4666), .Z0_t (Midori_rounds_round_Constant[11]), .Z0_f (new_AGEMA_signal_5033) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U128 ( .A0_t (Midori_rounds_constant_MUX_n125), .A0_f (new_AGEMA_signal_4075), .B0_t (Midori_rounds_constant_MUX_n126), .B0_f (new_AGEMA_signal_4062), .Z0_t (Midori_rounds_constant_MUX_n128), .Z0_f (new_AGEMA_signal_4666) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U126 ( .A0_t (Midori_rounds_constant_MUX_n124), .A0_f (new_AGEMA_signal_4667), .B0_t (Midori_rounds_constant_MUX_n123), .B0_f (new_AGEMA_signal_3613), .Z0_t (Midori_rounds_constant_MUX_n129), .Z0_f (new_AGEMA_signal_4923) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U125 ( .A0_t (Midori_rounds_constant_MUX_n122), .A0_f (new_AGEMA_signal_4060), .B0_t (Midori_rounds_constant_MUX_n120), .B0_f (new_AGEMA_signal_4084), .Z0_t (Midori_rounds_constant_MUX_n124), .Z0_f (new_AGEMA_signal_4667) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U124 ( .A0_t (Midori_rounds_constant_MUX_n119), .A0_f (new_AGEMA_signal_2597), .B0_t (Midori_rounds_constant_MUX_n118), .B0_f (new_AGEMA_signal_3614), .Z0_t (Midori_rounds_constant_MUX_n122), .Z0_f (new_AGEMA_signal_4060) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U123 ( .A0_t (Midori_rounds_constant_MUX_n117), .A0_f (new_AGEMA_signal_5480), .B0_t (Midori_rounds_constant_MUX_n116), .B0_f (new_AGEMA_signal_5034), .Z0_t (Midori_rounds_round_Constant[12]), .Z0_f (new_AGEMA_signal_5730) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U122 ( .A0_t (Midori_rounds_constant_MUX_n115), .A0_f (new_AGEMA_signal_4674), .B0_t (Midori_rounds_constant_MUX_n114), .B0_f (new_AGEMA_signal_4927), .Z0_t (Midori_rounds_constant_MUX_n116), .Z0_f (new_AGEMA_signal_5034) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U121 ( .A0_t (Midori_rounds_constant_MUX_n113), .A0_f (new_AGEMA_signal_5352), .B0_t (Midori_rounds_constant_MUX_n110), .B0_f (new_AGEMA_signal_5192), .Z0_t (Midori_rounds_round_Constant[7]), .Z0_f (new_AGEMA_signal_5475) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U120 ( .A0_t (Midori_rounds_constant_MUX_n109), .A0_f (new_AGEMA_signal_4677), .B0_t (Midori_rounds_constant_MUX_n108), .B0_f (new_AGEMA_signal_5036), .Z0_t (Midori_rounds_constant_MUX_n110), .Z0_f (new_AGEMA_signal_5192) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U118 ( .A0_t (Midori_rounds_constant_MUX_n133), .A0_f (new_AGEMA_signal_5198), .B0_t (Midori_rounds_constant_MUX_n115), .B0_f (new_AGEMA_signal_4674), .Z0_t (Midori_rounds_constant_MUX_n113), .Z0_f (new_AGEMA_signal_5352) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U117 ( .A0_t (Midori_rounds_constant_MUX_n103), .A0_f (new_AGEMA_signal_4679), .B0_t (Midori_rounds_constant_MUX_n107), .B0_f (new_AGEMA_signal_5193), .Z0_t (Midori_rounds_round_Constant[15]), .Z0_f (new_AGEMA_signal_5353) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U116 ( .A0_t (Midori_rounds_constant_MUX_n136), .A0_f (new_AGEMA_signal_4928), .B0_t (Midori_rounds_constant_MUX_n106), .B0_f (new_AGEMA_signal_5035), .Z0_t (Midori_rounds_constant_MUX_n107), .Z0_f (new_AGEMA_signal_5193) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U115 ( .A0_t (Midori_rounds_constant_MUX_n83), .A0_f (new_AGEMA_signal_4678), .B0_t (Midori_rounds_constant_MUX_n104), .B0_f (new_AGEMA_signal_4932), .Z0_t (Midori_rounds_constant_MUX_n106), .Z0_f (new_AGEMA_signal_5035) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U113 ( .A0_t (Midori_rounds_constant_MUX_n102), .A0_f (new_AGEMA_signal_5194), .B0_t (Midori_rounds_constant_MUX_n130), .B0_f (new_AGEMA_signal_5042), .Z0_t (Midori_rounds_round_Constant[14]), .Z0_f (new_AGEMA_signal_5354) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U112 ( .A0_t (Midori_rounds_constant_MUX_n101), .A0_f (new_AGEMA_signal_5043), .B0_t (Midori_rounds_constant_MUX_n108), .B0_f (new_AGEMA_signal_5036), .Z0_t (Midori_rounds_constant_MUX_n102), .Z0_f (new_AGEMA_signal_5194) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U111 ( .A0_t (Midori_rounds_constant_MUX_n100), .A0_f (new_AGEMA_signal_4929), .B0_t (Midori_rounds_constant_MUX_n99), .B0_f (new_AGEMA_signal_4924), .Z0_t (Midori_rounds_constant_MUX_n108), .Z0_f (new_AGEMA_signal_5036) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U110 ( .A0_t (Midori_rounds_constant_MUX_n103), .A0_f (new_AGEMA_signal_4679), .B0_t (Midori_rounds_constant_MUX_n137), .B0_f (new_AGEMA_signal_4671), .Z0_t (Midori_rounds_constant_MUX_n99), .Z0_f (new_AGEMA_signal_4924) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U109 ( .A0_t (Midori_rounds_constant_MUX_n98), .A0_f (new_AGEMA_signal_5195), .B0_t (Midori_rounds_constant_MUX_n97), .B0_f (new_AGEMA_signal_4072), .Z0_t (Midori_rounds_round_Constant[10]), .Z0_f (new_AGEMA_signal_5355) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U108 ( .A0_t (Midori_rounds_constant_MUX_n96), .A0_f (new_AGEMA_signal_4074), .B0_t (Midori_rounds_constant_MUX_n95), .B0_f (new_AGEMA_signal_5037), .Z0_t (Midori_rounds_constant_MUX_n98), .Z0_f (new_AGEMA_signal_5195) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U107 ( .A0_t (round_Signal[0]), .A0_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_constant_MUX_n94), .B0_f (new_AGEMA_signal_4925), .Z0_t (Midori_rounds_constant_MUX_n95), .Z0_f (new_AGEMA_signal_5037) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U106 ( .A0_t (Midori_rounds_constant_MUX_n93), .A0_f (new_AGEMA_signal_3621), .B0_t (Midori_rounds_constant_MUX_n92), .B0_f (new_AGEMA_signal_4668), .Z0_t (Midori_rounds_constant_MUX_n94), .Z0_f (new_AGEMA_signal_4925) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U105 ( .A0_t (Midori_rounds_constant_MUX_n118), .A0_f (new_AGEMA_signal_3614), .B0_t (Midori_rounds_constant_MUX_n91), .B0_f (new_AGEMA_signal_4061), .Z0_t (Midori_rounds_constant_MUX_n92), .Z0_f (new_AGEMA_signal_4668) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U104 ( .A0_t (enc_dec_t), .A0_f (enc_dec_f), .B0_t (Midori_rounds_constant_MUX_n123), .B0_f (new_AGEMA_signal_3613), .Z0_t (Midori_rounds_constant_MUX_n91), .Z0_f (new_AGEMA_signal_4061) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U103 ( .A0_t (Midori_rounds_constant_MUX_n35), .A0_f (new_AGEMA_signal_2592), .B0_t (Midori_rounds_constant_MUX_n88), .B0_f (new_AGEMA_signal_2595), .Z0_t (Midori_rounds_constant_MUX_n123), .Z0_f (new_AGEMA_signal_3613) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U102 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (Midori_rounds_constant_MUX_n86), .B0_f (new_AGEMA_signal_2596), .Z0_t (Midori_rounds_constant_MUX_n118), .Z0_f (new_AGEMA_signal_3614) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U101 ( .A0_t (Midori_rounds_constant_MUX_n85), .A0_f (new_AGEMA_signal_5038), .B0_t (Midori_rounds_constant_MUX_n125), .B0_f (new_AGEMA_signal_4075), .Z0_t (Midori_rounds_round_Constant[6]), .Z0_f (new_AGEMA_signal_5196) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U100 ( .A0_t (Midori_rounds_constant_MUX_n114), .A0_f (new_AGEMA_signal_4927), .B0_t (Midori_rounds_constant_MUX_n84), .B0_f (new_AGEMA_signal_4926), .Z0_t (Midori_rounds_constant_MUX_n85), .Z0_f (new_AGEMA_signal_5038) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U99 ( .A0_t (Midori_rounds_constant_MUX_n83), .A0_f (new_AGEMA_signal_4678), .B0_t (Midori_rounds_constant_MUX_n131), .B0_f (new_AGEMA_signal_4672), .Z0_t (Midori_rounds_constant_MUX_n84), .Z0_f (new_AGEMA_signal_4926) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U97 ( .A0_t (Midori_rounds_constant_MUX_n82), .A0_f (new_AGEMA_signal_4670), .B0_t (Midori_rounds_constant_MUX_n81), .B0_f (new_AGEMA_signal_4673), .Z0_t (Midori_rounds_constant_MUX_n114), .Z0_f (new_AGEMA_signal_4927) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U96 ( .A0_t (Midori_rounds_constant_MUX_n80), .A0_f (new_AGEMA_signal_5200), .B0_t (Midori_rounds_constant_MUX_n79), .B0_f (new_AGEMA_signal_5039), .Z0_t (Midori_rounds_round_Constant[5]), .Z0_f (new_AGEMA_signal_5356) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U95 ( .A0_t (Midori_rounds_constant_MUX_n137), .A0_f (new_AGEMA_signal_4671), .B0_t (Midori_rounds_constant_MUX_n78), .B0_f (new_AGEMA_signal_4930), .Z0_t (Midori_rounds_constant_MUX_n79), .Z0_f (new_AGEMA_signal_5039) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U94 ( .A0_t (Midori_rounds_constant_MUX_n77), .A0_f (new_AGEMA_signal_5731), .B0_t (Midori_rounds_constant_MUX_n76), .B0_f (new_AGEMA_signal_5041), .Z0_t (Midori_rounds_round_Constant[1]), .Z0_f (new_AGEMA_signal_5863) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U93 ( .A0_t (Midori_rounds_constant_MUX_n136), .A0_f (new_AGEMA_signal_4928), .B0_t (Midori_rounds_constant_MUX_n75), .B0_f (new_AGEMA_signal_5476), .Z0_t (Midori_rounds_constant_MUX_n77), .Z0_f (new_AGEMA_signal_5731) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U92 ( .A0_t (Midori_rounds_constant_MUX_n74), .A0_f (new_AGEMA_signal_5360), .B0_t (Midori_rounds_constant_MUX_n131), .B0_f (new_AGEMA_signal_4672), .Z0_t (Midori_rounds_constant_MUX_n75), .Z0_f (new_AGEMA_signal_5476) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U91 ( .A0_t (Midori_rounds_constant_MUX_n73), .A0_f (new_AGEMA_signal_4063), .B0_t (Midori_rounds_constant_MUX_n72), .B0_f (new_AGEMA_signal_4669), .Z0_t (Midori_rounds_constant_MUX_n136), .Z0_f (new_AGEMA_signal_4928) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U90 ( .A0_t (Midori_rounds_constant_MUX_n126), .A0_f (new_AGEMA_signal_4062), .B0_t (enc_dec_t), .B0_f (enc_dec_f), .Z0_t (Midori_rounds_constant_MUX_n72), .Z0_f (new_AGEMA_signal_4669) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U88 ( .A0_t (round_Signal[0]), .A0_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_constant_MUX_n70), .B0_f (new_AGEMA_signal_3619), .Z0_t (Midori_rounds_constant_MUX_n126), .Z0_f (new_AGEMA_signal_4062) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U87 ( .A0_t (Midori_rounds_constant_MUX_n69), .A0_f (new_AGEMA_signal_2598), .B0_t (Midori_rounds_constant_MUX_n111), .B0_f (new_AGEMA_signal_3623), .Z0_t (Midori_rounds_constant_MUX_n73), .Z0_f (new_AGEMA_signal_4063) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U86 ( .A0_t (Midori_rounds_constant_MUX_n100), .A0_f (new_AGEMA_signal_4929), .B0_t (Midori_rounds_constant_MUX_n68), .B0_f (new_AGEMA_signal_5357), .Z0_t (Midori_rounds_round_Constant[13]), .Z0_f (new_AGEMA_signal_5477) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U85 ( .A0_t (Midori_rounds_constant_MUX_n76), .A0_f (new_AGEMA_signal_5041), .B0_t (Midori_rounds_constant_MUX_n66), .B0_f (new_AGEMA_signal_5197), .Z0_t (Midori_rounds_constant_MUX_n68), .Z0_f (new_AGEMA_signal_5357) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U83 ( .A0_t (Midori_rounds_constant_MUX_n42), .A0_f (new_AGEMA_signal_4676), .B0_t (Midori_rounds_constant_MUX_n82), .B0_f (new_AGEMA_signal_4670), .Z0_t (Midori_rounds_constant_MUX_n100), .Z0_f (new_AGEMA_signal_4929) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U82 ( .A0_t (round_Signal[0]), .A0_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_constant_MUX_n64), .B0_f (new_AGEMA_signal_4064), .Z0_t (Midori_rounds_constant_MUX_n82), .Z0_f (new_AGEMA_signal_4670) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U81 ( .A0_t (Midori_rounds_constant_MUX_n70), .A0_f (new_AGEMA_signal_3619), .B0_t (Midori_rounds_constant_MUX_n62), .B0_f (new_AGEMA_signal_3615), .Z0_t (Midori_rounds_constant_MUX_n64), .Z0_f (new_AGEMA_signal_4064) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U80 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (Midori_rounds_constant_MUX_n69), .B0_f (new_AGEMA_signal_2598), .Z0_t (Midori_rounds_constant_MUX_n62), .Z0_f (new_AGEMA_signal_3615) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U79 ( .A0_t (Midori_rounds_constant_MUX_n117), .A0_f (new_AGEMA_signal_5480), .B0_t (Midori_rounds_constant_MUX_n61), .B0_f (new_AGEMA_signal_5358), .Z0_t (Midori_rounds_round_Constant[4]), .Z0_f (new_AGEMA_signal_5732) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U78 ( .A0_t (Midori_rounds_constant_MUX_n137), .A0_f (new_AGEMA_signal_4671), .B0_t (Midori_rounds_constant_MUX_n66), .B0_f (new_AGEMA_signal_5197), .Z0_t (Midori_rounds_constant_MUX_n61), .Z0_f (new_AGEMA_signal_5358) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U77 ( .A0_t (Midori_rounds_constant_MUX_n60), .A0_f (new_AGEMA_signal_4675), .B0_t (Midori_rounds_constant_MUX_n130), .B0_f (new_AGEMA_signal_5042), .Z0_t (Midori_rounds_constant_MUX_n66), .Z0_f (new_AGEMA_signal_5197) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U76 ( .A0_t (Midori_rounds_constant_MUX_n59), .A0_f (new_AGEMA_signal_4066), .B0_t (Midori_rounds_constant_MUX_n58), .B0_f (new_AGEMA_signal_4065), .Z0_t (Midori_rounds_constant_MUX_n137), .Z0_f (new_AGEMA_signal_4671) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U75 ( .A0_t (Midori_rounds_constant_MUX_n88), .A0_f (new_AGEMA_signal_2595), .B0_t (Midori_rounds_constant_MUX_n121), .B0_f (new_AGEMA_signal_3616), .Z0_t (Midori_rounds_constant_MUX_n58), .Z0_f (new_AGEMA_signal_4065) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U74 ( .A0_t (Midori_rounds_constant_MUX_n57), .A0_f (new_AGEMA_signal_3620), .B0_t (Midori_rounds_constant_MUX_n56), .B0_f (new_AGEMA_signal_2600), .Z0_t (Midori_rounds_constant_MUX_n59), .Z0_f (new_AGEMA_signal_4066) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U73 ( .A0_t (Midori_rounds_constant_MUX_n55), .A0_f (new_AGEMA_signal_2594), .B0_t (round_Signal[2]), .B0_f (new_AGEMA_signal_2585), .Z0_t (Midori_rounds_constant_MUX_n121), .Z0_f (new_AGEMA_signal_3616) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U72 ( .A0_t (Midori_rounds_constant_MUX_n139), .A0_f (new_AGEMA_signal_5359), .B0_t (Midori_rounds_constant_MUX_n54), .B0_f (new_AGEMA_signal_5040), .Z0_t (Midori_rounds_round_Constant[2]), .Z0_f (new_AGEMA_signal_5478) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U71 ( .A0_t (Midori_rounds_constant_MUX_n42), .A0_f (new_AGEMA_signal_4676), .B0_t (Midori_rounds_constant_MUX_n78), .B0_f (new_AGEMA_signal_4930), .Z0_t (Midori_rounds_constant_MUX_n54), .Z0_f (new_AGEMA_signal_5040) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U70 ( .A0_t (Midori_rounds_constant_MUX_n60), .A0_f (new_AGEMA_signal_4675), .B0_t (Midori_rounds_constant_MUX_n131), .B0_f (new_AGEMA_signal_4672), .Z0_t (Midori_rounds_constant_MUX_n78), .Z0_f (new_AGEMA_signal_4930) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U69 ( .A0_t (Midori_rounds_constant_MUX_n53), .A0_f (new_AGEMA_signal_4068), .B0_t (Midori_rounds_constant_MUX_n52), .B0_f (new_AGEMA_signal_4067), .Z0_t (Midori_rounds_constant_MUX_n131), .Z0_f (new_AGEMA_signal_4672) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U68 ( .A0_t (Midori_rounds_constant_MUX_n119), .A0_f (new_AGEMA_signal_2597), .B0_t (Midori_rounds_constant_MUX_n51), .B0_f (new_AGEMA_signal_3617), .Z0_t (Midori_rounds_constant_MUX_n52), .Z0_f (new_AGEMA_signal_4067) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U67 ( .A0_t (Midori_rounds_constant_MUX_n88), .A0_f (new_AGEMA_signal_2595), .B0_t (Midori_rounds_constant_MUX_n50), .B0_f (new_AGEMA_signal_3622), .Z0_t (Midori_rounds_constant_MUX_n53), .Z0_f (new_AGEMA_signal_4068) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U66 ( .A0_t (Midori_rounds_constant_MUX_n133), .A0_f (new_AGEMA_signal_5198), .B0_t (Midori_rounds_constant_MUX_n81), .B0_f (new_AGEMA_signal_4673), .Z0_t (Midori_rounds_constant_MUX_n139), .Z0_f (new_AGEMA_signal_5359) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U65 ( .A0_t (Midori_rounds_constant_MUX_n125), .A0_f (new_AGEMA_signal_4075), .B0_t (Midori_rounds_constant_MUX_n76), .B0_f (new_AGEMA_signal_5041), .Z0_t (Midori_rounds_constant_MUX_n133), .Z0_f (new_AGEMA_signal_5198) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U64 ( .A0_t (round_Signal[1]), .A0_f (new_AGEMA_signal_2581), .B0_t (Midori_rounds_constant_MUX_n112), .B0_f (new_AGEMA_signal_4935), .Z0_t (Midori_rounds_constant_MUX_n76), .Z0_f (new_AGEMA_signal_5041) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U63 ( .A0_t (Midori_rounds_constant_MUX_n104), .A0_f (new_AGEMA_signal_4932), .B0_t (Midori_rounds_constant_MUX_n74), .B0_f (new_AGEMA_signal_5360), .Z0_t (Midori_rounds_round_Constant[0]), .Z0_f (new_AGEMA_signal_5479) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U62 ( .A0_t (Midori_rounds_constant_MUX_n109), .A0_f (new_AGEMA_signal_4677), .B0_t (Midori_rounds_constant_MUX_n49), .B0_f (new_AGEMA_signal_5199), .Z0_t (Midori_rounds_constant_MUX_n74), .Z0_f (new_AGEMA_signal_5360) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U61 ( .A0_t (Midori_rounds_constant_MUX_n48), .A0_f (new_AGEMA_signal_4931), .B0_t (Midori_rounds_constant_MUX_n130), .B0_f (new_AGEMA_signal_5042), .Z0_t (Midori_rounds_constant_MUX_n49), .Z0_f (new_AGEMA_signal_5199) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U60 ( .A0_t (round_Signal[1]), .A0_f (new_AGEMA_signal_2581), .B0_t (Midori_rounds_constant_MUX_n43), .B0_f (new_AGEMA_signal_4934), .Z0_t (Midori_rounds_constant_MUX_n130), .Z0_f (new_AGEMA_signal_5042) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U59 ( .A0_t (Midori_rounds_constant_MUX_n42), .A0_f (new_AGEMA_signal_4676), .B0_t (Midori_rounds_constant_MUX_n81), .B0_f (new_AGEMA_signal_4673), .Z0_t (Midori_rounds_constant_MUX_n48), .Z0_f (new_AGEMA_signal_4931) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U58 ( .A0_t (Midori_rounds_constant_MUX_n47), .A0_f (new_AGEMA_signal_4070), .B0_t (Midori_rounds_constant_MUX_n46), .B0_f (new_AGEMA_signal_4069), .Z0_t (Midori_rounds_constant_MUX_n81), .Z0_f (new_AGEMA_signal_4673) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U57 ( .A0_t (Midori_rounds_constant_MUX_n86), .A0_f (new_AGEMA_signal_2596), .B0_t (Midori_rounds_constant_MUX_n50), .B0_f (new_AGEMA_signal_3622), .Z0_t (Midori_rounds_constant_MUX_n46), .Z0_f (new_AGEMA_signal_4069) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U55 ( .A0_t (Midori_rounds_constant_MUX_n57), .A0_f (new_AGEMA_signal_3620), .B0_t (Midori_rounds_constant_MUX_n119), .B0_f (new_AGEMA_signal_2597), .Z0_t (Midori_rounds_constant_MUX_n47), .Z0_f (new_AGEMA_signal_4070) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U52 ( .A0_t (Midori_rounds_constant_MUX_n60), .A0_f (new_AGEMA_signal_4675), .B0_t (Midori_rounds_constant_MUX_n115), .B0_f (new_AGEMA_signal_4674), .Z0_t (Midori_rounds_constant_MUX_n104), .Z0_f (new_AGEMA_signal_4932) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U51 ( .A0_t (Midori_rounds_constant_MUX_n97), .A0_f (new_AGEMA_signal_4072), .B0_t (Midori_rounds_constant_MUX_n40), .B0_f (new_AGEMA_signal_4071), .Z0_t (Midori_rounds_constant_MUX_n115), .Z0_f (new_AGEMA_signal_4674) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U50 ( .A0_t (Midori_rounds_constant_MUX_n88), .A0_f (new_AGEMA_signal_2595), .B0_t (Midori_rounds_constant_MUX_n36), .B0_f (new_AGEMA_signal_3618), .Z0_t (Midori_rounds_constant_MUX_n40), .Z0_f (new_AGEMA_signal_4071) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U49 ( .A0_t (Midori_rounds_constant_MUX_n51), .A0_f (new_AGEMA_signal_3617), .B0_t (Midori_rounds_constant_MUX_n34), .B0_f (new_AGEMA_signal_2599), .Z0_t (Midori_rounds_constant_MUX_n97), .Z0_f (new_AGEMA_signal_4072) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U47 ( .A0_t (Midori_rounds_constant_MUX_n96), .A0_f (new_AGEMA_signal_4074), .B0_t (Midori_rounds_constant_MUX_n37), .B0_f (new_AGEMA_signal_4073), .Z0_t (Midori_rounds_constant_MUX_n60), .Z0_f (new_AGEMA_signal_4675) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U46 ( .A0_t (Midori_rounds_constant_MUX_n36), .A0_f (new_AGEMA_signal_3618), .B0_t (Midori_rounds_constant_MUX_n35), .B0_f (new_AGEMA_signal_2592), .Z0_t (Midori_rounds_constant_MUX_n37), .Z0_f (new_AGEMA_signal_4073) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U45 ( .A0_t (Midori_rounds_constant_MUX_n34), .A0_f (new_AGEMA_signal_2599), .B0_t (Midori_rounds_constant_MUX_n70), .B0_f (new_AGEMA_signal_3619), .Z0_t (Midori_rounds_constant_MUX_n96), .Z0_f (new_AGEMA_signal_4074) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U44 ( .A0_t (Midori_rounds_constant_MUX_n117), .A0_f (new_AGEMA_signal_5480), .B0_t (Midori_rounds_constant_MUX_n125), .B0_f (new_AGEMA_signal_4075), .Z0_t (Midori_rounds_round_Constant[8]), .Z0_f (new_AGEMA_signal_5733) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U43 ( .A0_t (round_Signal[0]), .A0_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_constant_MUX_n51), .B0_f (new_AGEMA_signal_3617), .Z0_t (Midori_rounds_constant_MUX_n125), .Z0_f (new_AGEMA_signal_4075) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U42 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (Midori_rounds_constant_MUX_n35), .B0_f (new_AGEMA_signal_2592), .Z0_t (Midori_rounds_constant_MUX_n51), .Z0_f (new_AGEMA_signal_3617) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U41 ( .A0_t (Midori_rounds_constant_MUX_n103), .A0_f (new_AGEMA_signal_4679), .B0_t (Midori_rounds_constant_MUX_n33), .B0_f (new_AGEMA_signal_5361), .Z0_t (Midori_rounds_constant_MUX_n117), .Z0_f (new_AGEMA_signal_5480) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U40 ( .A0_t (Midori_rounds_constant_MUX_n80), .A0_f (new_AGEMA_signal_5200), .B0_t (Midori_rounds_constant_MUX_n42), .B0_f (new_AGEMA_signal_4676), .Z0_t (Midori_rounds_constant_MUX_n33), .Z0_f (new_AGEMA_signal_5361) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U39 ( .A0_t (Midori_rounds_constant_MUX_n32), .A0_f (new_AGEMA_signal_4077), .B0_t (Midori_rounds_constant_MUX_n31), .B0_f (new_AGEMA_signal_4076), .Z0_t (Midori_rounds_constant_MUX_n42), .Z0_f (new_AGEMA_signal_4676) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U38 ( .A0_t (Midori_rounds_constant_MUX_n57), .A0_f (new_AGEMA_signal_3620), .B0_t (Midori_rounds_constant_MUX_n34), .B0_f (new_AGEMA_signal_2599), .Z0_t (Midori_rounds_constant_MUX_n31), .Z0_f (new_AGEMA_signal_4076) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U37 ( .A0_t (Midori_rounds_constant_MUX_n86), .A0_f (new_AGEMA_signal_2596), .B0_t (Midori_rounds_constant_MUX_n36), .B0_f (new_AGEMA_signal_3618), .Z0_t (Midori_rounds_constant_MUX_n32), .Z0_f (new_AGEMA_signal_4077) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U36 ( .A0_t (Midori_rounds_constant_MUX_n101), .A0_f (new_AGEMA_signal_5043), .B0_t (Midori_rounds_constant_MUX_n109), .B0_f (new_AGEMA_signal_4677), .Z0_t (Midori_rounds_constant_MUX_n80), .Z0_f (new_AGEMA_signal_5200) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U35 ( .A0_t (Midori_rounds_constant_MUX_n30), .A0_f (new_AGEMA_signal_4079), .B0_t (Midori_rounds_constant_MUX_n29), .B0_f (new_AGEMA_signal_4078), .Z0_t (Midori_rounds_constant_MUX_n109), .Z0_f (new_AGEMA_signal_4677) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U34 ( .A0_t (Midori_rounds_constant_MUX_n93), .A0_f (new_AGEMA_signal_3621), .B0_t (Midori_rounds_constant_MUX_n34), .B0_f (new_AGEMA_signal_2599), .Z0_t (Midori_rounds_constant_MUX_n29), .Z0_f (new_AGEMA_signal_4078) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U32 ( .A0_t (Midori_rounds_constant_MUX_n36), .A0_f (new_AGEMA_signal_3618), .B0_t (Midori_rounds_constant_MUX_n69), .B0_f (new_AGEMA_signal_2598), .Z0_t (Midori_rounds_constant_MUX_n30), .Z0_f (new_AGEMA_signal_4079) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U30 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (Midori_rounds_constant_MUX_n119), .B0_f (new_AGEMA_signal_2597), .Z0_t (Midori_rounds_constant_MUX_n36), .Z0_f (new_AGEMA_signal_3618) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U29 ( .A0_t (Midori_rounds_constant_MUX_n28), .A0_f (new_AGEMA_signal_4933), .B0_t (Midori_rounds_constant_MUX_n27), .B0_f (new_AGEMA_signal_4080), .Z0_t (Midori_rounds_constant_MUX_n101), .Z0_f (new_AGEMA_signal_5043) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U28 ( .A0_t (Midori_rounds_constant_MUX_n35), .A0_f (new_AGEMA_signal_2592), .B0_t (Midori_rounds_constant_MUX_n50), .B0_f (new_AGEMA_signal_3622), .Z0_t (Midori_rounds_constant_MUX_n27), .Z0_f (new_AGEMA_signal_4080) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U26 ( .A0_t (round_Signal[3]), .A0_f (new_AGEMA_signal_2584), .B0_t (round_Signal[1]), .B0_f (new_AGEMA_signal_2581), .Z0_t (Midori_rounds_constant_MUX_n35), .Z0_f (new_AGEMA_signal_2592) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U25 ( .A0_t (Midori_rounds_constant_MUX_n83), .A0_f (new_AGEMA_signal_4678), .B0_t (Midori_rounds_constant_MUX_n25), .B0_f (new_AGEMA_signal_4081), .Z0_t (Midori_rounds_constant_MUX_n28), .Z0_f (new_AGEMA_signal_4933) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U24 ( .A0_t (Midori_rounds_constant_MUX_n119), .A0_f (new_AGEMA_signal_2597), .B0_t (Midori_rounds_constant_MUX_n70), .B0_f (new_AGEMA_signal_3619), .Z0_t (Midori_rounds_constant_MUX_n25), .Z0_f (new_AGEMA_signal_4081) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U22 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (Midori_rounds_constant_MUX_n88), .B0_f (new_AGEMA_signal_2595), .Z0_t (Midori_rounds_constant_MUX_n70), .Z0_f (new_AGEMA_signal_3619) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U21 ( .A0_t (Midori_rounds_constant_MUX_n24), .A0_f (new_AGEMA_signal_4083), .B0_t (Midori_rounds_constant_MUX_n23), .B0_f (new_AGEMA_signal_4082), .Z0_t (Midori_rounds_constant_MUX_n83), .Z0_f (new_AGEMA_signal_4678) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U20 ( .A0_t (Midori_rounds_constant_MUX_n55), .A0_f (new_AGEMA_signal_2594), .B0_t (Midori_rounds_constant_MUX_n57), .B0_f (new_AGEMA_signal_3620), .Z0_t (Midori_rounds_constant_MUX_n23), .Z0_f (new_AGEMA_signal_4082) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U18 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (Midori_rounds_constant_MUX_n69), .B0_f (new_AGEMA_signal_2598), .Z0_t (Midori_rounds_constant_MUX_n57), .Z0_f (new_AGEMA_signal_3620) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U17 ( .A0_t (enc_dec_t), .A0_f (enc_dec_f), .B0_t (round_Signal[0]), .B0_f (new_AGEMA_signal_2582), .Z0_t (Midori_rounds_constant_MUX_n55), .Z0_f (new_AGEMA_signal_2594) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U16 ( .A0_t (Midori_rounds_constant_MUX_n111), .A0_f (new_AGEMA_signal_3623), .B0_t (Midori_rounds_constant_MUX_n88), .B0_f (new_AGEMA_signal_2595), .Z0_t (Midori_rounds_constant_MUX_n24), .Z0_f (new_AGEMA_signal_4083) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U15 ( .A0_t (round_Signal[1]), .A0_f (new_AGEMA_signal_2581), .B0_t (round_Signal[3]), .B0_f (new_AGEMA_signal_2584), .Z0_t (Midori_rounds_constant_MUX_n88), .Z0_f (new_AGEMA_signal_2595) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U13 ( .A0_t (Midori_rounds_constant_MUX_n22), .A0_f (new_AGEMA_signal_4085), .B0_t (Midori_rounds_constant_MUX_n120), .B0_f (new_AGEMA_signal_4084), .Z0_t (Midori_rounds_constant_MUX_n103), .Z0_f (new_AGEMA_signal_4679) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U12 ( .A0_t (Midori_rounds_constant_MUX_n119), .A0_f (new_AGEMA_signal_2597), .B0_t (Midori_rounds_constant_MUX_n93), .B0_f (new_AGEMA_signal_3621), .Z0_t (Midori_rounds_constant_MUX_n120), .Z0_f (new_AGEMA_signal_4084) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U11 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (Midori_rounds_constant_MUX_n86), .B0_f (new_AGEMA_signal_2596), .Z0_t (Midori_rounds_constant_MUX_n93), .Z0_f (new_AGEMA_signal_3621) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U10 ( .A0_t (round_Signal[3]), .A0_f (new_AGEMA_signal_2584), .B0_t (round_Signal[1]), .B0_f (new_AGEMA_signal_2581), .Z0_t (Midori_rounds_constant_MUX_n86), .Z0_f (new_AGEMA_signal_2596) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U8 ( .A0_t (round_Signal[0]), .A0_f (new_AGEMA_signal_2582), .B0_t (enc_dec_t), .B0_f (enc_dec_f), .Z0_t (Midori_rounds_constant_MUX_n119), .Z0_f (new_AGEMA_signal_2597) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U7 ( .A0_t (Midori_rounds_constant_MUX_n50), .A0_f (new_AGEMA_signal_3622), .B0_t (Midori_rounds_constant_MUX_n69), .B0_f (new_AGEMA_signal_2598), .Z0_t (Midori_rounds_constant_MUX_n22), .Z0_f (new_AGEMA_signal_4085) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U6 ( .A0_t (round_Signal[3]), .A0_f (new_AGEMA_signal_2584), .B0_t (round_Signal[1]), .B0_f (new_AGEMA_signal_2581), .Z0_t (Midori_rounds_constant_MUX_n69), .Z0_f (new_AGEMA_signal_2598) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U5 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (Midori_rounds_constant_MUX_n34), .B0_f (new_AGEMA_signal_2599), .Z0_t (Midori_rounds_constant_MUX_n50), .Z0_f (new_AGEMA_signal_3622) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U4 ( .A0_t (enc_dec_t), .A0_f (enc_dec_f), .B0_t (round_Signal[0]), .B0_f (new_AGEMA_signal_2582), .Z0_t (Midori_rounds_constant_MUX_n34), .Z0_f (new_AGEMA_signal_2599) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U2 ( .A0_t (round_Signal[2]), .A0_f (new_AGEMA_signal_2585), .B0_t (Midori_rounds_constant_MUX_n56), .B0_f (new_AGEMA_signal_2600), .Z0_t (Midori_rounds_constant_MUX_n111), .Z0_f (new_AGEMA_signal_3623) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U1 ( .A0_t (round_Signal[0]), .A0_f (new_AGEMA_signal_2582), .B0_t (enc_dec_t), .B0_f (enc_dec_f), .Z0_t (Midori_rounds_constant_MUX_n56), .Z0_f (new_AGEMA_signal_2600) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) Midori_rounds_constant_MUX_U53_XOR1_U1 ( .A0_t (Midori_rounds_constant_MUX_n121), .A0_f (new_AGEMA_signal_3616), .B0_t (Midori_rounds_constant_MUX_n111), .B0_f (new_AGEMA_signal_3623), .Z0_t (Midori_rounds_constant_MUX_U53_X), .Z0_f (new_AGEMA_signal_4086) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U53_AND1_U1 ( .A0_t (round_Signal[3]), .A0_f (new_AGEMA_signal_2584), .B0_t (Midori_rounds_constant_MUX_U53_X), .B0_f (new_AGEMA_signal_4086), .Z0_t (Midori_rounds_constant_MUX_U53_Y), .Z0_f (new_AGEMA_signal_4680) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) Midori_rounds_constant_MUX_U53_XOR2_U1 ( .A0_t (Midori_rounds_constant_MUX_U53_Y), .A0_f (new_AGEMA_signal_4680), .B0_t (Midori_rounds_constant_MUX_n121), .B0_f (new_AGEMA_signal_3616), .Z0_t (Midori_rounds_constant_MUX_n43), .Z0_f (new_AGEMA_signal_4934) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) Midori_rounds_constant_MUX_U119_XOR1_U1 ( .A0_t (Midori_rounds_constant_MUX_n111), .A0_f (new_AGEMA_signal_3623), .B0_t (Midori_rounds_constant_MUX_n121), .B0_f (new_AGEMA_signal_3616), .Z0_t (Midori_rounds_constant_MUX_U119_X), .Z0_f (new_AGEMA_signal_4087) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U119_AND1_U1 ( .A0_t (round_Signal[3]), .A0_f (new_AGEMA_signal_2584), .B0_t (Midori_rounds_constant_MUX_U119_X), .B0_f (new_AGEMA_signal_4087), .Z0_t (Midori_rounds_constant_MUX_U119_Y), .Z0_f (new_AGEMA_signal_4681) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) Midori_rounds_constant_MUX_U119_XOR2_U1 ( .A0_t (Midori_rounds_constant_MUX_U119_Y), .A0_f (new_AGEMA_signal_4681), .B0_t (Midori_rounds_constant_MUX_n111), .B0_f (new_AGEMA_signal_3623), .Z0_t (Midori_rounds_constant_MUX_n112), .Z0_f (new_AGEMA_signal_4935) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_0_U1_XOR1_U1 ( .A0_t (key_s0_t[64]), .A0_f (key_s0_f[64]), .A1_t (key_s1_t[64]), .A1_f (key_s1_f[64]), .B0_t (key_s0_t[0]), .B0_f (key_s0_f[0]), .B1_t (key_s1_t[0]), .B1_f (key_s1_f[0]), .Z0_t (Midori_rounds_MUXInst_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_2601), .Z1_t (new_AGEMA_signal_2602), .Z1_f (new_AGEMA_signal_2603) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_2601), .B1_t (new_AGEMA_signal_2602), .B1_f (new_AGEMA_signal_2603), .Z0_t (Midori_rounds_MUXInst_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_3624), .Z1_t (new_AGEMA_signal_3625), .Z1_f (new_AGEMA_signal_3626) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_0_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_3624), .A1_t (new_AGEMA_signal_3625), .A1_f (new_AGEMA_signal_3626), .B0_t (key_s0_t[64]), .B0_f (key_s0_f[64]), .B1_t (key_s1_t[64]), .B1_f (key_s1_f[64]), .Z0_t (Midori_rounds_SelectedKey[0]), .Z0_f (new_AGEMA_signal_4088), .Z1_t (new_AGEMA_signal_4089), .Z1_f (new_AGEMA_signal_4090) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_1_U1_XOR1_U1 ( .A0_t (key_s0_t[65]), .A0_f (key_s0_f[65]), .A1_t (key_s1_t[65]), .A1_f (key_s1_f[65]), .B0_t (key_s0_t[1]), .B0_f (key_s0_f[1]), .B1_t (key_s1_t[1]), .B1_f (key_s1_f[1]), .Z0_t (Midori_rounds_MUXInst_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_2604), .Z1_t (new_AGEMA_signal_2605), .Z1_f (new_AGEMA_signal_2606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_2604), .B1_t (new_AGEMA_signal_2605), .B1_f (new_AGEMA_signal_2606), .Z0_t (Midori_rounds_MUXInst_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_3627), .Z1_t (new_AGEMA_signal_3628), .Z1_f (new_AGEMA_signal_3629) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_1_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_3627), .A1_t (new_AGEMA_signal_3628), .A1_f (new_AGEMA_signal_3629), .B0_t (key_s0_t[65]), .B0_f (key_s0_f[65]), .B1_t (key_s1_t[65]), .B1_f (key_s1_f[65]), .Z0_t (Midori_rounds_SelectedKey[1]), .Z0_f (new_AGEMA_signal_4091), .Z1_t (new_AGEMA_signal_4092), .Z1_f (new_AGEMA_signal_4093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_2_U1_XOR1_U1 ( .A0_t (key_s0_t[66]), .A0_f (key_s0_f[66]), .A1_t (key_s1_t[66]), .A1_f (key_s1_f[66]), .B0_t (key_s0_t[2]), .B0_f (key_s0_f[2]), .B1_t (key_s1_t[2]), .B1_f (key_s1_f[2]), .Z0_t (Midori_rounds_MUXInst_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_2607), .Z1_t (new_AGEMA_signal_2608), .Z1_f (new_AGEMA_signal_2609) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_2607), .B1_t (new_AGEMA_signal_2608), .B1_f (new_AGEMA_signal_2609), .Z0_t (Midori_rounds_MUXInst_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_3630), .Z1_t (new_AGEMA_signal_3631), .Z1_f (new_AGEMA_signal_3632) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_2_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_3630), .A1_t (new_AGEMA_signal_3631), .A1_f (new_AGEMA_signal_3632), .B0_t (key_s0_t[66]), .B0_f (key_s0_f[66]), .B1_t (key_s1_t[66]), .B1_f (key_s1_f[66]), .Z0_t (Midori_rounds_SelectedKey[2]), .Z0_f (new_AGEMA_signal_4094), .Z1_t (new_AGEMA_signal_4095), .Z1_f (new_AGEMA_signal_4096) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_3_U1_XOR1_U1 ( .A0_t (key_s0_t[67]), .A0_f (key_s0_f[67]), .A1_t (key_s1_t[67]), .A1_f (key_s1_f[67]), .B0_t (key_s0_t[3]), .B0_f (key_s0_f[3]), .B1_t (key_s1_t[3]), .B1_f (key_s1_f[3]), .Z0_t (Midori_rounds_MUXInst_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_2610), .Z1_t (new_AGEMA_signal_2611), .Z1_f (new_AGEMA_signal_2612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_2610), .B1_t (new_AGEMA_signal_2611), .B1_f (new_AGEMA_signal_2612), .Z0_t (Midori_rounds_MUXInst_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_3633), .Z1_t (new_AGEMA_signal_3634), .Z1_f (new_AGEMA_signal_3635) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_3_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_3633), .A1_t (new_AGEMA_signal_3634), .A1_f (new_AGEMA_signal_3635), .B0_t (key_s0_t[67]), .B0_f (key_s0_f[67]), .B1_t (key_s1_t[67]), .B1_f (key_s1_f[67]), .Z0_t (Midori_rounds_SelectedKey[3]), .Z0_f (new_AGEMA_signal_4097), .Z1_t (new_AGEMA_signal_4098), .Z1_f (new_AGEMA_signal_4099) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_4_U1_XOR1_U1 ( .A0_t (key_s0_t[68]), .A0_f (key_s0_f[68]), .A1_t (key_s1_t[68]), .A1_f (key_s1_f[68]), .B0_t (key_s0_t[4]), .B0_f (key_s0_f[4]), .B1_t (key_s1_t[4]), .B1_f (key_s1_f[4]), .Z0_t (Midori_rounds_MUXInst_mux_inst_4_U1_X), .Z0_f (new_AGEMA_signal_2613), .Z1_t (new_AGEMA_signal_2614), .Z1_f (new_AGEMA_signal_2615) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_4_U1_X), .B0_f (new_AGEMA_signal_2613), .B1_t (new_AGEMA_signal_2614), .B1_f (new_AGEMA_signal_2615), .Z0_t (Midori_rounds_MUXInst_mux_inst_4_U1_Y), .Z0_f (new_AGEMA_signal_3636), .Z1_t (new_AGEMA_signal_3637), .Z1_f (new_AGEMA_signal_3638) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_4_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_4_U1_Y), .A0_f (new_AGEMA_signal_3636), .A1_t (new_AGEMA_signal_3637), .A1_f (new_AGEMA_signal_3638), .B0_t (key_s0_t[68]), .B0_f (key_s0_f[68]), .B1_t (key_s1_t[68]), .B1_f (key_s1_f[68]), .Z0_t (Midori_rounds_SelectedKey[4]), .Z0_f (new_AGEMA_signal_4100), .Z1_t (new_AGEMA_signal_4101), .Z1_f (new_AGEMA_signal_4102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_5_U1_XOR1_U1 ( .A0_t (key_s0_t[69]), .A0_f (key_s0_f[69]), .A1_t (key_s1_t[69]), .A1_f (key_s1_f[69]), .B0_t (key_s0_t[5]), .B0_f (key_s0_f[5]), .B1_t (key_s1_t[5]), .B1_f (key_s1_f[5]), .Z0_t (Midori_rounds_MUXInst_mux_inst_5_U1_X), .Z0_f (new_AGEMA_signal_2616), .Z1_t (new_AGEMA_signal_2617), .Z1_f (new_AGEMA_signal_2618) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_5_U1_X), .B0_f (new_AGEMA_signal_2616), .B1_t (new_AGEMA_signal_2617), .B1_f (new_AGEMA_signal_2618), .Z0_t (Midori_rounds_MUXInst_mux_inst_5_U1_Y), .Z0_f (new_AGEMA_signal_3639), .Z1_t (new_AGEMA_signal_3640), .Z1_f (new_AGEMA_signal_3641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_5_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_5_U1_Y), .A0_f (new_AGEMA_signal_3639), .A1_t (new_AGEMA_signal_3640), .A1_f (new_AGEMA_signal_3641), .B0_t (key_s0_t[69]), .B0_f (key_s0_f[69]), .B1_t (key_s1_t[69]), .B1_f (key_s1_f[69]), .Z0_t (Midori_rounds_SelectedKey[5]), .Z0_f (new_AGEMA_signal_4103), .Z1_t (new_AGEMA_signal_4104), .Z1_f (new_AGEMA_signal_4105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_6_U1_XOR1_U1 ( .A0_t (key_s0_t[70]), .A0_f (key_s0_f[70]), .A1_t (key_s1_t[70]), .A1_f (key_s1_f[70]), .B0_t (key_s0_t[6]), .B0_f (key_s0_f[6]), .B1_t (key_s1_t[6]), .B1_f (key_s1_f[6]), .Z0_t (Midori_rounds_MUXInst_mux_inst_6_U1_X), .Z0_f (new_AGEMA_signal_2619), .Z1_t (new_AGEMA_signal_2620), .Z1_f (new_AGEMA_signal_2621) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_6_U1_X), .B0_f (new_AGEMA_signal_2619), .B1_t (new_AGEMA_signal_2620), .B1_f (new_AGEMA_signal_2621), .Z0_t (Midori_rounds_MUXInst_mux_inst_6_U1_Y), .Z0_f (new_AGEMA_signal_3642), .Z1_t (new_AGEMA_signal_3643), .Z1_f (new_AGEMA_signal_3644) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_6_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_6_U1_Y), .A0_f (new_AGEMA_signal_3642), .A1_t (new_AGEMA_signal_3643), .A1_f (new_AGEMA_signal_3644), .B0_t (key_s0_t[70]), .B0_f (key_s0_f[70]), .B1_t (key_s1_t[70]), .B1_f (key_s1_f[70]), .Z0_t (Midori_rounds_SelectedKey[6]), .Z0_f (new_AGEMA_signal_4106), .Z1_t (new_AGEMA_signal_4107), .Z1_f (new_AGEMA_signal_4108) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_7_U1_XOR1_U1 ( .A0_t (key_s0_t[71]), .A0_f (key_s0_f[71]), .A1_t (key_s1_t[71]), .A1_f (key_s1_f[71]), .B0_t (key_s0_t[7]), .B0_f (key_s0_f[7]), .B1_t (key_s1_t[7]), .B1_f (key_s1_f[7]), .Z0_t (Midori_rounds_MUXInst_mux_inst_7_U1_X), .Z0_f (new_AGEMA_signal_2622), .Z1_t (new_AGEMA_signal_2623), .Z1_f (new_AGEMA_signal_2624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_7_U1_X), .B0_f (new_AGEMA_signal_2622), .B1_t (new_AGEMA_signal_2623), .B1_f (new_AGEMA_signal_2624), .Z0_t (Midori_rounds_MUXInst_mux_inst_7_U1_Y), .Z0_f (new_AGEMA_signal_3645), .Z1_t (new_AGEMA_signal_3646), .Z1_f (new_AGEMA_signal_3647) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_7_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_7_U1_Y), .A0_f (new_AGEMA_signal_3645), .A1_t (new_AGEMA_signal_3646), .A1_f (new_AGEMA_signal_3647), .B0_t (key_s0_t[71]), .B0_f (key_s0_f[71]), .B1_t (key_s1_t[71]), .B1_f (key_s1_f[71]), .Z0_t (Midori_rounds_SelectedKey[7]), .Z0_f (new_AGEMA_signal_4109), .Z1_t (new_AGEMA_signal_4110), .Z1_f (new_AGEMA_signal_4111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_8_U1_XOR1_U1 ( .A0_t (key_s0_t[72]), .A0_f (key_s0_f[72]), .A1_t (key_s1_t[72]), .A1_f (key_s1_f[72]), .B0_t (key_s0_t[8]), .B0_f (key_s0_f[8]), .B1_t (key_s1_t[8]), .B1_f (key_s1_f[8]), .Z0_t (Midori_rounds_MUXInst_mux_inst_8_U1_X), .Z0_f (new_AGEMA_signal_2625), .Z1_t (new_AGEMA_signal_2626), .Z1_f (new_AGEMA_signal_2627) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_8_U1_X), .B0_f (new_AGEMA_signal_2625), .B1_t (new_AGEMA_signal_2626), .B1_f (new_AGEMA_signal_2627), .Z0_t (Midori_rounds_MUXInst_mux_inst_8_U1_Y), .Z0_f (new_AGEMA_signal_3648), .Z1_t (new_AGEMA_signal_3649), .Z1_f (new_AGEMA_signal_3650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_8_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_8_U1_Y), .A0_f (new_AGEMA_signal_3648), .A1_t (new_AGEMA_signal_3649), .A1_f (new_AGEMA_signal_3650), .B0_t (key_s0_t[72]), .B0_f (key_s0_f[72]), .B1_t (key_s1_t[72]), .B1_f (key_s1_f[72]), .Z0_t (Midori_rounds_SelectedKey[8]), .Z0_f (new_AGEMA_signal_4112), .Z1_t (new_AGEMA_signal_4113), .Z1_f (new_AGEMA_signal_4114) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_9_U1_XOR1_U1 ( .A0_t (key_s0_t[73]), .A0_f (key_s0_f[73]), .A1_t (key_s1_t[73]), .A1_f (key_s1_f[73]), .B0_t (key_s0_t[9]), .B0_f (key_s0_f[9]), .B1_t (key_s1_t[9]), .B1_f (key_s1_f[9]), .Z0_t (Midori_rounds_MUXInst_mux_inst_9_U1_X), .Z0_f (new_AGEMA_signal_2628), .Z1_t (new_AGEMA_signal_2629), .Z1_f (new_AGEMA_signal_2630) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_9_U1_X), .B0_f (new_AGEMA_signal_2628), .B1_t (new_AGEMA_signal_2629), .B1_f (new_AGEMA_signal_2630), .Z0_t (Midori_rounds_MUXInst_mux_inst_9_U1_Y), .Z0_f (new_AGEMA_signal_3651), .Z1_t (new_AGEMA_signal_3652), .Z1_f (new_AGEMA_signal_3653) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_9_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_9_U1_Y), .A0_f (new_AGEMA_signal_3651), .A1_t (new_AGEMA_signal_3652), .A1_f (new_AGEMA_signal_3653), .B0_t (key_s0_t[73]), .B0_f (key_s0_f[73]), .B1_t (key_s1_t[73]), .B1_f (key_s1_f[73]), .Z0_t (Midori_rounds_SelectedKey[9]), .Z0_f (new_AGEMA_signal_4115), .Z1_t (new_AGEMA_signal_4116), .Z1_f (new_AGEMA_signal_4117) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_10_U1_XOR1_U1 ( .A0_t (key_s0_t[74]), .A0_f (key_s0_f[74]), .A1_t (key_s1_t[74]), .A1_f (key_s1_f[74]), .B0_t (key_s0_t[10]), .B0_f (key_s0_f[10]), .B1_t (key_s1_t[10]), .B1_f (key_s1_f[10]), .Z0_t (Midori_rounds_MUXInst_mux_inst_10_U1_X), .Z0_f (new_AGEMA_signal_2631), .Z1_t (new_AGEMA_signal_2632), .Z1_f (new_AGEMA_signal_2633) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_10_U1_X), .B0_f (new_AGEMA_signal_2631), .B1_t (new_AGEMA_signal_2632), .B1_f (new_AGEMA_signal_2633), .Z0_t (Midori_rounds_MUXInst_mux_inst_10_U1_Y), .Z0_f (new_AGEMA_signal_3654), .Z1_t (new_AGEMA_signal_3655), .Z1_f (new_AGEMA_signal_3656) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_10_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_10_U1_Y), .A0_f (new_AGEMA_signal_3654), .A1_t (new_AGEMA_signal_3655), .A1_f (new_AGEMA_signal_3656), .B0_t (key_s0_t[74]), .B0_f (key_s0_f[74]), .B1_t (key_s1_t[74]), .B1_f (key_s1_f[74]), .Z0_t (Midori_rounds_SelectedKey[10]), .Z0_f (new_AGEMA_signal_4118), .Z1_t (new_AGEMA_signal_4119), .Z1_f (new_AGEMA_signal_4120) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_11_U1_XOR1_U1 ( .A0_t (key_s0_t[75]), .A0_f (key_s0_f[75]), .A1_t (key_s1_t[75]), .A1_f (key_s1_f[75]), .B0_t (key_s0_t[11]), .B0_f (key_s0_f[11]), .B1_t (key_s1_t[11]), .B1_f (key_s1_f[11]), .Z0_t (Midori_rounds_MUXInst_mux_inst_11_U1_X), .Z0_f (new_AGEMA_signal_2634), .Z1_t (new_AGEMA_signal_2635), .Z1_f (new_AGEMA_signal_2636) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_11_U1_X), .B0_f (new_AGEMA_signal_2634), .B1_t (new_AGEMA_signal_2635), .B1_f (new_AGEMA_signal_2636), .Z0_t (Midori_rounds_MUXInst_mux_inst_11_U1_Y), .Z0_f (new_AGEMA_signal_3657), .Z1_t (new_AGEMA_signal_3658), .Z1_f (new_AGEMA_signal_3659) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_11_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_11_U1_Y), .A0_f (new_AGEMA_signal_3657), .A1_t (new_AGEMA_signal_3658), .A1_f (new_AGEMA_signal_3659), .B0_t (key_s0_t[75]), .B0_f (key_s0_f[75]), .B1_t (key_s1_t[75]), .B1_f (key_s1_f[75]), .Z0_t (Midori_rounds_SelectedKey[11]), .Z0_f (new_AGEMA_signal_4121), .Z1_t (new_AGEMA_signal_4122), .Z1_f (new_AGEMA_signal_4123) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_12_U1_XOR1_U1 ( .A0_t (key_s0_t[76]), .A0_f (key_s0_f[76]), .A1_t (key_s1_t[76]), .A1_f (key_s1_f[76]), .B0_t (key_s0_t[12]), .B0_f (key_s0_f[12]), .B1_t (key_s1_t[12]), .B1_f (key_s1_f[12]), .Z0_t (Midori_rounds_MUXInst_mux_inst_12_U1_X), .Z0_f (new_AGEMA_signal_2637), .Z1_t (new_AGEMA_signal_2638), .Z1_f (new_AGEMA_signal_2639) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_12_U1_X), .B0_f (new_AGEMA_signal_2637), .B1_t (new_AGEMA_signal_2638), .B1_f (new_AGEMA_signal_2639), .Z0_t (Midori_rounds_MUXInst_mux_inst_12_U1_Y), .Z0_f (new_AGEMA_signal_3660), .Z1_t (new_AGEMA_signal_3661), .Z1_f (new_AGEMA_signal_3662) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_12_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_12_U1_Y), .A0_f (new_AGEMA_signal_3660), .A1_t (new_AGEMA_signal_3661), .A1_f (new_AGEMA_signal_3662), .B0_t (key_s0_t[76]), .B0_f (key_s0_f[76]), .B1_t (key_s1_t[76]), .B1_f (key_s1_f[76]), .Z0_t (Midori_rounds_SelectedKey[12]), .Z0_f (new_AGEMA_signal_4124), .Z1_t (new_AGEMA_signal_4125), .Z1_f (new_AGEMA_signal_4126) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_13_U1_XOR1_U1 ( .A0_t (key_s0_t[77]), .A0_f (key_s0_f[77]), .A1_t (key_s1_t[77]), .A1_f (key_s1_f[77]), .B0_t (key_s0_t[13]), .B0_f (key_s0_f[13]), .B1_t (key_s1_t[13]), .B1_f (key_s1_f[13]), .Z0_t (Midori_rounds_MUXInst_mux_inst_13_U1_X), .Z0_f (new_AGEMA_signal_2640), .Z1_t (new_AGEMA_signal_2641), .Z1_f (new_AGEMA_signal_2642) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_13_U1_X), .B0_f (new_AGEMA_signal_2640), .B1_t (new_AGEMA_signal_2641), .B1_f (new_AGEMA_signal_2642), .Z0_t (Midori_rounds_MUXInst_mux_inst_13_U1_Y), .Z0_f (new_AGEMA_signal_3663), .Z1_t (new_AGEMA_signal_3664), .Z1_f (new_AGEMA_signal_3665) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_13_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_13_U1_Y), .A0_f (new_AGEMA_signal_3663), .A1_t (new_AGEMA_signal_3664), .A1_f (new_AGEMA_signal_3665), .B0_t (key_s0_t[77]), .B0_f (key_s0_f[77]), .B1_t (key_s1_t[77]), .B1_f (key_s1_f[77]), .Z0_t (Midori_rounds_SelectedKey[13]), .Z0_f (new_AGEMA_signal_4127), .Z1_t (new_AGEMA_signal_4128), .Z1_f (new_AGEMA_signal_4129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_14_U1_XOR1_U1 ( .A0_t (key_s0_t[78]), .A0_f (key_s0_f[78]), .A1_t (key_s1_t[78]), .A1_f (key_s1_f[78]), .B0_t (key_s0_t[14]), .B0_f (key_s0_f[14]), .B1_t (key_s1_t[14]), .B1_f (key_s1_f[14]), .Z0_t (Midori_rounds_MUXInst_mux_inst_14_U1_X), .Z0_f (new_AGEMA_signal_2643), .Z1_t (new_AGEMA_signal_2644), .Z1_f (new_AGEMA_signal_2645) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_14_U1_X), .B0_f (new_AGEMA_signal_2643), .B1_t (new_AGEMA_signal_2644), .B1_f (new_AGEMA_signal_2645), .Z0_t (Midori_rounds_MUXInst_mux_inst_14_U1_Y), .Z0_f (new_AGEMA_signal_3666), .Z1_t (new_AGEMA_signal_3667), .Z1_f (new_AGEMA_signal_3668) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_14_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_14_U1_Y), .A0_f (new_AGEMA_signal_3666), .A1_t (new_AGEMA_signal_3667), .A1_f (new_AGEMA_signal_3668), .B0_t (key_s0_t[78]), .B0_f (key_s0_f[78]), .B1_t (key_s1_t[78]), .B1_f (key_s1_f[78]), .Z0_t (Midori_rounds_SelectedKey[14]), .Z0_f (new_AGEMA_signal_4130), .Z1_t (new_AGEMA_signal_4131), .Z1_f (new_AGEMA_signal_4132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_15_U1_XOR1_U1 ( .A0_t (key_s0_t[79]), .A0_f (key_s0_f[79]), .A1_t (key_s1_t[79]), .A1_f (key_s1_f[79]), .B0_t (key_s0_t[15]), .B0_f (key_s0_f[15]), .B1_t (key_s1_t[15]), .B1_f (key_s1_f[15]), .Z0_t (Midori_rounds_MUXInst_mux_inst_15_U1_X), .Z0_f (new_AGEMA_signal_2646), .Z1_t (new_AGEMA_signal_2647), .Z1_f (new_AGEMA_signal_2648) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_15_U1_X), .B0_f (new_AGEMA_signal_2646), .B1_t (new_AGEMA_signal_2647), .B1_f (new_AGEMA_signal_2648), .Z0_t (Midori_rounds_MUXInst_mux_inst_15_U1_Y), .Z0_f (new_AGEMA_signal_3669), .Z1_t (new_AGEMA_signal_3670), .Z1_f (new_AGEMA_signal_3671) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_15_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_15_U1_Y), .A0_f (new_AGEMA_signal_3669), .A1_t (new_AGEMA_signal_3670), .A1_f (new_AGEMA_signal_3671), .B0_t (key_s0_t[79]), .B0_f (key_s0_f[79]), .B1_t (key_s1_t[79]), .B1_f (key_s1_f[79]), .Z0_t (Midori_rounds_SelectedKey[15]), .Z0_f (new_AGEMA_signal_4133), .Z1_t (new_AGEMA_signal_4134), .Z1_f (new_AGEMA_signal_4135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_16_U1_XOR1_U1 ( .A0_t (key_s0_t[80]), .A0_f (key_s0_f[80]), .A1_t (key_s1_t[80]), .A1_f (key_s1_f[80]), .B0_t (key_s0_t[16]), .B0_f (key_s0_f[16]), .B1_t (key_s1_t[16]), .B1_f (key_s1_f[16]), .Z0_t (Midori_rounds_MUXInst_mux_inst_16_U1_X), .Z0_f (new_AGEMA_signal_2649), .Z1_t (new_AGEMA_signal_2650), .Z1_f (new_AGEMA_signal_2651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_16_U1_X), .B0_f (new_AGEMA_signal_2649), .B1_t (new_AGEMA_signal_2650), .B1_f (new_AGEMA_signal_2651), .Z0_t (Midori_rounds_MUXInst_mux_inst_16_U1_Y), .Z0_f (new_AGEMA_signal_3672), .Z1_t (new_AGEMA_signal_3673), .Z1_f (new_AGEMA_signal_3674) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_16_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_16_U1_Y), .A0_f (new_AGEMA_signal_3672), .A1_t (new_AGEMA_signal_3673), .A1_f (new_AGEMA_signal_3674), .B0_t (key_s0_t[80]), .B0_f (key_s0_f[80]), .B1_t (key_s1_t[80]), .B1_f (key_s1_f[80]), .Z0_t (Midori_rounds_SelectedKey[16]), .Z0_f (new_AGEMA_signal_4136), .Z1_t (new_AGEMA_signal_4137), .Z1_f (new_AGEMA_signal_4138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_17_U1_XOR1_U1 ( .A0_t (key_s0_t[81]), .A0_f (key_s0_f[81]), .A1_t (key_s1_t[81]), .A1_f (key_s1_f[81]), .B0_t (key_s0_t[17]), .B0_f (key_s0_f[17]), .B1_t (key_s1_t[17]), .B1_f (key_s1_f[17]), .Z0_t (Midori_rounds_MUXInst_mux_inst_17_U1_X), .Z0_f (new_AGEMA_signal_2652), .Z1_t (new_AGEMA_signal_2653), .Z1_f (new_AGEMA_signal_2654) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_17_U1_X), .B0_f (new_AGEMA_signal_2652), .B1_t (new_AGEMA_signal_2653), .B1_f (new_AGEMA_signal_2654), .Z0_t (Midori_rounds_MUXInst_mux_inst_17_U1_Y), .Z0_f (new_AGEMA_signal_3675), .Z1_t (new_AGEMA_signal_3676), .Z1_f (new_AGEMA_signal_3677) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_17_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_17_U1_Y), .A0_f (new_AGEMA_signal_3675), .A1_t (new_AGEMA_signal_3676), .A1_f (new_AGEMA_signal_3677), .B0_t (key_s0_t[81]), .B0_f (key_s0_f[81]), .B1_t (key_s1_t[81]), .B1_f (key_s1_f[81]), .Z0_t (Midori_rounds_SelectedKey[17]), .Z0_f (new_AGEMA_signal_4139), .Z1_t (new_AGEMA_signal_4140), .Z1_f (new_AGEMA_signal_4141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_18_U1_XOR1_U1 ( .A0_t (key_s0_t[82]), .A0_f (key_s0_f[82]), .A1_t (key_s1_t[82]), .A1_f (key_s1_f[82]), .B0_t (key_s0_t[18]), .B0_f (key_s0_f[18]), .B1_t (key_s1_t[18]), .B1_f (key_s1_f[18]), .Z0_t (Midori_rounds_MUXInst_mux_inst_18_U1_X), .Z0_f (new_AGEMA_signal_2655), .Z1_t (new_AGEMA_signal_2656), .Z1_f (new_AGEMA_signal_2657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_18_U1_X), .B0_f (new_AGEMA_signal_2655), .B1_t (new_AGEMA_signal_2656), .B1_f (new_AGEMA_signal_2657), .Z0_t (Midori_rounds_MUXInst_mux_inst_18_U1_Y), .Z0_f (new_AGEMA_signal_3678), .Z1_t (new_AGEMA_signal_3679), .Z1_f (new_AGEMA_signal_3680) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_18_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_18_U1_Y), .A0_f (new_AGEMA_signal_3678), .A1_t (new_AGEMA_signal_3679), .A1_f (new_AGEMA_signal_3680), .B0_t (key_s0_t[82]), .B0_f (key_s0_f[82]), .B1_t (key_s1_t[82]), .B1_f (key_s1_f[82]), .Z0_t (Midori_rounds_SelectedKey[18]), .Z0_f (new_AGEMA_signal_4142), .Z1_t (new_AGEMA_signal_4143), .Z1_f (new_AGEMA_signal_4144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_19_U1_XOR1_U1 ( .A0_t (key_s0_t[83]), .A0_f (key_s0_f[83]), .A1_t (key_s1_t[83]), .A1_f (key_s1_f[83]), .B0_t (key_s0_t[19]), .B0_f (key_s0_f[19]), .B1_t (key_s1_t[19]), .B1_f (key_s1_f[19]), .Z0_t (Midori_rounds_MUXInst_mux_inst_19_U1_X), .Z0_f (new_AGEMA_signal_2658), .Z1_t (new_AGEMA_signal_2659), .Z1_f (new_AGEMA_signal_2660) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_19_U1_X), .B0_f (new_AGEMA_signal_2658), .B1_t (new_AGEMA_signal_2659), .B1_f (new_AGEMA_signal_2660), .Z0_t (Midori_rounds_MUXInst_mux_inst_19_U1_Y), .Z0_f (new_AGEMA_signal_3681), .Z1_t (new_AGEMA_signal_3682), .Z1_f (new_AGEMA_signal_3683) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_19_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_19_U1_Y), .A0_f (new_AGEMA_signal_3681), .A1_t (new_AGEMA_signal_3682), .A1_f (new_AGEMA_signal_3683), .B0_t (key_s0_t[83]), .B0_f (key_s0_f[83]), .B1_t (key_s1_t[83]), .B1_f (key_s1_f[83]), .Z0_t (Midori_rounds_SelectedKey[19]), .Z0_f (new_AGEMA_signal_4145), .Z1_t (new_AGEMA_signal_4146), .Z1_f (new_AGEMA_signal_4147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_20_U1_XOR1_U1 ( .A0_t (key_s0_t[84]), .A0_f (key_s0_f[84]), .A1_t (key_s1_t[84]), .A1_f (key_s1_f[84]), .B0_t (key_s0_t[20]), .B0_f (key_s0_f[20]), .B1_t (key_s1_t[20]), .B1_f (key_s1_f[20]), .Z0_t (Midori_rounds_MUXInst_mux_inst_20_U1_X), .Z0_f (new_AGEMA_signal_2661), .Z1_t (new_AGEMA_signal_2662), .Z1_f (new_AGEMA_signal_2663) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_20_U1_X), .B0_f (new_AGEMA_signal_2661), .B1_t (new_AGEMA_signal_2662), .B1_f (new_AGEMA_signal_2663), .Z0_t (Midori_rounds_MUXInst_mux_inst_20_U1_Y), .Z0_f (new_AGEMA_signal_3684), .Z1_t (new_AGEMA_signal_3685), .Z1_f (new_AGEMA_signal_3686) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_20_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_20_U1_Y), .A0_f (new_AGEMA_signal_3684), .A1_t (new_AGEMA_signal_3685), .A1_f (new_AGEMA_signal_3686), .B0_t (key_s0_t[84]), .B0_f (key_s0_f[84]), .B1_t (key_s1_t[84]), .B1_f (key_s1_f[84]), .Z0_t (Midori_rounds_SelectedKey[20]), .Z0_f (new_AGEMA_signal_4148), .Z1_t (new_AGEMA_signal_4149), .Z1_f (new_AGEMA_signal_4150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_21_U1_XOR1_U1 ( .A0_t (key_s0_t[85]), .A0_f (key_s0_f[85]), .A1_t (key_s1_t[85]), .A1_f (key_s1_f[85]), .B0_t (key_s0_t[21]), .B0_f (key_s0_f[21]), .B1_t (key_s1_t[21]), .B1_f (key_s1_f[21]), .Z0_t (Midori_rounds_MUXInst_mux_inst_21_U1_X), .Z0_f (new_AGEMA_signal_2664), .Z1_t (new_AGEMA_signal_2665), .Z1_f (new_AGEMA_signal_2666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_21_U1_X), .B0_f (new_AGEMA_signal_2664), .B1_t (new_AGEMA_signal_2665), .B1_f (new_AGEMA_signal_2666), .Z0_t (Midori_rounds_MUXInst_mux_inst_21_U1_Y), .Z0_f (new_AGEMA_signal_3687), .Z1_t (new_AGEMA_signal_3688), .Z1_f (new_AGEMA_signal_3689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_21_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_21_U1_Y), .A0_f (new_AGEMA_signal_3687), .A1_t (new_AGEMA_signal_3688), .A1_f (new_AGEMA_signal_3689), .B0_t (key_s0_t[85]), .B0_f (key_s0_f[85]), .B1_t (key_s1_t[85]), .B1_f (key_s1_f[85]), .Z0_t (Midori_rounds_SelectedKey[21]), .Z0_f (new_AGEMA_signal_4151), .Z1_t (new_AGEMA_signal_4152), .Z1_f (new_AGEMA_signal_4153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_22_U1_XOR1_U1 ( .A0_t (key_s0_t[86]), .A0_f (key_s0_f[86]), .A1_t (key_s1_t[86]), .A1_f (key_s1_f[86]), .B0_t (key_s0_t[22]), .B0_f (key_s0_f[22]), .B1_t (key_s1_t[22]), .B1_f (key_s1_f[22]), .Z0_t (Midori_rounds_MUXInst_mux_inst_22_U1_X), .Z0_f (new_AGEMA_signal_2667), .Z1_t (new_AGEMA_signal_2668), .Z1_f (new_AGEMA_signal_2669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_22_U1_X), .B0_f (new_AGEMA_signal_2667), .B1_t (new_AGEMA_signal_2668), .B1_f (new_AGEMA_signal_2669), .Z0_t (Midori_rounds_MUXInst_mux_inst_22_U1_Y), .Z0_f (new_AGEMA_signal_3690), .Z1_t (new_AGEMA_signal_3691), .Z1_f (new_AGEMA_signal_3692) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_22_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_22_U1_Y), .A0_f (new_AGEMA_signal_3690), .A1_t (new_AGEMA_signal_3691), .A1_f (new_AGEMA_signal_3692), .B0_t (key_s0_t[86]), .B0_f (key_s0_f[86]), .B1_t (key_s1_t[86]), .B1_f (key_s1_f[86]), .Z0_t (Midori_rounds_SelectedKey[22]), .Z0_f (new_AGEMA_signal_4154), .Z1_t (new_AGEMA_signal_4155), .Z1_f (new_AGEMA_signal_4156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_23_U1_XOR1_U1 ( .A0_t (key_s0_t[87]), .A0_f (key_s0_f[87]), .A1_t (key_s1_t[87]), .A1_f (key_s1_f[87]), .B0_t (key_s0_t[23]), .B0_f (key_s0_f[23]), .B1_t (key_s1_t[23]), .B1_f (key_s1_f[23]), .Z0_t (Midori_rounds_MUXInst_mux_inst_23_U1_X), .Z0_f (new_AGEMA_signal_2670), .Z1_t (new_AGEMA_signal_2671), .Z1_f (new_AGEMA_signal_2672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_23_U1_X), .B0_f (new_AGEMA_signal_2670), .B1_t (new_AGEMA_signal_2671), .B1_f (new_AGEMA_signal_2672), .Z0_t (Midori_rounds_MUXInst_mux_inst_23_U1_Y), .Z0_f (new_AGEMA_signal_3693), .Z1_t (new_AGEMA_signal_3694), .Z1_f (new_AGEMA_signal_3695) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_23_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_23_U1_Y), .A0_f (new_AGEMA_signal_3693), .A1_t (new_AGEMA_signal_3694), .A1_f (new_AGEMA_signal_3695), .B0_t (key_s0_t[87]), .B0_f (key_s0_f[87]), .B1_t (key_s1_t[87]), .B1_f (key_s1_f[87]), .Z0_t (Midori_rounds_SelectedKey[23]), .Z0_f (new_AGEMA_signal_4157), .Z1_t (new_AGEMA_signal_4158), .Z1_f (new_AGEMA_signal_4159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_24_U1_XOR1_U1 ( .A0_t (key_s0_t[88]), .A0_f (key_s0_f[88]), .A1_t (key_s1_t[88]), .A1_f (key_s1_f[88]), .B0_t (key_s0_t[24]), .B0_f (key_s0_f[24]), .B1_t (key_s1_t[24]), .B1_f (key_s1_f[24]), .Z0_t (Midori_rounds_MUXInst_mux_inst_24_U1_X), .Z0_f (new_AGEMA_signal_2673), .Z1_t (new_AGEMA_signal_2674), .Z1_f (new_AGEMA_signal_2675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_24_U1_X), .B0_f (new_AGEMA_signal_2673), .B1_t (new_AGEMA_signal_2674), .B1_f (new_AGEMA_signal_2675), .Z0_t (Midori_rounds_MUXInst_mux_inst_24_U1_Y), .Z0_f (new_AGEMA_signal_3696), .Z1_t (new_AGEMA_signal_3697), .Z1_f (new_AGEMA_signal_3698) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_24_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_24_U1_Y), .A0_f (new_AGEMA_signal_3696), .A1_t (new_AGEMA_signal_3697), .A1_f (new_AGEMA_signal_3698), .B0_t (key_s0_t[88]), .B0_f (key_s0_f[88]), .B1_t (key_s1_t[88]), .B1_f (key_s1_f[88]), .Z0_t (Midori_rounds_SelectedKey[24]), .Z0_f (new_AGEMA_signal_4160), .Z1_t (new_AGEMA_signal_4161), .Z1_f (new_AGEMA_signal_4162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_25_U1_XOR1_U1 ( .A0_t (key_s0_t[89]), .A0_f (key_s0_f[89]), .A1_t (key_s1_t[89]), .A1_f (key_s1_f[89]), .B0_t (key_s0_t[25]), .B0_f (key_s0_f[25]), .B1_t (key_s1_t[25]), .B1_f (key_s1_f[25]), .Z0_t (Midori_rounds_MUXInst_mux_inst_25_U1_X), .Z0_f (new_AGEMA_signal_2676), .Z1_t (new_AGEMA_signal_2677), .Z1_f (new_AGEMA_signal_2678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_25_U1_X), .B0_f (new_AGEMA_signal_2676), .B1_t (new_AGEMA_signal_2677), .B1_f (new_AGEMA_signal_2678), .Z0_t (Midori_rounds_MUXInst_mux_inst_25_U1_Y), .Z0_f (new_AGEMA_signal_3699), .Z1_t (new_AGEMA_signal_3700), .Z1_f (new_AGEMA_signal_3701) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_25_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_25_U1_Y), .A0_f (new_AGEMA_signal_3699), .A1_t (new_AGEMA_signal_3700), .A1_f (new_AGEMA_signal_3701), .B0_t (key_s0_t[89]), .B0_f (key_s0_f[89]), .B1_t (key_s1_t[89]), .B1_f (key_s1_f[89]), .Z0_t (Midori_rounds_SelectedKey[25]), .Z0_f (new_AGEMA_signal_4163), .Z1_t (new_AGEMA_signal_4164), .Z1_f (new_AGEMA_signal_4165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_26_U1_XOR1_U1 ( .A0_t (key_s0_t[90]), .A0_f (key_s0_f[90]), .A1_t (key_s1_t[90]), .A1_f (key_s1_f[90]), .B0_t (key_s0_t[26]), .B0_f (key_s0_f[26]), .B1_t (key_s1_t[26]), .B1_f (key_s1_f[26]), .Z0_t (Midori_rounds_MUXInst_mux_inst_26_U1_X), .Z0_f (new_AGEMA_signal_2679), .Z1_t (new_AGEMA_signal_2680), .Z1_f (new_AGEMA_signal_2681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_26_U1_X), .B0_f (new_AGEMA_signal_2679), .B1_t (new_AGEMA_signal_2680), .B1_f (new_AGEMA_signal_2681), .Z0_t (Midori_rounds_MUXInst_mux_inst_26_U1_Y), .Z0_f (new_AGEMA_signal_3702), .Z1_t (new_AGEMA_signal_3703), .Z1_f (new_AGEMA_signal_3704) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_26_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_26_U1_Y), .A0_f (new_AGEMA_signal_3702), .A1_t (new_AGEMA_signal_3703), .A1_f (new_AGEMA_signal_3704), .B0_t (key_s0_t[90]), .B0_f (key_s0_f[90]), .B1_t (key_s1_t[90]), .B1_f (key_s1_f[90]), .Z0_t (Midori_rounds_SelectedKey[26]), .Z0_f (new_AGEMA_signal_4166), .Z1_t (new_AGEMA_signal_4167), .Z1_f (new_AGEMA_signal_4168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_27_U1_XOR1_U1 ( .A0_t (key_s0_t[91]), .A0_f (key_s0_f[91]), .A1_t (key_s1_t[91]), .A1_f (key_s1_f[91]), .B0_t (key_s0_t[27]), .B0_f (key_s0_f[27]), .B1_t (key_s1_t[27]), .B1_f (key_s1_f[27]), .Z0_t (Midori_rounds_MUXInst_mux_inst_27_U1_X), .Z0_f (new_AGEMA_signal_2682), .Z1_t (new_AGEMA_signal_2683), .Z1_f (new_AGEMA_signal_2684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_27_U1_X), .B0_f (new_AGEMA_signal_2682), .B1_t (new_AGEMA_signal_2683), .B1_f (new_AGEMA_signal_2684), .Z0_t (Midori_rounds_MUXInst_mux_inst_27_U1_Y), .Z0_f (new_AGEMA_signal_3705), .Z1_t (new_AGEMA_signal_3706), .Z1_f (new_AGEMA_signal_3707) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_27_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_27_U1_Y), .A0_f (new_AGEMA_signal_3705), .A1_t (new_AGEMA_signal_3706), .A1_f (new_AGEMA_signal_3707), .B0_t (key_s0_t[91]), .B0_f (key_s0_f[91]), .B1_t (key_s1_t[91]), .B1_f (key_s1_f[91]), .Z0_t (Midori_rounds_SelectedKey[27]), .Z0_f (new_AGEMA_signal_4169), .Z1_t (new_AGEMA_signal_4170), .Z1_f (new_AGEMA_signal_4171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_28_U1_XOR1_U1 ( .A0_t (key_s0_t[92]), .A0_f (key_s0_f[92]), .A1_t (key_s1_t[92]), .A1_f (key_s1_f[92]), .B0_t (key_s0_t[28]), .B0_f (key_s0_f[28]), .B1_t (key_s1_t[28]), .B1_f (key_s1_f[28]), .Z0_t (Midori_rounds_MUXInst_mux_inst_28_U1_X), .Z0_f (new_AGEMA_signal_2685), .Z1_t (new_AGEMA_signal_2686), .Z1_f (new_AGEMA_signal_2687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_28_U1_X), .B0_f (new_AGEMA_signal_2685), .B1_t (new_AGEMA_signal_2686), .B1_f (new_AGEMA_signal_2687), .Z0_t (Midori_rounds_MUXInst_mux_inst_28_U1_Y), .Z0_f (new_AGEMA_signal_3708), .Z1_t (new_AGEMA_signal_3709), .Z1_f (new_AGEMA_signal_3710) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_28_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_28_U1_Y), .A0_f (new_AGEMA_signal_3708), .A1_t (new_AGEMA_signal_3709), .A1_f (new_AGEMA_signal_3710), .B0_t (key_s0_t[92]), .B0_f (key_s0_f[92]), .B1_t (key_s1_t[92]), .B1_f (key_s1_f[92]), .Z0_t (Midori_rounds_SelectedKey[28]), .Z0_f (new_AGEMA_signal_4172), .Z1_t (new_AGEMA_signal_4173), .Z1_f (new_AGEMA_signal_4174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_29_U1_XOR1_U1 ( .A0_t (key_s0_t[93]), .A0_f (key_s0_f[93]), .A1_t (key_s1_t[93]), .A1_f (key_s1_f[93]), .B0_t (key_s0_t[29]), .B0_f (key_s0_f[29]), .B1_t (key_s1_t[29]), .B1_f (key_s1_f[29]), .Z0_t (Midori_rounds_MUXInst_mux_inst_29_U1_X), .Z0_f (new_AGEMA_signal_2688), .Z1_t (new_AGEMA_signal_2689), .Z1_f (new_AGEMA_signal_2690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_29_U1_X), .B0_f (new_AGEMA_signal_2688), .B1_t (new_AGEMA_signal_2689), .B1_f (new_AGEMA_signal_2690), .Z0_t (Midori_rounds_MUXInst_mux_inst_29_U1_Y), .Z0_f (new_AGEMA_signal_3711), .Z1_t (new_AGEMA_signal_3712), .Z1_f (new_AGEMA_signal_3713) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_29_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_29_U1_Y), .A0_f (new_AGEMA_signal_3711), .A1_t (new_AGEMA_signal_3712), .A1_f (new_AGEMA_signal_3713), .B0_t (key_s0_t[93]), .B0_f (key_s0_f[93]), .B1_t (key_s1_t[93]), .B1_f (key_s1_f[93]), .Z0_t (Midori_rounds_SelectedKey[29]), .Z0_f (new_AGEMA_signal_4175), .Z1_t (new_AGEMA_signal_4176), .Z1_f (new_AGEMA_signal_4177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_30_U1_XOR1_U1 ( .A0_t (key_s0_t[94]), .A0_f (key_s0_f[94]), .A1_t (key_s1_t[94]), .A1_f (key_s1_f[94]), .B0_t (key_s0_t[30]), .B0_f (key_s0_f[30]), .B1_t (key_s1_t[30]), .B1_f (key_s1_f[30]), .Z0_t (Midori_rounds_MUXInst_mux_inst_30_U1_X), .Z0_f (new_AGEMA_signal_2691), .Z1_t (new_AGEMA_signal_2692), .Z1_f (new_AGEMA_signal_2693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_30_U1_X), .B0_f (new_AGEMA_signal_2691), .B1_t (new_AGEMA_signal_2692), .B1_f (new_AGEMA_signal_2693), .Z0_t (Midori_rounds_MUXInst_mux_inst_30_U1_Y), .Z0_f (new_AGEMA_signal_3714), .Z1_t (new_AGEMA_signal_3715), .Z1_f (new_AGEMA_signal_3716) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_30_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_30_U1_Y), .A0_f (new_AGEMA_signal_3714), .A1_t (new_AGEMA_signal_3715), .A1_f (new_AGEMA_signal_3716), .B0_t (key_s0_t[94]), .B0_f (key_s0_f[94]), .B1_t (key_s1_t[94]), .B1_f (key_s1_f[94]), .Z0_t (Midori_rounds_SelectedKey[30]), .Z0_f (new_AGEMA_signal_4178), .Z1_t (new_AGEMA_signal_4179), .Z1_f (new_AGEMA_signal_4180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_31_U1_XOR1_U1 ( .A0_t (key_s0_t[95]), .A0_f (key_s0_f[95]), .A1_t (key_s1_t[95]), .A1_f (key_s1_f[95]), .B0_t (key_s0_t[31]), .B0_f (key_s0_f[31]), .B1_t (key_s1_t[31]), .B1_f (key_s1_f[31]), .Z0_t (Midori_rounds_MUXInst_mux_inst_31_U1_X), .Z0_f (new_AGEMA_signal_2694), .Z1_t (new_AGEMA_signal_2695), .Z1_f (new_AGEMA_signal_2696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_31_U1_X), .B0_f (new_AGEMA_signal_2694), .B1_t (new_AGEMA_signal_2695), .B1_f (new_AGEMA_signal_2696), .Z0_t (Midori_rounds_MUXInst_mux_inst_31_U1_Y), .Z0_f (new_AGEMA_signal_3717), .Z1_t (new_AGEMA_signal_3718), .Z1_f (new_AGEMA_signal_3719) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_31_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_31_U1_Y), .A0_f (new_AGEMA_signal_3717), .A1_t (new_AGEMA_signal_3718), .A1_f (new_AGEMA_signal_3719), .B0_t (key_s0_t[95]), .B0_f (key_s0_f[95]), .B1_t (key_s1_t[95]), .B1_f (key_s1_f[95]), .Z0_t (Midori_rounds_SelectedKey[31]), .Z0_f (new_AGEMA_signal_4181), .Z1_t (new_AGEMA_signal_4182), .Z1_f (new_AGEMA_signal_4183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_32_U1_XOR1_U1 ( .A0_t (key_s0_t[96]), .A0_f (key_s0_f[96]), .A1_t (key_s1_t[96]), .A1_f (key_s1_f[96]), .B0_t (key_s0_t[32]), .B0_f (key_s0_f[32]), .B1_t (key_s1_t[32]), .B1_f (key_s1_f[32]), .Z0_t (Midori_rounds_MUXInst_mux_inst_32_U1_X), .Z0_f (new_AGEMA_signal_2697), .Z1_t (new_AGEMA_signal_2698), .Z1_f (new_AGEMA_signal_2699) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_32_U1_X), .B0_f (new_AGEMA_signal_2697), .B1_t (new_AGEMA_signal_2698), .B1_f (new_AGEMA_signal_2699), .Z0_t (Midori_rounds_MUXInst_mux_inst_32_U1_Y), .Z0_f (new_AGEMA_signal_3720), .Z1_t (new_AGEMA_signal_3721), .Z1_f (new_AGEMA_signal_3722) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_32_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_32_U1_Y), .A0_f (new_AGEMA_signal_3720), .A1_t (new_AGEMA_signal_3721), .A1_f (new_AGEMA_signal_3722), .B0_t (key_s0_t[96]), .B0_f (key_s0_f[96]), .B1_t (key_s1_t[96]), .B1_f (key_s1_f[96]), .Z0_t (Midori_rounds_SelectedKey[32]), .Z0_f (new_AGEMA_signal_4184), .Z1_t (new_AGEMA_signal_4185), .Z1_f (new_AGEMA_signal_4186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_33_U1_XOR1_U1 ( .A0_t (key_s0_t[97]), .A0_f (key_s0_f[97]), .A1_t (key_s1_t[97]), .A1_f (key_s1_f[97]), .B0_t (key_s0_t[33]), .B0_f (key_s0_f[33]), .B1_t (key_s1_t[33]), .B1_f (key_s1_f[33]), .Z0_t (Midori_rounds_MUXInst_mux_inst_33_U1_X), .Z0_f (new_AGEMA_signal_2700), .Z1_t (new_AGEMA_signal_2701), .Z1_f (new_AGEMA_signal_2702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_33_U1_X), .B0_f (new_AGEMA_signal_2700), .B1_t (new_AGEMA_signal_2701), .B1_f (new_AGEMA_signal_2702), .Z0_t (Midori_rounds_MUXInst_mux_inst_33_U1_Y), .Z0_f (new_AGEMA_signal_3723), .Z1_t (new_AGEMA_signal_3724), .Z1_f (new_AGEMA_signal_3725) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_33_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_33_U1_Y), .A0_f (new_AGEMA_signal_3723), .A1_t (new_AGEMA_signal_3724), .A1_f (new_AGEMA_signal_3725), .B0_t (key_s0_t[97]), .B0_f (key_s0_f[97]), .B1_t (key_s1_t[97]), .B1_f (key_s1_f[97]), .Z0_t (Midori_rounds_SelectedKey[33]), .Z0_f (new_AGEMA_signal_4187), .Z1_t (new_AGEMA_signal_4188), .Z1_f (new_AGEMA_signal_4189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_34_U1_XOR1_U1 ( .A0_t (key_s0_t[98]), .A0_f (key_s0_f[98]), .A1_t (key_s1_t[98]), .A1_f (key_s1_f[98]), .B0_t (key_s0_t[34]), .B0_f (key_s0_f[34]), .B1_t (key_s1_t[34]), .B1_f (key_s1_f[34]), .Z0_t (Midori_rounds_MUXInst_mux_inst_34_U1_X), .Z0_f (new_AGEMA_signal_2703), .Z1_t (new_AGEMA_signal_2704), .Z1_f (new_AGEMA_signal_2705) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_34_U1_X), .B0_f (new_AGEMA_signal_2703), .B1_t (new_AGEMA_signal_2704), .B1_f (new_AGEMA_signal_2705), .Z0_t (Midori_rounds_MUXInst_mux_inst_34_U1_Y), .Z0_f (new_AGEMA_signal_3726), .Z1_t (new_AGEMA_signal_3727), .Z1_f (new_AGEMA_signal_3728) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_34_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_34_U1_Y), .A0_f (new_AGEMA_signal_3726), .A1_t (new_AGEMA_signal_3727), .A1_f (new_AGEMA_signal_3728), .B0_t (key_s0_t[98]), .B0_f (key_s0_f[98]), .B1_t (key_s1_t[98]), .B1_f (key_s1_f[98]), .Z0_t (Midori_rounds_SelectedKey[34]), .Z0_f (new_AGEMA_signal_4190), .Z1_t (new_AGEMA_signal_4191), .Z1_f (new_AGEMA_signal_4192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_35_U1_XOR1_U1 ( .A0_t (key_s0_t[99]), .A0_f (key_s0_f[99]), .A1_t (key_s1_t[99]), .A1_f (key_s1_f[99]), .B0_t (key_s0_t[35]), .B0_f (key_s0_f[35]), .B1_t (key_s1_t[35]), .B1_f (key_s1_f[35]), .Z0_t (Midori_rounds_MUXInst_mux_inst_35_U1_X), .Z0_f (new_AGEMA_signal_2706), .Z1_t (new_AGEMA_signal_2707), .Z1_f (new_AGEMA_signal_2708) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_35_U1_X), .B0_f (new_AGEMA_signal_2706), .B1_t (new_AGEMA_signal_2707), .B1_f (new_AGEMA_signal_2708), .Z0_t (Midori_rounds_MUXInst_mux_inst_35_U1_Y), .Z0_f (new_AGEMA_signal_3729), .Z1_t (new_AGEMA_signal_3730), .Z1_f (new_AGEMA_signal_3731) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_35_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_35_U1_Y), .A0_f (new_AGEMA_signal_3729), .A1_t (new_AGEMA_signal_3730), .A1_f (new_AGEMA_signal_3731), .B0_t (key_s0_t[99]), .B0_f (key_s0_f[99]), .B1_t (key_s1_t[99]), .B1_f (key_s1_f[99]), .Z0_t (Midori_rounds_SelectedKey[35]), .Z0_f (new_AGEMA_signal_4193), .Z1_t (new_AGEMA_signal_4194), .Z1_f (new_AGEMA_signal_4195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_36_U1_XOR1_U1 ( .A0_t (key_s0_t[100]), .A0_f (key_s0_f[100]), .A1_t (key_s1_t[100]), .A1_f (key_s1_f[100]), .B0_t (key_s0_t[36]), .B0_f (key_s0_f[36]), .B1_t (key_s1_t[36]), .B1_f (key_s1_f[36]), .Z0_t (Midori_rounds_MUXInst_mux_inst_36_U1_X), .Z0_f (new_AGEMA_signal_2709), .Z1_t (new_AGEMA_signal_2710), .Z1_f (new_AGEMA_signal_2711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_36_U1_X), .B0_f (new_AGEMA_signal_2709), .B1_t (new_AGEMA_signal_2710), .B1_f (new_AGEMA_signal_2711), .Z0_t (Midori_rounds_MUXInst_mux_inst_36_U1_Y), .Z0_f (new_AGEMA_signal_3732), .Z1_t (new_AGEMA_signal_3733), .Z1_f (new_AGEMA_signal_3734) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_36_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_36_U1_Y), .A0_f (new_AGEMA_signal_3732), .A1_t (new_AGEMA_signal_3733), .A1_f (new_AGEMA_signal_3734), .B0_t (key_s0_t[100]), .B0_f (key_s0_f[100]), .B1_t (key_s1_t[100]), .B1_f (key_s1_f[100]), .Z0_t (Midori_rounds_SelectedKey[36]), .Z0_f (new_AGEMA_signal_4196), .Z1_t (new_AGEMA_signal_4197), .Z1_f (new_AGEMA_signal_4198) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_37_U1_XOR1_U1 ( .A0_t (key_s0_t[101]), .A0_f (key_s0_f[101]), .A1_t (key_s1_t[101]), .A1_f (key_s1_f[101]), .B0_t (key_s0_t[37]), .B0_f (key_s0_f[37]), .B1_t (key_s1_t[37]), .B1_f (key_s1_f[37]), .Z0_t (Midori_rounds_MUXInst_mux_inst_37_U1_X), .Z0_f (new_AGEMA_signal_2712), .Z1_t (new_AGEMA_signal_2713), .Z1_f (new_AGEMA_signal_2714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_37_U1_X), .B0_f (new_AGEMA_signal_2712), .B1_t (new_AGEMA_signal_2713), .B1_f (new_AGEMA_signal_2714), .Z0_t (Midori_rounds_MUXInst_mux_inst_37_U1_Y), .Z0_f (new_AGEMA_signal_3735), .Z1_t (new_AGEMA_signal_3736), .Z1_f (new_AGEMA_signal_3737) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_37_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_37_U1_Y), .A0_f (new_AGEMA_signal_3735), .A1_t (new_AGEMA_signal_3736), .A1_f (new_AGEMA_signal_3737), .B0_t (key_s0_t[101]), .B0_f (key_s0_f[101]), .B1_t (key_s1_t[101]), .B1_f (key_s1_f[101]), .Z0_t (Midori_rounds_SelectedKey[37]), .Z0_f (new_AGEMA_signal_4199), .Z1_t (new_AGEMA_signal_4200), .Z1_f (new_AGEMA_signal_4201) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_38_U1_XOR1_U1 ( .A0_t (key_s0_t[102]), .A0_f (key_s0_f[102]), .A1_t (key_s1_t[102]), .A1_f (key_s1_f[102]), .B0_t (key_s0_t[38]), .B0_f (key_s0_f[38]), .B1_t (key_s1_t[38]), .B1_f (key_s1_f[38]), .Z0_t (Midori_rounds_MUXInst_mux_inst_38_U1_X), .Z0_f (new_AGEMA_signal_2715), .Z1_t (new_AGEMA_signal_2716), .Z1_f (new_AGEMA_signal_2717) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_38_U1_X), .B0_f (new_AGEMA_signal_2715), .B1_t (new_AGEMA_signal_2716), .B1_f (new_AGEMA_signal_2717), .Z0_t (Midori_rounds_MUXInst_mux_inst_38_U1_Y), .Z0_f (new_AGEMA_signal_3738), .Z1_t (new_AGEMA_signal_3739), .Z1_f (new_AGEMA_signal_3740) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_38_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_38_U1_Y), .A0_f (new_AGEMA_signal_3738), .A1_t (new_AGEMA_signal_3739), .A1_f (new_AGEMA_signal_3740), .B0_t (key_s0_t[102]), .B0_f (key_s0_f[102]), .B1_t (key_s1_t[102]), .B1_f (key_s1_f[102]), .Z0_t (Midori_rounds_SelectedKey[38]), .Z0_f (new_AGEMA_signal_4202), .Z1_t (new_AGEMA_signal_4203), .Z1_f (new_AGEMA_signal_4204) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_39_U1_XOR1_U1 ( .A0_t (key_s0_t[103]), .A0_f (key_s0_f[103]), .A1_t (key_s1_t[103]), .A1_f (key_s1_f[103]), .B0_t (key_s0_t[39]), .B0_f (key_s0_f[39]), .B1_t (key_s1_t[39]), .B1_f (key_s1_f[39]), .Z0_t (Midori_rounds_MUXInst_mux_inst_39_U1_X), .Z0_f (new_AGEMA_signal_2718), .Z1_t (new_AGEMA_signal_2719), .Z1_f (new_AGEMA_signal_2720) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_39_U1_X), .B0_f (new_AGEMA_signal_2718), .B1_t (new_AGEMA_signal_2719), .B1_f (new_AGEMA_signal_2720), .Z0_t (Midori_rounds_MUXInst_mux_inst_39_U1_Y), .Z0_f (new_AGEMA_signal_3741), .Z1_t (new_AGEMA_signal_3742), .Z1_f (new_AGEMA_signal_3743) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_39_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_39_U1_Y), .A0_f (new_AGEMA_signal_3741), .A1_t (new_AGEMA_signal_3742), .A1_f (new_AGEMA_signal_3743), .B0_t (key_s0_t[103]), .B0_f (key_s0_f[103]), .B1_t (key_s1_t[103]), .B1_f (key_s1_f[103]), .Z0_t (Midori_rounds_SelectedKey[39]), .Z0_f (new_AGEMA_signal_4205), .Z1_t (new_AGEMA_signal_4206), .Z1_f (new_AGEMA_signal_4207) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_40_U1_XOR1_U1 ( .A0_t (key_s0_t[104]), .A0_f (key_s0_f[104]), .A1_t (key_s1_t[104]), .A1_f (key_s1_f[104]), .B0_t (key_s0_t[40]), .B0_f (key_s0_f[40]), .B1_t (key_s1_t[40]), .B1_f (key_s1_f[40]), .Z0_t (Midori_rounds_MUXInst_mux_inst_40_U1_X), .Z0_f (new_AGEMA_signal_2721), .Z1_t (new_AGEMA_signal_2722), .Z1_f (new_AGEMA_signal_2723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_40_U1_X), .B0_f (new_AGEMA_signal_2721), .B1_t (new_AGEMA_signal_2722), .B1_f (new_AGEMA_signal_2723), .Z0_t (Midori_rounds_MUXInst_mux_inst_40_U1_Y), .Z0_f (new_AGEMA_signal_3744), .Z1_t (new_AGEMA_signal_3745), .Z1_f (new_AGEMA_signal_3746) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_40_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_40_U1_Y), .A0_f (new_AGEMA_signal_3744), .A1_t (new_AGEMA_signal_3745), .A1_f (new_AGEMA_signal_3746), .B0_t (key_s0_t[104]), .B0_f (key_s0_f[104]), .B1_t (key_s1_t[104]), .B1_f (key_s1_f[104]), .Z0_t (Midori_rounds_SelectedKey[40]), .Z0_f (new_AGEMA_signal_4208), .Z1_t (new_AGEMA_signal_4209), .Z1_f (new_AGEMA_signal_4210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_41_U1_XOR1_U1 ( .A0_t (key_s0_t[105]), .A0_f (key_s0_f[105]), .A1_t (key_s1_t[105]), .A1_f (key_s1_f[105]), .B0_t (key_s0_t[41]), .B0_f (key_s0_f[41]), .B1_t (key_s1_t[41]), .B1_f (key_s1_f[41]), .Z0_t (Midori_rounds_MUXInst_mux_inst_41_U1_X), .Z0_f (new_AGEMA_signal_2724), .Z1_t (new_AGEMA_signal_2725), .Z1_f (new_AGEMA_signal_2726) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_41_U1_X), .B0_f (new_AGEMA_signal_2724), .B1_t (new_AGEMA_signal_2725), .B1_f (new_AGEMA_signal_2726), .Z0_t (Midori_rounds_MUXInst_mux_inst_41_U1_Y), .Z0_f (new_AGEMA_signal_3747), .Z1_t (new_AGEMA_signal_3748), .Z1_f (new_AGEMA_signal_3749) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_41_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_41_U1_Y), .A0_f (new_AGEMA_signal_3747), .A1_t (new_AGEMA_signal_3748), .A1_f (new_AGEMA_signal_3749), .B0_t (key_s0_t[105]), .B0_f (key_s0_f[105]), .B1_t (key_s1_t[105]), .B1_f (key_s1_f[105]), .Z0_t (Midori_rounds_SelectedKey[41]), .Z0_f (new_AGEMA_signal_4211), .Z1_t (new_AGEMA_signal_4212), .Z1_f (new_AGEMA_signal_4213) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_42_U1_XOR1_U1 ( .A0_t (key_s0_t[106]), .A0_f (key_s0_f[106]), .A1_t (key_s1_t[106]), .A1_f (key_s1_f[106]), .B0_t (key_s0_t[42]), .B0_f (key_s0_f[42]), .B1_t (key_s1_t[42]), .B1_f (key_s1_f[42]), .Z0_t (Midori_rounds_MUXInst_mux_inst_42_U1_X), .Z0_f (new_AGEMA_signal_2727), .Z1_t (new_AGEMA_signal_2728), .Z1_f (new_AGEMA_signal_2729) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_42_U1_X), .B0_f (new_AGEMA_signal_2727), .B1_t (new_AGEMA_signal_2728), .B1_f (new_AGEMA_signal_2729), .Z0_t (Midori_rounds_MUXInst_mux_inst_42_U1_Y), .Z0_f (new_AGEMA_signal_3750), .Z1_t (new_AGEMA_signal_3751), .Z1_f (new_AGEMA_signal_3752) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_42_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_42_U1_Y), .A0_f (new_AGEMA_signal_3750), .A1_t (new_AGEMA_signal_3751), .A1_f (new_AGEMA_signal_3752), .B0_t (key_s0_t[106]), .B0_f (key_s0_f[106]), .B1_t (key_s1_t[106]), .B1_f (key_s1_f[106]), .Z0_t (Midori_rounds_SelectedKey[42]), .Z0_f (new_AGEMA_signal_4214), .Z1_t (new_AGEMA_signal_4215), .Z1_f (new_AGEMA_signal_4216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_43_U1_XOR1_U1 ( .A0_t (key_s0_t[107]), .A0_f (key_s0_f[107]), .A1_t (key_s1_t[107]), .A1_f (key_s1_f[107]), .B0_t (key_s0_t[43]), .B0_f (key_s0_f[43]), .B1_t (key_s1_t[43]), .B1_f (key_s1_f[43]), .Z0_t (Midori_rounds_MUXInst_mux_inst_43_U1_X), .Z0_f (new_AGEMA_signal_2730), .Z1_t (new_AGEMA_signal_2731), .Z1_f (new_AGEMA_signal_2732) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_43_U1_X), .B0_f (new_AGEMA_signal_2730), .B1_t (new_AGEMA_signal_2731), .B1_f (new_AGEMA_signal_2732), .Z0_t (Midori_rounds_MUXInst_mux_inst_43_U1_Y), .Z0_f (new_AGEMA_signal_3753), .Z1_t (new_AGEMA_signal_3754), .Z1_f (new_AGEMA_signal_3755) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_43_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_43_U1_Y), .A0_f (new_AGEMA_signal_3753), .A1_t (new_AGEMA_signal_3754), .A1_f (new_AGEMA_signal_3755), .B0_t (key_s0_t[107]), .B0_f (key_s0_f[107]), .B1_t (key_s1_t[107]), .B1_f (key_s1_f[107]), .Z0_t (Midori_rounds_SelectedKey[43]), .Z0_f (new_AGEMA_signal_4217), .Z1_t (new_AGEMA_signal_4218), .Z1_f (new_AGEMA_signal_4219) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_44_U1_XOR1_U1 ( .A0_t (key_s0_t[108]), .A0_f (key_s0_f[108]), .A1_t (key_s1_t[108]), .A1_f (key_s1_f[108]), .B0_t (key_s0_t[44]), .B0_f (key_s0_f[44]), .B1_t (key_s1_t[44]), .B1_f (key_s1_f[44]), .Z0_t (Midori_rounds_MUXInst_mux_inst_44_U1_X), .Z0_f (new_AGEMA_signal_2733), .Z1_t (new_AGEMA_signal_2734), .Z1_f (new_AGEMA_signal_2735) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_44_U1_X), .B0_f (new_AGEMA_signal_2733), .B1_t (new_AGEMA_signal_2734), .B1_f (new_AGEMA_signal_2735), .Z0_t (Midori_rounds_MUXInst_mux_inst_44_U1_Y), .Z0_f (new_AGEMA_signal_3756), .Z1_t (new_AGEMA_signal_3757), .Z1_f (new_AGEMA_signal_3758) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_44_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_44_U1_Y), .A0_f (new_AGEMA_signal_3756), .A1_t (new_AGEMA_signal_3757), .A1_f (new_AGEMA_signal_3758), .B0_t (key_s0_t[108]), .B0_f (key_s0_f[108]), .B1_t (key_s1_t[108]), .B1_f (key_s1_f[108]), .Z0_t (Midori_rounds_SelectedKey[44]), .Z0_f (new_AGEMA_signal_4220), .Z1_t (new_AGEMA_signal_4221), .Z1_f (new_AGEMA_signal_4222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_45_U1_XOR1_U1 ( .A0_t (key_s0_t[109]), .A0_f (key_s0_f[109]), .A1_t (key_s1_t[109]), .A1_f (key_s1_f[109]), .B0_t (key_s0_t[45]), .B0_f (key_s0_f[45]), .B1_t (key_s1_t[45]), .B1_f (key_s1_f[45]), .Z0_t (Midori_rounds_MUXInst_mux_inst_45_U1_X), .Z0_f (new_AGEMA_signal_2736), .Z1_t (new_AGEMA_signal_2737), .Z1_f (new_AGEMA_signal_2738) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_45_U1_X), .B0_f (new_AGEMA_signal_2736), .B1_t (new_AGEMA_signal_2737), .B1_f (new_AGEMA_signal_2738), .Z0_t (Midori_rounds_MUXInst_mux_inst_45_U1_Y), .Z0_f (new_AGEMA_signal_3759), .Z1_t (new_AGEMA_signal_3760), .Z1_f (new_AGEMA_signal_3761) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_45_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_45_U1_Y), .A0_f (new_AGEMA_signal_3759), .A1_t (new_AGEMA_signal_3760), .A1_f (new_AGEMA_signal_3761), .B0_t (key_s0_t[109]), .B0_f (key_s0_f[109]), .B1_t (key_s1_t[109]), .B1_f (key_s1_f[109]), .Z0_t (Midori_rounds_SelectedKey[45]), .Z0_f (new_AGEMA_signal_4223), .Z1_t (new_AGEMA_signal_4224), .Z1_f (new_AGEMA_signal_4225) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_46_U1_XOR1_U1 ( .A0_t (key_s0_t[110]), .A0_f (key_s0_f[110]), .A1_t (key_s1_t[110]), .A1_f (key_s1_f[110]), .B0_t (key_s0_t[46]), .B0_f (key_s0_f[46]), .B1_t (key_s1_t[46]), .B1_f (key_s1_f[46]), .Z0_t (Midori_rounds_MUXInst_mux_inst_46_U1_X), .Z0_f (new_AGEMA_signal_2739), .Z1_t (new_AGEMA_signal_2740), .Z1_f (new_AGEMA_signal_2741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_46_U1_X), .B0_f (new_AGEMA_signal_2739), .B1_t (new_AGEMA_signal_2740), .B1_f (new_AGEMA_signal_2741), .Z0_t (Midori_rounds_MUXInst_mux_inst_46_U1_Y), .Z0_f (new_AGEMA_signal_3762), .Z1_t (new_AGEMA_signal_3763), .Z1_f (new_AGEMA_signal_3764) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_46_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_46_U1_Y), .A0_f (new_AGEMA_signal_3762), .A1_t (new_AGEMA_signal_3763), .A1_f (new_AGEMA_signal_3764), .B0_t (key_s0_t[110]), .B0_f (key_s0_f[110]), .B1_t (key_s1_t[110]), .B1_f (key_s1_f[110]), .Z0_t (Midori_rounds_SelectedKey[46]), .Z0_f (new_AGEMA_signal_4226), .Z1_t (new_AGEMA_signal_4227), .Z1_f (new_AGEMA_signal_4228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_47_U1_XOR1_U1 ( .A0_t (key_s0_t[111]), .A0_f (key_s0_f[111]), .A1_t (key_s1_t[111]), .A1_f (key_s1_f[111]), .B0_t (key_s0_t[47]), .B0_f (key_s0_f[47]), .B1_t (key_s1_t[47]), .B1_f (key_s1_f[47]), .Z0_t (Midori_rounds_MUXInst_mux_inst_47_U1_X), .Z0_f (new_AGEMA_signal_2742), .Z1_t (new_AGEMA_signal_2743), .Z1_f (new_AGEMA_signal_2744) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_47_U1_X), .B0_f (new_AGEMA_signal_2742), .B1_t (new_AGEMA_signal_2743), .B1_f (new_AGEMA_signal_2744), .Z0_t (Midori_rounds_MUXInst_mux_inst_47_U1_Y), .Z0_f (new_AGEMA_signal_3765), .Z1_t (new_AGEMA_signal_3766), .Z1_f (new_AGEMA_signal_3767) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_47_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_47_U1_Y), .A0_f (new_AGEMA_signal_3765), .A1_t (new_AGEMA_signal_3766), .A1_f (new_AGEMA_signal_3767), .B0_t (key_s0_t[111]), .B0_f (key_s0_f[111]), .B1_t (key_s1_t[111]), .B1_f (key_s1_f[111]), .Z0_t (Midori_rounds_SelectedKey[47]), .Z0_f (new_AGEMA_signal_4229), .Z1_t (new_AGEMA_signal_4230), .Z1_f (new_AGEMA_signal_4231) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_48_U1_XOR1_U1 ( .A0_t (key_s0_t[112]), .A0_f (key_s0_f[112]), .A1_t (key_s1_t[112]), .A1_f (key_s1_f[112]), .B0_t (key_s0_t[48]), .B0_f (key_s0_f[48]), .B1_t (key_s1_t[48]), .B1_f (key_s1_f[48]), .Z0_t (Midori_rounds_MUXInst_mux_inst_48_U1_X), .Z0_f (new_AGEMA_signal_2745), .Z1_t (new_AGEMA_signal_2746), .Z1_f (new_AGEMA_signal_2747) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_48_U1_X), .B0_f (new_AGEMA_signal_2745), .B1_t (new_AGEMA_signal_2746), .B1_f (new_AGEMA_signal_2747), .Z0_t (Midori_rounds_MUXInst_mux_inst_48_U1_Y), .Z0_f (new_AGEMA_signal_3768), .Z1_t (new_AGEMA_signal_3769), .Z1_f (new_AGEMA_signal_3770) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_48_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_48_U1_Y), .A0_f (new_AGEMA_signal_3768), .A1_t (new_AGEMA_signal_3769), .A1_f (new_AGEMA_signal_3770), .B0_t (key_s0_t[112]), .B0_f (key_s0_f[112]), .B1_t (key_s1_t[112]), .B1_f (key_s1_f[112]), .Z0_t (Midori_rounds_SelectedKey[48]), .Z0_f (new_AGEMA_signal_4232), .Z1_t (new_AGEMA_signal_4233), .Z1_f (new_AGEMA_signal_4234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_49_U1_XOR1_U1 ( .A0_t (key_s0_t[113]), .A0_f (key_s0_f[113]), .A1_t (key_s1_t[113]), .A1_f (key_s1_f[113]), .B0_t (key_s0_t[49]), .B0_f (key_s0_f[49]), .B1_t (key_s1_t[49]), .B1_f (key_s1_f[49]), .Z0_t (Midori_rounds_MUXInst_mux_inst_49_U1_X), .Z0_f (new_AGEMA_signal_2748), .Z1_t (new_AGEMA_signal_2749), .Z1_f (new_AGEMA_signal_2750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_49_U1_X), .B0_f (new_AGEMA_signal_2748), .B1_t (new_AGEMA_signal_2749), .B1_f (new_AGEMA_signal_2750), .Z0_t (Midori_rounds_MUXInst_mux_inst_49_U1_Y), .Z0_f (new_AGEMA_signal_3771), .Z1_t (new_AGEMA_signal_3772), .Z1_f (new_AGEMA_signal_3773) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_49_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_49_U1_Y), .A0_f (new_AGEMA_signal_3771), .A1_t (new_AGEMA_signal_3772), .A1_f (new_AGEMA_signal_3773), .B0_t (key_s0_t[113]), .B0_f (key_s0_f[113]), .B1_t (key_s1_t[113]), .B1_f (key_s1_f[113]), .Z0_t (Midori_rounds_SelectedKey[49]), .Z0_f (new_AGEMA_signal_4235), .Z1_t (new_AGEMA_signal_4236), .Z1_f (new_AGEMA_signal_4237) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_50_U1_XOR1_U1 ( .A0_t (key_s0_t[114]), .A0_f (key_s0_f[114]), .A1_t (key_s1_t[114]), .A1_f (key_s1_f[114]), .B0_t (key_s0_t[50]), .B0_f (key_s0_f[50]), .B1_t (key_s1_t[50]), .B1_f (key_s1_f[50]), .Z0_t (Midori_rounds_MUXInst_mux_inst_50_U1_X), .Z0_f (new_AGEMA_signal_2751), .Z1_t (new_AGEMA_signal_2752), .Z1_f (new_AGEMA_signal_2753) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_50_U1_X), .B0_f (new_AGEMA_signal_2751), .B1_t (new_AGEMA_signal_2752), .B1_f (new_AGEMA_signal_2753), .Z0_t (Midori_rounds_MUXInst_mux_inst_50_U1_Y), .Z0_f (new_AGEMA_signal_3774), .Z1_t (new_AGEMA_signal_3775), .Z1_f (new_AGEMA_signal_3776) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_50_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_50_U1_Y), .A0_f (new_AGEMA_signal_3774), .A1_t (new_AGEMA_signal_3775), .A1_f (new_AGEMA_signal_3776), .B0_t (key_s0_t[114]), .B0_f (key_s0_f[114]), .B1_t (key_s1_t[114]), .B1_f (key_s1_f[114]), .Z0_t (Midori_rounds_SelectedKey[50]), .Z0_f (new_AGEMA_signal_4238), .Z1_t (new_AGEMA_signal_4239), .Z1_f (new_AGEMA_signal_4240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_51_U1_XOR1_U1 ( .A0_t (key_s0_t[115]), .A0_f (key_s0_f[115]), .A1_t (key_s1_t[115]), .A1_f (key_s1_f[115]), .B0_t (key_s0_t[51]), .B0_f (key_s0_f[51]), .B1_t (key_s1_t[51]), .B1_f (key_s1_f[51]), .Z0_t (Midori_rounds_MUXInst_mux_inst_51_U1_X), .Z0_f (new_AGEMA_signal_2754), .Z1_t (new_AGEMA_signal_2755), .Z1_f (new_AGEMA_signal_2756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_51_U1_X), .B0_f (new_AGEMA_signal_2754), .B1_t (new_AGEMA_signal_2755), .B1_f (new_AGEMA_signal_2756), .Z0_t (Midori_rounds_MUXInst_mux_inst_51_U1_Y), .Z0_f (new_AGEMA_signal_3777), .Z1_t (new_AGEMA_signal_3778), .Z1_f (new_AGEMA_signal_3779) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_51_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_51_U1_Y), .A0_f (new_AGEMA_signal_3777), .A1_t (new_AGEMA_signal_3778), .A1_f (new_AGEMA_signal_3779), .B0_t (key_s0_t[115]), .B0_f (key_s0_f[115]), .B1_t (key_s1_t[115]), .B1_f (key_s1_f[115]), .Z0_t (Midori_rounds_SelectedKey[51]), .Z0_f (new_AGEMA_signal_4241), .Z1_t (new_AGEMA_signal_4242), .Z1_f (new_AGEMA_signal_4243) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_52_U1_XOR1_U1 ( .A0_t (key_s0_t[116]), .A0_f (key_s0_f[116]), .A1_t (key_s1_t[116]), .A1_f (key_s1_f[116]), .B0_t (key_s0_t[52]), .B0_f (key_s0_f[52]), .B1_t (key_s1_t[52]), .B1_f (key_s1_f[52]), .Z0_t (Midori_rounds_MUXInst_mux_inst_52_U1_X), .Z0_f (new_AGEMA_signal_2757), .Z1_t (new_AGEMA_signal_2758), .Z1_f (new_AGEMA_signal_2759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_52_U1_X), .B0_f (new_AGEMA_signal_2757), .B1_t (new_AGEMA_signal_2758), .B1_f (new_AGEMA_signal_2759), .Z0_t (Midori_rounds_MUXInst_mux_inst_52_U1_Y), .Z0_f (new_AGEMA_signal_3780), .Z1_t (new_AGEMA_signal_3781), .Z1_f (new_AGEMA_signal_3782) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_52_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_52_U1_Y), .A0_f (new_AGEMA_signal_3780), .A1_t (new_AGEMA_signal_3781), .A1_f (new_AGEMA_signal_3782), .B0_t (key_s0_t[116]), .B0_f (key_s0_f[116]), .B1_t (key_s1_t[116]), .B1_f (key_s1_f[116]), .Z0_t (Midori_rounds_SelectedKey[52]), .Z0_f (new_AGEMA_signal_4244), .Z1_t (new_AGEMA_signal_4245), .Z1_f (new_AGEMA_signal_4246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_53_U1_XOR1_U1 ( .A0_t (key_s0_t[117]), .A0_f (key_s0_f[117]), .A1_t (key_s1_t[117]), .A1_f (key_s1_f[117]), .B0_t (key_s0_t[53]), .B0_f (key_s0_f[53]), .B1_t (key_s1_t[53]), .B1_f (key_s1_f[53]), .Z0_t (Midori_rounds_MUXInst_mux_inst_53_U1_X), .Z0_f (new_AGEMA_signal_2760), .Z1_t (new_AGEMA_signal_2761), .Z1_f (new_AGEMA_signal_2762) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_53_U1_X), .B0_f (new_AGEMA_signal_2760), .B1_t (new_AGEMA_signal_2761), .B1_f (new_AGEMA_signal_2762), .Z0_t (Midori_rounds_MUXInst_mux_inst_53_U1_Y), .Z0_f (new_AGEMA_signal_3783), .Z1_t (new_AGEMA_signal_3784), .Z1_f (new_AGEMA_signal_3785) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_53_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_53_U1_Y), .A0_f (new_AGEMA_signal_3783), .A1_t (new_AGEMA_signal_3784), .A1_f (new_AGEMA_signal_3785), .B0_t (key_s0_t[117]), .B0_f (key_s0_f[117]), .B1_t (key_s1_t[117]), .B1_f (key_s1_f[117]), .Z0_t (Midori_rounds_SelectedKey[53]), .Z0_f (new_AGEMA_signal_4247), .Z1_t (new_AGEMA_signal_4248), .Z1_f (new_AGEMA_signal_4249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_54_U1_XOR1_U1 ( .A0_t (key_s0_t[118]), .A0_f (key_s0_f[118]), .A1_t (key_s1_t[118]), .A1_f (key_s1_f[118]), .B0_t (key_s0_t[54]), .B0_f (key_s0_f[54]), .B1_t (key_s1_t[54]), .B1_f (key_s1_f[54]), .Z0_t (Midori_rounds_MUXInst_mux_inst_54_U1_X), .Z0_f (new_AGEMA_signal_2763), .Z1_t (new_AGEMA_signal_2764), .Z1_f (new_AGEMA_signal_2765) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_54_U1_X), .B0_f (new_AGEMA_signal_2763), .B1_t (new_AGEMA_signal_2764), .B1_f (new_AGEMA_signal_2765), .Z0_t (Midori_rounds_MUXInst_mux_inst_54_U1_Y), .Z0_f (new_AGEMA_signal_3786), .Z1_t (new_AGEMA_signal_3787), .Z1_f (new_AGEMA_signal_3788) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_54_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_54_U1_Y), .A0_f (new_AGEMA_signal_3786), .A1_t (new_AGEMA_signal_3787), .A1_f (new_AGEMA_signal_3788), .B0_t (key_s0_t[118]), .B0_f (key_s0_f[118]), .B1_t (key_s1_t[118]), .B1_f (key_s1_f[118]), .Z0_t (Midori_rounds_SelectedKey[54]), .Z0_f (new_AGEMA_signal_4250), .Z1_t (new_AGEMA_signal_4251), .Z1_f (new_AGEMA_signal_4252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_55_U1_XOR1_U1 ( .A0_t (key_s0_t[119]), .A0_f (key_s0_f[119]), .A1_t (key_s1_t[119]), .A1_f (key_s1_f[119]), .B0_t (key_s0_t[55]), .B0_f (key_s0_f[55]), .B1_t (key_s1_t[55]), .B1_f (key_s1_f[55]), .Z0_t (Midori_rounds_MUXInst_mux_inst_55_U1_X), .Z0_f (new_AGEMA_signal_2766), .Z1_t (new_AGEMA_signal_2767), .Z1_f (new_AGEMA_signal_2768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_55_U1_X), .B0_f (new_AGEMA_signal_2766), .B1_t (new_AGEMA_signal_2767), .B1_f (new_AGEMA_signal_2768), .Z0_t (Midori_rounds_MUXInst_mux_inst_55_U1_Y), .Z0_f (new_AGEMA_signal_3789), .Z1_t (new_AGEMA_signal_3790), .Z1_f (new_AGEMA_signal_3791) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_55_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_55_U1_Y), .A0_f (new_AGEMA_signal_3789), .A1_t (new_AGEMA_signal_3790), .A1_f (new_AGEMA_signal_3791), .B0_t (key_s0_t[119]), .B0_f (key_s0_f[119]), .B1_t (key_s1_t[119]), .B1_f (key_s1_f[119]), .Z0_t (Midori_rounds_SelectedKey[55]), .Z0_f (new_AGEMA_signal_4253), .Z1_t (new_AGEMA_signal_4254), .Z1_f (new_AGEMA_signal_4255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_56_U1_XOR1_U1 ( .A0_t (key_s0_t[120]), .A0_f (key_s0_f[120]), .A1_t (key_s1_t[120]), .A1_f (key_s1_f[120]), .B0_t (key_s0_t[56]), .B0_f (key_s0_f[56]), .B1_t (key_s1_t[56]), .B1_f (key_s1_f[56]), .Z0_t (Midori_rounds_MUXInst_mux_inst_56_U1_X), .Z0_f (new_AGEMA_signal_2769), .Z1_t (new_AGEMA_signal_2770), .Z1_f (new_AGEMA_signal_2771) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_56_U1_X), .B0_f (new_AGEMA_signal_2769), .B1_t (new_AGEMA_signal_2770), .B1_f (new_AGEMA_signal_2771), .Z0_t (Midori_rounds_MUXInst_mux_inst_56_U1_Y), .Z0_f (new_AGEMA_signal_3792), .Z1_t (new_AGEMA_signal_3793), .Z1_f (new_AGEMA_signal_3794) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_56_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_56_U1_Y), .A0_f (new_AGEMA_signal_3792), .A1_t (new_AGEMA_signal_3793), .A1_f (new_AGEMA_signal_3794), .B0_t (key_s0_t[120]), .B0_f (key_s0_f[120]), .B1_t (key_s1_t[120]), .B1_f (key_s1_f[120]), .Z0_t (Midori_rounds_SelectedKey[56]), .Z0_f (new_AGEMA_signal_4256), .Z1_t (new_AGEMA_signal_4257), .Z1_f (new_AGEMA_signal_4258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_57_U1_XOR1_U1 ( .A0_t (key_s0_t[121]), .A0_f (key_s0_f[121]), .A1_t (key_s1_t[121]), .A1_f (key_s1_f[121]), .B0_t (key_s0_t[57]), .B0_f (key_s0_f[57]), .B1_t (key_s1_t[57]), .B1_f (key_s1_f[57]), .Z0_t (Midori_rounds_MUXInst_mux_inst_57_U1_X), .Z0_f (new_AGEMA_signal_2772), .Z1_t (new_AGEMA_signal_2773), .Z1_f (new_AGEMA_signal_2774) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_57_U1_X), .B0_f (new_AGEMA_signal_2772), .B1_t (new_AGEMA_signal_2773), .B1_f (new_AGEMA_signal_2774), .Z0_t (Midori_rounds_MUXInst_mux_inst_57_U1_Y), .Z0_f (new_AGEMA_signal_3795), .Z1_t (new_AGEMA_signal_3796), .Z1_f (new_AGEMA_signal_3797) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_57_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_57_U1_Y), .A0_f (new_AGEMA_signal_3795), .A1_t (new_AGEMA_signal_3796), .A1_f (new_AGEMA_signal_3797), .B0_t (key_s0_t[121]), .B0_f (key_s0_f[121]), .B1_t (key_s1_t[121]), .B1_f (key_s1_f[121]), .Z0_t (Midori_rounds_SelectedKey[57]), .Z0_f (new_AGEMA_signal_4259), .Z1_t (new_AGEMA_signal_4260), .Z1_f (new_AGEMA_signal_4261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_58_U1_XOR1_U1 ( .A0_t (key_s0_t[122]), .A0_f (key_s0_f[122]), .A1_t (key_s1_t[122]), .A1_f (key_s1_f[122]), .B0_t (key_s0_t[58]), .B0_f (key_s0_f[58]), .B1_t (key_s1_t[58]), .B1_f (key_s1_f[58]), .Z0_t (Midori_rounds_MUXInst_mux_inst_58_U1_X), .Z0_f (new_AGEMA_signal_2775), .Z1_t (new_AGEMA_signal_2776), .Z1_f (new_AGEMA_signal_2777) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_58_U1_X), .B0_f (new_AGEMA_signal_2775), .B1_t (new_AGEMA_signal_2776), .B1_f (new_AGEMA_signal_2777), .Z0_t (Midori_rounds_MUXInst_mux_inst_58_U1_Y), .Z0_f (new_AGEMA_signal_3798), .Z1_t (new_AGEMA_signal_3799), .Z1_f (new_AGEMA_signal_3800) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_58_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_58_U1_Y), .A0_f (new_AGEMA_signal_3798), .A1_t (new_AGEMA_signal_3799), .A1_f (new_AGEMA_signal_3800), .B0_t (key_s0_t[122]), .B0_f (key_s0_f[122]), .B1_t (key_s1_t[122]), .B1_f (key_s1_f[122]), .Z0_t (Midori_rounds_SelectedKey[58]), .Z0_f (new_AGEMA_signal_4262), .Z1_t (new_AGEMA_signal_4263), .Z1_f (new_AGEMA_signal_4264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_59_U1_XOR1_U1 ( .A0_t (key_s0_t[123]), .A0_f (key_s0_f[123]), .A1_t (key_s1_t[123]), .A1_f (key_s1_f[123]), .B0_t (key_s0_t[59]), .B0_f (key_s0_f[59]), .B1_t (key_s1_t[59]), .B1_f (key_s1_f[59]), .Z0_t (Midori_rounds_MUXInst_mux_inst_59_U1_X), .Z0_f (new_AGEMA_signal_2778), .Z1_t (new_AGEMA_signal_2779), .Z1_f (new_AGEMA_signal_2780) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_59_U1_X), .B0_f (new_AGEMA_signal_2778), .B1_t (new_AGEMA_signal_2779), .B1_f (new_AGEMA_signal_2780), .Z0_t (Midori_rounds_MUXInst_mux_inst_59_U1_Y), .Z0_f (new_AGEMA_signal_3801), .Z1_t (new_AGEMA_signal_3802), .Z1_f (new_AGEMA_signal_3803) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_59_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_59_U1_Y), .A0_f (new_AGEMA_signal_3801), .A1_t (new_AGEMA_signal_3802), .A1_f (new_AGEMA_signal_3803), .B0_t (key_s0_t[123]), .B0_f (key_s0_f[123]), .B1_t (key_s1_t[123]), .B1_f (key_s1_f[123]), .Z0_t (Midori_rounds_SelectedKey[59]), .Z0_f (new_AGEMA_signal_4265), .Z1_t (new_AGEMA_signal_4266), .Z1_f (new_AGEMA_signal_4267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_60_U1_XOR1_U1 ( .A0_t (key_s0_t[124]), .A0_f (key_s0_f[124]), .A1_t (key_s1_t[124]), .A1_f (key_s1_f[124]), .B0_t (key_s0_t[60]), .B0_f (key_s0_f[60]), .B1_t (key_s1_t[60]), .B1_f (key_s1_f[60]), .Z0_t (Midori_rounds_MUXInst_mux_inst_60_U1_X), .Z0_f (new_AGEMA_signal_2781), .Z1_t (new_AGEMA_signal_2782), .Z1_f (new_AGEMA_signal_2783) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_60_U1_X), .B0_f (new_AGEMA_signal_2781), .B1_t (new_AGEMA_signal_2782), .B1_f (new_AGEMA_signal_2783), .Z0_t (Midori_rounds_MUXInst_mux_inst_60_U1_Y), .Z0_f (new_AGEMA_signal_3804), .Z1_t (new_AGEMA_signal_3805), .Z1_f (new_AGEMA_signal_3806) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_60_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_60_U1_Y), .A0_f (new_AGEMA_signal_3804), .A1_t (new_AGEMA_signal_3805), .A1_f (new_AGEMA_signal_3806), .B0_t (key_s0_t[124]), .B0_f (key_s0_f[124]), .B1_t (key_s1_t[124]), .B1_f (key_s1_f[124]), .Z0_t (Midori_rounds_SelectedKey[60]), .Z0_f (new_AGEMA_signal_4268), .Z1_t (new_AGEMA_signal_4269), .Z1_f (new_AGEMA_signal_4270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_61_U1_XOR1_U1 ( .A0_t (key_s0_t[125]), .A0_f (key_s0_f[125]), .A1_t (key_s1_t[125]), .A1_f (key_s1_f[125]), .B0_t (key_s0_t[61]), .B0_f (key_s0_f[61]), .B1_t (key_s1_t[61]), .B1_f (key_s1_f[61]), .Z0_t (Midori_rounds_MUXInst_mux_inst_61_U1_X), .Z0_f (new_AGEMA_signal_2784), .Z1_t (new_AGEMA_signal_2785), .Z1_f (new_AGEMA_signal_2786) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_61_U1_X), .B0_f (new_AGEMA_signal_2784), .B1_t (new_AGEMA_signal_2785), .B1_f (new_AGEMA_signal_2786), .Z0_t (Midori_rounds_MUXInst_mux_inst_61_U1_Y), .Z0_f (new_AGEMA_signal_3807), .Z1_t (new_AGEMA_signal_3808), .Z1_f (new_AGEMA_signal_3809) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_61_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_61_U1_Y), .A0_f (new_AGEMA_signal_3807), .A1_t (new_AGEMA_signal_3808), .A1_f (new_AGEMA_signal_3809), .B0_t (key_s0_t[125]), .B0_f (key_s0_f[125]), .B1_t (key_s1_t[125]), .B1_f (key_s1_f[125]), .Z0_t (Midori_rounds_SelectedKey[61]), .Z0_f (new_AGEMA_signal_4271), .Z1_t (new_AGEMA_signal_4272), .Z1_f (new_AGEMA_signal_4273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_62_U1_XOR1_U1 ( .A0_t (key_s0_t[126]), .A0_f (key_s0_f[126]), .A1_t (key_s1_t[126]), .A1_f (key_s1_f[126]), .B0_t (key_s0_t[62]), .B0_f (key_s0_f[62]), .B1_t (key_s1_t[62]), .B1_f (key_s1_f[62]), .Z0_t (Midori_rounds_MUXInst_mux_inst_62_U1_X), .Z0_f (new_AGEMA_signal_2787), .Z1_t (new_AGEMA_signal_2788), .Z1_f (new_AGEMA_signal_2789) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_62_U1_X), .B0_f (new_AGEMA_signal_2787), .B1_t (new_AGEMA_signal_2788), .B1_f (new_AGEMA_signal_2789), .Z0_t (Midori_rounds_MUXInst_mux_inst_62_U1_Y), .Z0_f (new_AGEMA_signal_3810), .Z1_t (new_AGEMA_signal_3811), .Z1_f (new_AGEMA_signal_3812) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_62_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_62_U1_Y), .A0_f (new_AGEMA_signal_3810), .A1_t (new_AGEMA_signal_3811), .A1_f (new_AGEMA_signal_3812), .B0_t (key_s0_t[126]), .B0_f (key_s0_f[126]), .B1_t (key_s1_t[126]), .B1_f (key_s1_f[126]), .Z0_t (Midori_rounds_SelectedKey[62]), .Z0_f (new_AGEMA_signal_4274), .Z1_t (new_AGEMA_signal_4275), .Z1_f (new_AGEMA_signal_4276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_63_U1_XOR1_U1 ( .A0_t (key_s0_t[127]), .A0_f (key_s0_f[127]), .A1_t (key_s1_t[127]), .A1_f (key_s1_f[127]), .B0_t (key_s0_t[63]), .B0_f (key_s0_f[63]), .B1_t (key_s1_t[63]), .B1_f (key_s1_f[63]), .Z0_t (Midori_rounds_MUXInst_mux_inst_63_U1_X), .Z0_f (new_AGEMA_signal_2790), .Z1_t (new_AGEMA_signal_2791), .Z1_f (new_AGEMA_signal_2792) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (round_Signal[0]), .A1_f (new_AGEMA_signal_2582), .B0_t (Midori_rounds_MUXInst_mux_inst_63_U1_X), .B0_f (new_AGEMA_signal_2790), .B1_t (new_AGEMA_signal_2791), .B1_f (new_AGEMA_signal_2792), .Z0_t (Midori_rounds_MUXInst_mux_inst_63_U1_Y), .Z0_f (new_AGEMA_signal_3813), .Z1_t (new_AGEMA_signal_3814), .Z1_f (new_AGEMA_signal_3815) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_63_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_63_U1_Y), .A0_f (new_AGEMA_signal_3813), .A1_t (new_AGEMA_signal_3814), .A1_f (new_AGEMA_signal_3815), .B0_t (key_s0_t[127]), .B0_f (key_s0_f[127]), .B1_t (key_s1_t[127]), .B1_f (key_s1_f[127]), .Z0_t (Midori_rounds_SelectedKey[63]), .Z0_f (new_AGEMA_signal_4277), .Z1_t (new_AGEMA_signal_4278), .Z1_f (new_AGEMA_signal_4279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[0]), .A0_f (new_AGEMA_signal_6980), .A1_t (new_AGEMA_signal_6981), .A1_f (new_AGEMA_signal_6982), .B0_t (Midori_add_Result_Start[0]), .B0_f (new_AGEMA_signal_3610), .B1_t (new_AGEMA_signal_3611), .B1_f (new_AGEMA_signal_3612), .Z0_t (Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_7010), .Z1_t (new_AGEMA_signal_7011), .Z1_f (new_AGEMA_signal_7012) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_X), .B0_f (new_AGEMA_signal_7010), .B1_t (new_AGEMA_signal_7011), .B1_f (new_AGEMA_signal_7012), .Z0_t (Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7058), .Z1_t (new_AGEMA_signal_7059), .Z1_f (new_AGEMA_signal_7060) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7058), .A1_t (new_AGEMA_signal_7059), .A1_f (new_AGEMA_signal_7060), .B0_t (Midori_rounds_round_Result[0]), .B0_f (new_AGEMA_signal_6980), .B1_t (new_AGEMA_signal_6981), .B1_f (new_AGEMA_signal_6982), .Z0_t (Midori_rounds_roundReg_out[0]), .Z0_f (new_AGEMA_signal_2805), .Z1_t (new_AGEMA_signal_2806), .Z1_f (new_AGEMA_signal_2807) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[1]), .A0_f (new_AGEMA_signal_6209), .A1_t (new_AGEMA_signal_6210), .A1_f (new_AGEMA_signal_6211), .B0_t (Midori_add_Result_Start[1]), .B0_f (new_AGEMA_signal_3604), .B1_t (new_AGEMA_signal_3605), .B1_f (new_AGEMA_signal_3606), .Z0_t (Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6353), .Z1_t (new_AGEMA_signal_6354), .Z1_f (new_AGEMA_signal_6355) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6353), .B1_t (new_AGEMA_signal_6354), .B1_f (new_AGEMA_signal_6355), .Z0_t (Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6533), .Z1_t (new_AGEMA_signal_6534), .Z1_f (new_AGEMA_signal_6535) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6533), .A1_t (new_AGEMA_signal_6534), .A1_f (new_AGEMA_signal_6535), .B0_t (Midori_rounds_round_Result[1]), .B0_f (new_AGEMA_signal_6209), .B1_t (new_AGEMA_signal_6210), .B1_f (new_AGEMA_signal_6211), .Z0_t (Midori_rounds_roundReg_out[1]), .Z0_f (new_AGEMA_signal_3816), .Z1_t (new_AGEMA_signal_3817), .Z1_f (new_AGEMA_signal_3818) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[2]), .A0_f (new_AGEMA_signal_6485), .A1_t (new_AGEMA_signal_6486), .A1_f (new_AGEMA_signal_6487), .B0_t (Midori_add_Result_Start[2]), .B0_f (new_AGEMA_signal_3598), .B1_t (new_AGEMA_signal_3599), .B1_f (new_AGEMA_signal_3600), .Z0_t (Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6536), .Z1_t (new_AGEMA_signal_6537), .Z1_f (new_AGEMA_signal_6538) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6536), .B1_t (new_AGEMA_signal_6537), .B1_f (new_AGEMA_signal_6538), .Z0_t (Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6707), .Z1_t (new_AGEMA_signal_6708), .Z1_f (new_AGEMA_signal_6709) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6707), .A1_t (new_AGEMA_signal_6708), .A1_f (new_AGEMA_signal_6709), .B0_t (Midori_rounds_round_Result[2]), .B0_f (new_AGEMA_signal_6485), .B1_t (new_AGEMA_signal_6486), .B1_f (new_AGEMA_signal_6487), .Z0_t (Midori_rounds_roundReg_out[2]), .Z0_f (new_AGEMA_signal_2796), .Z1_t (new_AGEMA_signal_2797), .Z1_f (new_AGEMA_signal_2798) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[3]), .A0_f (new_AGEMA_signal_6215), .A1_t (new_AGEMA_signal_6216), .A1_f (new_AGEMA_signal_6217), .B0_t (Midori_add_Result_Start[3]), .B0_f (new_AGEMA_signal_3592), .B1_t (new_AGEMA_signal_3593), .B1_f (new_AGEMA_signal_3594), .Z0_t (Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6356), .Z1_t (new_AGEMA_signal_6357), .Z1_f (new_AGEMA_signal_6358) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6356), .B1_t (new_AGEMA_signal_6357), .B1_f (new_AGEMA_signal_6358), .Z0_t (Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6539), .Z1_t (new_AGEMA_signal_6540), .Z1_f (new_AGEMA_signal_6541) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6539), .A1_t (new_AGEMA_signal_6540), .A1_f (new_AGEMA_signal_6541), .B0_t (Midori_rounds_round_Result[3]), .B0_f (new_AGEMA_signal_6215), .B1_t (new_AGEMA_signal_6216), .B1_f (new_AGEMA_signal_6217), .Z0_t (Midori_rounds_roundReg_out[3]), .Z0_f (new_AGEMA_signal_2793), .Z1_t (new_AGEMA_signal_2794), .Z1_f (new_AGEMA_signal_2795) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[4]), .A0_f (new_AGEMA_signal_6917), .A1_t (new_AGEMA_signal_6918), .A1_f (new_AGEMA_signal_6919), .B0_t (Midori_add_Result_Start[4]), .B0_f (new_AGEMA_signal_3586), .B1_t (new_AGEMA_signal_3587), .B1_f (new_AGEMA_signal_3588), .Z0_t (Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6962), .Z1_t (new_AGEMA_signal_6963), .Z1_f (new_AGEMA_signal_6964) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6962), .B1_t (new_AGEMA_signal_6963), .B1_f (new_AGEMA_signal_6964), .Z0_t (Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7013), .Z1_t (new_AGEMA_signal_7014), .Z1_f (new_AGEMA_signal_7015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7013), .A1_t (new_AGEMA_signal_7014), .A1_f (new_AGEMA_signal_7015), .B0_t (Midori_rounds_round_Result[4]), .B0_f (new_AGEMA_signal_6917), .B1_t (new_AGEMA_signal_6918), .B1_f (new_AGEMA_signal_6919), .Z0_t (Midori_rounds_roundReg_out[4]), .Z0_f (new_AGEMA_signal_2829), .Z1_t (new_AGEMA_signal_2830), .Z1_f (new_AGEMA_signal_2831) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[5]), .A0_f (new_AGEMA_signal_6218), .A1_t (new_AGEMA_signal_6219), .A1_f (new_AGEMA_signal_6220), .B0_t (Midori_add_Result_Start[5]), .B0_f (new_AGEMA_signal_3580), .B1_t (new_AGEMA_signal_3581), .B1_f (new_AGEMA_signal_3582), .Z0_t (Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6359), .Z1_t (new_AGEMA_signal_6360), .Z1_f (new_AGEMA_signal_6361) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6359), .B1_t (new_AGEMA_signal_6360), .B1_f (new_AGEMA_signal_6361), .Z0_t (Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6542), .Z1_t (new_AGEMA_signal_6543), .Z1_f (new_AGEMA_signal_6544) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6542), .A1_t (new_AGEMA_signal_6543), .A1_f (new_AGEMA_signal_6544), .B0_t (Midori_rounds_round_Result[5]), .B0_f (new_AGEMA_signal_6218), .B1_t (new_AGEMA_signal_6219), .B1_f (new_AGEMA_signal_6220), .Z0_t (Midori_rounds_roundReg_out[5]), .Z0_f (new_AGEMA_signal_3837), .Z1_t (new_AGEMA_signal_3838), .Z1_f (new_AGEMA_signal_3839) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[6]), .A0_f (new_AGEMA_signal_6488), .A1_t (new_AGEMA_signal_6489), .A1_f (new_AGEMA_signal_6490), .B0_t (Midori_add_Result_Start[6]), .B0_f (new_AGEMA_signal_3574), .B1_t (new_AGEMA_signal_3575), .B1_f (new_AGEMA_signal_3576), .Z0_t (Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6545), .Z1_t (new_AGEMA_signal_6546), .Z1_f (new_AGEMA_signal_6547) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6545), .B1_t (new_AGEMA_signal_6546), .B1_f (new_AGEMA_signal_6547), .Z0_t (Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6710), .Z1_t (new_AGEMA_signal_6711), .Z1_f (new_AGEMA_signal_6712) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6710), .A1_t (new_AGEMA_signal_6711), .A1_f (new_AGEMA_signal_6712), .B0_t (Midori_rounds_round_Result[6]), .B0_f (new_AGEMA_signal_6488), .B1_t (new_AGEMA_signal_6489), .B1_f (new_AGEMA_signal_6490), .Z0_t (Midori_rounds_roundReg_out[6]), .Z0_f (new_AGEMA_signal_2820), .Z1_t (new_AGEMA_signal_2821), .Z1_f (new_AGEMA_signal_2822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[7]), .A0_f (new_AGEMA_signal_6224), .A1_t (new_AGEMA_signal_6225), .A1_f (new_AGEMA_signal_6226), .B0_t (Midori_add_Result_Start[7]), .B0_f (new_AGEMA_signal_3568), .B1_t (new_AGEMA_signal_3569), .B1_f (new_AGEMA_signal_3570), .Z0_t (Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6362), .Z1_t (new_AGEMA_signal_6363), .Z1_f (new_AGEMA_signal_6364) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6362), .B1_t (new_AGEMA_signal_6363), .B1_f (new_AGEMA_signal_6364), .Z0_t (Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6548), .Z1_t (new_AGEMA_signal_6549), .Z1_f (new_AGEMA_signal_6550) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6548), .A1_t (new_AGEMA_signal_6549), .A1_f (new_AGEMA_signal_6550), .B0_t (Midori_rounds_round_Result[7]), .B0_f (new_AGEMA_signal_6224), .B1_t (new_AGEMA_signal_6225), .B1_f (new_AGEMA_signal_6226), .Z0_t (Midori_rounds_roundReg_out[7]), .Z0_f (new_AGEMA_signal_2823), .Z1_t (new_AGEMA_signal_2824), .Z1_f (new_AGEMA_signal_2825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[8]), .A0_f (new_AGEMA_signal_7052), .A1_t (new_AGEMA_signal_7053), .A1_f (new_AGEMA_signal_7054), .B0_t (Midori_add_Result_Start[8]), .B0_f (new_AGEMA_signal_3562), .B1_t (new_AGEMA_signal_3563), .B1_f (new_AGEMA_signal_3564), .Z0_t (Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_7061), .Z1_t (new_AGEMA_signal_7062), .Z1_f (new_AGEMA_signal_7063) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_X), .B0_f (new_AGEMA_signal_7061), .B1_t (new_AGEMA_signal_7062), .B1_f (new_AGEMA_signal_7063), .Z0_t (Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7088), .Z1_t (new_AGEMA_signal_7089), .Z1_f (new_AGEMA_signal_7090) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7088), .A1_t (new_AGEMA_signal_7089), .A1_f (new_AGEMA_signal_7090), .B0_t (Midori_rounds_round_Result[8]), .B0_f (new_AGEMA_signal_7052), .B1_t (new_AGEMA_signal_7053), .B1_f (new_AGEMA_signal_7054), .Z0_t (Midori_rounds_roundReg_out[8]), .Z0_f (new_AGEMA_signal_2856), .Z1_t (new_AGEMA_signal_2857), .Z1_f (new_AGEMA_signal_2858) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[9]), .A0_f (new_AGEMA_signal_6227), .A1_t (new_AGEMA_signal_6228), .A1_f (new_AGEMA_signal_6229), .B0_t (Midori_add_Result_Start[9]), .B0_f (new_AGEMA_signal_3556), .B1_t (new_AGEMA_signal_3557), .B1_f (new_AGEMA_signal_3558), .Z0_t (Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6365), .Z1_t (new_AGEMA_signal_6366), .Z1_f (new_AGEMA_signal_6367) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6365), .B1_t (new_AGEMA_signal_6366), .B1_f (new_AGEMA_signal_6367), .Z0_t (Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6551), .Z1_t (new_AGEMA_signal_6552), .Z1_f (new_AGEMA_signal_6553) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6551), .A1_t (new_AGEMA_signal_6552), .A1_f (new_AGEMA_signal_6553), .B0_t (Midori_rounds_round_Result[9]), .B0_f (new_AGEMA_signal_6227), .B1_t (new_AGEMA_signal_6228), .B1_f (new_AGEMA_signal_6229), .Z0_t (Midori_rounds_roundReg_out[9]), .Z0_f (new_AGEMA_signal_3852), .Z1_t (new_AGEMA_signal_3853), .Z1_f (new_AGEMA_signal_3854) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[10]), .A0_f (new_AGEMA_signal_6491), .A1_t (new_AGEMA_signal_6492), .A1_f (new_AGEMA_signal_6493), .B0_t (Midori_add_Result_Start[10]), .B0_f (new_AGEMA_signal_3550), .B1_t (new_AGEMA_signal_3551), .B1_f (new_AGEMA_signal_3552), .Z0_t (Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6554), .Z1_t (new_AGEMA_signal_6555), .Z1_f (new_AGEMA_signal_6556) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6554), .B1_t (new_AGEMA_signal_6555), .B1_f (new_AGEMA_signal_6556), .Z0_t (Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6713), .Z1_t (new_AGEMA_signal_6714), .Z1_f (new_AGEMA_signal_6715) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6713), .A1_t (new_AGEMA_signal_6714), .A1_f (new_AGEMA_signal_6715), .B0_t (Midori_rounds_round_Result[10]), .B0_f (new_AGEMA_signal_6491), .B1_t (new_AGEMA_signal_6492), .B1_f (new_AGEMA_signal_6493), .Z0_t (Midori_rounds_roundReg_out[10]), .Z0_f (new_AGEMA_signal_2847), .Z1_t (new_AGEMA_signal_2848), .Z1_f (new_AGEMA_signal_2849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[11]), .A0_f (new_AGEMA_signal_6233), .A1_t (new_AGEMA_signal_6234), .A1_f (new_AGEMA_signal_6235), .B0_t (Midori_add_Result_Start[11]), .B0_f (new_AGEMA_signal_3544), .B1_t (new_AGEMA_signal_3545), .B1_f (new_AGEMA_signal_3546), .Z0_t (Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6368), .Z1_t (new_AGEMA_signal_6369), .Z1_f (new_AGEMA_signal_6370) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6368), .B1_t (new_AGEMA_signal_6369), .B1_f (new_AGEMA_signal_6370), .Z0_t (Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6557), .Z1_t (new_AGEMA_signal_6558), .Z1_f (new_AGEMA_signal_6559) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6557), .A1_t (new_AGEMA_signal_6558), .A1_f (new_AGEMA_signal_6559), .B0_t (Midori_rounds_round_Result[11]), .B0_f (new_AGEMA_signal_6233), .B1_t (new_AGEMA_signal_6234), .B1_f (new_AGEMA_signal_6235), .Z0_t (Midori_rounds_roundReg_out[11]), .Z0_f (new_AGEMA_signal_2850), .Z1_t (new_AGEMA_signal_2851), .Z1_f (new_AGEMA_signal_2852) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[12]), .A0_f (new_AGEMA_signal_7055), .A1_t (new_AGEMA_signal_7056), .A1_f (new_AGEMA_signal_7057), .B0_t (Midori_add_Result_Start[12]), .B0_f (new_AGEMA_signal_3538), .B1_t (new_AGEMA_signal_3539), .B1_f (new_AGEMA_signal_3540), .Z0_t (Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_7064), .Z1_t (new_AGEMA_signal_7065), .Z1_f (new_AGEMA_signal_7066) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_X), .B0_f (new_AGEMA_signal_7064), .B1_t (new_AGEMA_signal_7065), .B1_f (new_AGEMA_signal_7066), .Z0_t (Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7091), .Z1_t (new_AGEMA_signal_7092), .Z1_f (new_AGEMA_signal_7093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7091), .A1_t (new_AGEMA_signal_7092), .A1_f (new_AGEMA_signal_7093), .B0_t (Midori_rounds_round_Result[12]), .B0_f (new_AGEMA_signal_7055), .B1_t (new_AGEMA_signal_7056), .B1_f (new_AGEMA_signal_7057), .Z0_t (Midori_rounds_roundReg_out[12]), .Z0_f (new_AGEMA_signal_2883), .Z1_t (new_AGEMA_signal_2884), .Z1_f (new_AGEMA_signal_2885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[13]), .A0_f (new_AGEMA_signal_6236), .A1_t (new_AGEMA_signal_6237), .A1_f (new_AGEMA_signal_6238), .B0_t (Midori_add_Result_Start[13]), .B0_f (new_AGEMA_signal_3532), .B1_t (new_AGEMA_signal_3533), .B1_f (new_AGEMA_signal_3534), .Z0_t (Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6371), .Z1_t (new_AGEMA_signal_6372), .Z1_f (new_AGEMA_signal_6373) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6371), .B1_t (new_AGEMA_signal_6372), .B1_f (new_AGEMA_signal_6373), .Z0_t (Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6560), .Z1_t (new_AGEMA_signal_6561), .Z1_f (new_AGEMA_signal_6562) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6560), .A1_t (new_AGEMA_signal_6561), .A1_f (new_AGEMA_signal_6562), .B0_t (Midori_rounds_round_Result[13]), .B0_f (new_AGEMA_signal_6236), .B1_t (new_AGEMA_signal_6237), .B1_f (new_AGEMA_signal_6238), .Z0_t (Midori_rounds_roundReg_out[13]), .Z0_f (new_AGEMA_signal_3867), .Z1_t (new_AGEMA_signal_3868), .Z1_f (new_AGEMA_signal_3869) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[14]), .A0_f (new_AGEMA_signal_6494), .A1_t (new_AGEMA_signal_6495), .A1_f (new_AGEMA_signal_6496), .B0_t (Midori_add_Result_Start[14]), .B0_f (new_AGEMA_signal_3526), .B1_t (new_AGEMA_signal_3527), .B1_f (new_AGEMA_signal_3528), .Z0_t (Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6563), .Z1_t (new_AGEMA_signal_6564), .Z1_f (new_AGEMA_signal_6565) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6563), .B1_t (new_AGEMA_signal_6564), .B1_f (new_AGEMA_signal_6565), .Z0_t (Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6716), .Z1_t (new_AGEMA_signal_6717), .Z1_f (new_AGEMA_signal_6718) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6716), .A1_t (new_AGEMA_signal_6717), .A1_f (new_AGEMA_signal_6718), .B0_t (Midori_rounds_round_Result[14]), .B0_f (new_AGEMA_signal_6494), .B1_t (new_AGEMA_signal_6495), .B1_f (new_AGEMA_signal_6496), .Z0_t (Midori_rounds_roundReg_out[14]), .Z0_f (new_AGEMA_signal_2874), .Z1_t (new_AGEMA_signal_2875), .Z1_f (new_AGEMA_signal_2876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[15]), .A0_f (new_AGEMA_signal_6242), .A1_t (new_AGEMA_signal_6243), .A1_f (new_AGEMA_signal_6244), .B0_t (Midori_add_Result_Start[15]), .B0_f (new_AGEMA_signal_3520), .B1_t (new_AGEMA_signal_3521), .B1_f (new_AGEMA_signal_3522), .Z0_t (Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6374), .Z1_t (new_AGEMA_signal_6375), .Z1_f (new_AGEMA_signal_6376) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6374), .B1_t (new_AGEMA_signal_6375), .B1_f (new_AGEMA_signal_6376), .Z0_t (Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6566), .Z1_t (new_AGEMA_signal_6567), .Z1_f (new_AGEMA_signal_6568) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6566), .A1_t (new_AGEMA_signal_6567), .A1_f (new_AGEMA_signal_6568), .B0_t (Midori_rounds_round_Result[15]), .B0_f (new_AGEMA_signal_6242), .B1_t (new_AGEMA_signal_6243), .B1_f (new_AGEMA_signal_6244), .Z0_t (Midori_rounds_roundReg_out[15]), .Z0_f (new_AGEMA_signal_2877), .Z1_t (new_AGEMA_signal_2878), .Z1_f (new_AGEMA_signal_2879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[16]), .A0_f (new_AGEMA_signal_6926), .A1_t (new_AGEMA_signal_6927), .A1_f (new_AGEMA_signal_6928), .B0_t (Midori_add_Result_Start[16]), .B0_f (new_AGEMA_signal_3514), .B1_t (new_AGEMA_signal_3515), .B1_f (new_AGEMA_signal_3516), .Z0_t (Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6965), .Z1_t (new_AGEMA_signal_6966), .Z1_f (new_AGEMA_signal_6967) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6965), .B1_t (new_AGEMA_signal_6966), .B1_f (new_AGEMA_signal_6967), .Z0_t (Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7016), .Z1_t (new_AGEMA_signal_7017), .Z1_f (new_AGEMA_signal_7018) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7016), .A1_t (new_AGEMA_signal_7017), .A1_f (new_AGEMA_signal_7018), .B0_t (Midori_rounds_round_Result[16]), .B0_f (new_AGEMA_signal_6926), .B1_t (new_AGEMA_signal_6927), .B1_f (new_AGEMA_signal_6928), .Z0_t (Midori_rounds_roundReg_out[16]), .Z0_f (new_AGEMA_signal_2910), .Z1_t (new_AGEMA_signal_2911), .Z1_f (new_AGEMA_signal_2912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[17]), .A0_f (new_AGEMA_signal_6245), .A1_t (new_AGEMA_signal_6246), .A1_f (new_AGEMA_signal_6247), .B0_t (Midori_add_Result_Start[17]), .B0_f (new_AGEMA_signal_3508), .B1_t (new_AGEMA_signal_3509), .B1_f (new_AGEMA_signal_3510), .Z0_t (Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6377), .Z1_t (new_AGEMA_signal_6378), .Z1_f (new_AGEMA_signal_6379) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6377), .B1_t (new_AGEMA_signal_6378), .B1_f (new_AGEMA_signal_6379), .Z0_t (Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6569), .Z1_t (new_AGEMA_signal_6570), .Z1_f (new_AGEMA_signal_6571) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6569), .A1_t (new_AGEMA_signal_6570), .A1_f (new_AGEMA_signal_6571), .B0_t (Midori_rounds_round_Result[17]), .B0_f (new_AGEMA_signal_6245), .B1_t (new_AGEMA_signal_6246), .B1_f (new_AGEMA_signal_6247), .Z0_t (Midori_rounds_roundReg_out[17]), .Z0_f (new_AGEMA_signal_3882), .Z1_t (new_AGEMA_signal_3883), .Z1_f (new_AGEMA_signal_3884) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[18]), .A0_f (new_AGEMA_signal_6497), .A1_t (new_AGEMA_signal_6498), .A1_f (new_AGEMA_signal_6499), .B0_t (Midori_add_Result_Start[18]), .B0_f (new_AGEMA_signal_3502), .B1_t (new_AGEMA_signal_3503), .B1_f (new_AGEMA_signal_3504), .Z0_t (Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6572), .Z1_t (new_AGEMA_signal_6573), .Z1_f (new_AGEMA_signal_6574) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6572), .B1_t (new_AGEMA_signal_6573), .B1_f (new_AGEMA_signal_6574), .Z0_t (Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6719), .Z1_t (new_AGEMA_signal_6720), .Z1_f (new_AGEMA_signal_6721) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6719), .A1_t (new_AGEMA_signal_6720), .A1_f (new_AGEMA_signal_6721), .B0_t (Midori_rounds_round_Result[18]), .B0_f (new_AGEMA_signal_6497), .B1_t (new_AGEMA_signal_6498), .B1_f (new_AGEMA_signal_6499), .Z0_t (Midori_rounds_roundReg_out[18]), .Z0_f (new_AGEMA_signal_2901), .Z1_t (new_AGEMA_signal_2902), .Z1_f (new_AGEMA_signal_2903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[19]), .A0_f (new_AGEMA_signal_6251), .A1_t (new_AGEMA_signal_6252), .A1_f (new_AGEMA_signal_6253), .B0_t (Midori_add_Result_Start[19]), .B0_f (new_AGEMA_signal_3496), .B1_t (new_AGEMA_signal_3497), .B1_f (new_AGEMA_signal_3498), .Z0_t (Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6380), .Z1_t (new_AGEMA_signal_6381), .Z1_f (new_AGEMA_signal_6382) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6380), .B1_t (new_AGEMA_signal_6381), .B1_f (new_AGEMA_signal_6382), .Z0_t (Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6575), .Z1_t (new_AGEMA_signal_6576), .Z1_f (new_AGEMA_signal_6577) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6575), .A1_t (new_AGEMA_signal_6576), .A1_f (new_AGEMA_signal_6577), .B0_t (Midori_rounds_round_Result[19]), .B0_f (new_AGEMA_signal_6251), .B1_t (new_AGEMA_signal_6252), .B1_f (new_AGEMA_signal_6253), .Z0_t (Midori_rounds_roundReg_out[19]), .Z0_f (new_AGEMA_signal_2904), .Z1_t (new_AGEMA_signal_2905), .Z1_f (new_AGEMA_signal_2906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[20]), .A0_f (new_AGEMA_signal_6929), .A1_t (new_AGEMA_signal_6930), .A1_f (new_AGEMA_signal_6931), .B0_t (Midori_add_Result_Start[20]), .B0_f (new_AGEMA_signal_3490), .B1_t (new_AGEMA_signal_3491), .B1_f (new_AGEMA_signal_3492), .Z0_t (Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6968), .Z1_t (new_AGEMA_signal_6969), .Z1_f (new_AGEMA_signal_6970) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6968), .B1_t (new_AGEMA_signal_6969), .B1_f (new_AGEMA_signal_6970), .Z0_t (Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7019), .Z1_t (new_AGEMA_signal_7020), .Z1_f (new_AGEMA_signal_7021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7019), .A1_t (new_AGEMA_signal_7020), .A1_f (new_AGEMA_signal_7021), .B0_t (Midori_rounds_round_Result[20]), .B0_f (new_AGEMA_signal_6929), .B1_t (new_AGEMA_signal_6930), .B1_f (new_AGEMA_signal_6931), .Z0_t (Midori_rounds_roundReg_out[20]), .Z0_f (new_AGEMA_signal_2937), .Z1_t (new_AGEMA_signal_2938), .Z1_f (new_AGEMA_signal_2939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[21]), .A0_f (new_AGEMA_signal_6254), .A1_t (new_AGEMA_signal_6255), .A1_f (new_AGEMA_signal_6256), .B0_t (Midori_add_Result_Start[21]), .B0_f (new_AGEMA_signal_3484), .B1_t (new_AGEMA_signal_3485), .B1_f (new_AGEMA_signal_3486), .Z0_t (Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6383), .Z1_t (new_AGEMA_signal_6384), .Z1_f (new_AGEMA_signal_6385) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6383), .B1_t (new_AGEMA_signal_6384), .B1_f (new_AGEMA_signal_6385), .Z0_t (Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6578), .Z1_t (new_AGEMA_signal_6579), .Z1_f (new_AGEMA_signal_6580) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6578), .A1_t (new_AGEMA_signal_6579), .A1_f (new_AGEMA_signal_6580), .B0_t (Midori_rounds_round_Result[21]), .B0_f (new_AGEMA_signal_6254), .B1_t (new_AGEMA_signal_6255), .B1_f (new_AGEMA_signal_6256), .Z0_t (Midori_rounds_roundReg_out[21]), .Z0_f (new_AGEMA_signal_3897), .Z1_t (new_AGEMA_signal_3898), .Z1_f (new_AGEMA_signal_3899) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[22]), .A0_f (new_AGEMA_signal_6500), .A1_t (new_AGEMA_signal_6501), .A1_f (new_AGEMA_signal_6502), .B0_t (Midori_add_Result_Start[22]), .B0_f (new_AGEMA_signal_3478), .B1_t (new_AGEMA_signal_3479), .B1_f (new_AGEMA_signal_3480), .Z0_t (Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6581), .Z1_t (new_AGEMA_signal_6582), .Z1_f (new_AGEMA_signal_6583) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6581), .B1_t (new_AGEMA_signal_6582), .B1_f (new_AGEMA_signal_6583), .Z0_t (Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6722), .Z1_t (new_AGEMA_signal_6723), .Z1_f (new_AGEMA_signal_6724) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6722), .A1_t (new_AGEMA_signal_6723), .A1_f (new_AGEMA_signal_6724), .B0_t (Midori_rounds_round_Result[22]), .B0_f (new_AGEMA_signal_6500), .B1_t (new_AGEMA_signal_6501), .B1_f (new_AGEMA_signal_6502), .Z0_t (Midori_rounds_roundReg_out[22]), .Z0_f (new_AGEMA_signal_2928), .Z1_t (new_AGEMA_signal_2929), .Z1_f (new_AGEMA_signal_2930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[23]), .A0_f (new_AGEMA_signal_6260), .A1_t (new_AGEMA_signal_6261), .A1_f (new_AGEMA_signal_6262), .B0_t (Midori_add_Result_Start[23]), .B0_f (new_AGEMA_signal_3472), .B1_t (new_AGEMA_signal_3473), .B1_f (new_AGEMA_signal_3474), .Z0_t (Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6386), .Z1_t (new_AGEMA_signal_6387), .Z1_f (new_AGEMA_signal_6388) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6386), .B1_t (new_AGEMA_signal_6387), .B1_f (new_AGEMA_signal_6388), .Z0_t (Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6584), .Z1_t (new_AGEMA_signal_6585), .Z1_f (new_AGEMA_signal_6586) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6584), .A1_t (new_AGEMA_signal_6585), .A1_f (new_AGEMA_signal_6586), .B0_t (Midori_rounds_round_Result[23]), .B0_f (new_AGEMA_signal_6260), .B1_t (new_AGEMA_signal_6261), .B1_f (new_AGEMA_signal_6262), .Z0_t (Midori_rounds_roundReg_out[23]), .Z0_f (new_AGEMA_signal_2931), .Z1_t (new_AGEMA_signal_2932), .Z1_f (new_AGEMA_signal_2933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[24]), .A0_f (new_AGEMA_signal_6989), .A1_t (new_AGEMA_signal_6990), .A1_f (new_AGEMA_signal_6991), .B0_t (Midori_add_Result_Start[24]), .B0_f (new_AGEMA_signal_3466), .B1_t (new_AGEMA_signal_3467), .B1_f (new_AGEMA_signal_3468), .Z0_t (Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_7022), .Z1_t (new_AGEMA_signal_7023), .Z1_f (new_AGEMA_signal_7024) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_X), .B0_f (new_AGEMA_signal_7022), .B1_t (new_AGEMA_signal_7023), .B1_f (new_AGEMA_signal_7024), .Z0_t (Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7067), .Z1_t (new_AGEMA_signal_7068), .Z1_f (new_AGEMA_signal_7069) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7067), .A1_t (new_AGEMA_signal_7068), .A1_f (new_AGEMA_signal_7069), .B0_t (Midori_rounds_round_Result[24]), .B0_f (new_AGEMA_signal_6989), .B1_t (new_AGEMA_signal_6990), .B1_f (new_AGEMA_signal_6991), .Z0_t (Midori_rounds_roundReg_out[24]), .Z0_f (new_AGEMA_signal_2964), .Z1_t (new_AGEMA_signal_2965), .Z1_f (new_AGEMA_signal_2966) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[25]), .A0_f (new_AGEMA_signal_6263), .A1_t (new_AGEMA_signal_6264), .A1_f (new_AGEMA_signal_6265), .B0_t (Midori_add_Result_Start[25]), .B0_f (new_AGEMA_signal_3460), .B1_t (new_AGEMA_signal_3461), .B1_f (new_AGEMA_signal_3462), .Z0_t (Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6389), .Z1_t (new_AGEMA_signal_6390), .Z1_f (new_AGEMA_signal_6391) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6389), .B1_t (new_AGEMA_signal_6390), .B1_f (new_AGEMA_signal_6391), .Z0_t (Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6587), .Z1_t (new_AGEMA_signal_6588), .Z1_f (new_AGEMA_signal_6589) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6587), .A1_t (new_AGEMA_signal_6588), .A1_f (new_AGEMA_signal_6589), .B0_t (Midori_rounds_round_Result[25]), .B0_f (new_AGEMA_signal_6263), .B1_t (new_AGEMA_signal_6264), .B1_f (new_AGEMA_signal_6265), .Z0_t (Midori_rounds_roundReg_out[25]), .Z0_f (new_AGEMA_signal_3912), .Z1_t (new_AGEMA_signal_3913), .Z1_f (new_AGEMA_signal_3914) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[26]), .A0_f (new_AGEMA_signal_6503), .A1_t (new_AGEMA_signal_6504), .A1_f (new_AGEMA_signal_6505), .B0_t (Midori_add_Result_Start[26]), .B0_f (new_AGEMA_signal_3454), .B1_t (new_AGEMA_signal_3455), .B1_f (new_AGEMA_signal_3456), .Z0_t (Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6590), .Z1_t (new_AGEMA_signal_6591), .Z1_f (new_AGEMA_signal_6592) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6590), .B1_t (new_AGEMA_signal_6591), .B1_f (new_AGEMA_signal_6592), .Z0_t (Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6725), .Z1_t (new_AGEMA_signal_6726), .Z1_f (new_AGEMA_signal_6727) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6725), .A1_t (new_AGEMA_signal_6726), .A1_f (new_AGEMA_signal_6727), .B0_t (Midori_rounds_round_Result[26]), .B0_f (new_AGEMA_signal_6503), .B1_t (new_AGEMA_signal_6504), .B1_f (new_AGEMA_signal_6505), .Z0_t (Midori_rounds_roundReg_out[26]), .Z0_f (new_AGEMA_signal_2955), .Z1_t (new_AGEMA_signal_2956), .Z1_f (new_AGEMA_signal_2957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[27]), .A0_f (new_AGEMA_signal_6269), .A1_t (new_AGEMA_signal_6270), .A1_f (new_AGEMA_signal_6271), .B0_t (Midori_add_Result_Start[27]), .B0_f (new_AGEMA_signal_3448), .B1_t (new_AGEMA_signal_3449), .B1_f (new_AGEMA_signal_3450), .Z0_t (Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6392), .Z1_t (new_AGEMA_signal_6393), .Z1_f (new_AGEMA_signal_6394) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6392), .B1_t (new_AGEMA_signal_6393), .B1_f (new_AGEMA_signal_6394), .Z0_t (Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6593), .Z1_t (new_AGEMA_signal_6594), .Z1_f (new_AGEMA_signal_6595) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6593), .A1_t (new_AGEMA_signal_6594), .A1_f (new_AGEMA_signal_6595), .B0_t (Midori_rounds_round_Result[27]), .B0_f (new_AGEMA_signal_6269), .B1_t (new_AGEMA_signal_6270), .B1_f (new_AGEMA_signal_6271), .Z0_t (Midori_rounds_roundReg_out[27]), .Z0_f (new_AGEMA_signal_2958), .Z1_t (new_AGEMA_signal_2959), .Z1_f (new_AGEMA_signal_2960) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[28]), .A0_f (new_AGEMA_signal_6992), .A1_t (new_AGEMA_signal_6993), .A1_f (new_AGEMA_signal_6994), .B0_t (Midori_add_Result_Start[28]), .B0_f (new_AGEMA_signal_3442), .B1_t (new_AGEMA_signal_3443), .B1_f (new_AGEMA_signal_3444), .Z0_t (Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_7025), .Z1_t (new_AGEMA_signal_7026), .Z1_f (new_AGEMA_signal_7027) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_X), .B0_f (new_AGEMA_signal_7025), .B1_t (new_AGEMA_signal_7026), .B1_f (new_AGEMA_signal_7027), .Z0_t (Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7070), .Z1_t (new_AGEMA_signal_7071), .Z1_f (new_AGEMA_signal_7072) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7070), .A1_t (new_AGEMA_signal_7071), .A1_f (new_AGEMA_signal_7072), .B0_t (Midori_rounds_round_Result[28]), .B0_f (new_AGEMA_signal_6992), .B1_t (new_AGEMA_signal_6993), .B1_f (new_AGEMA_signal_6994), .Z0_t (Midori_rounds_roundReg_out[28]), .Z0_f (new_AGEMA_signal_2994), .Z1_t (new_AGEMA_signal_2995), .Z1_f (new_AGEMA_signal_2996) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[29]), .A0_f (new_AGEMA_signal_6272), .A1_t (new_AGEMA_signal_6273), .A1_f (new_AGEMA_signal_6274), .B0_t (Midori_add_Result_Start[29]), .B0_f (new_AGEMA_signal_3436), .B1_t (new_AGEMA_signal_3437), .B1_f (new_AGEMA_signal_3438), .Z0_t (Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6395), .Z1_t (new_AGEMA_signal_6396), .Z1_f (new_AGEMA_signal_6397) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6395), .B1_t (new_AGEMA_signal_6396), .B1_f (new_AGEMA_signal_6397), .Z0_t (Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6596), .Z1_t (new_AGEMA_signal_6597), .Z1_f (new_AGEMA_signal_6598) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6596), .A1_t (new_AGEMA_signal_6597), .A1_f (new_AGEMA_signal_6598), .B0_t (Midori_rounds_round_Result[29]), .B0_f (new_AGEMA_signal_6272), .B1_t (new_AGEMA_signal_6273), .B1_f (new_AGEMA_signal_6274), .Z0_t (Midori_rounds_roundReg_out[29]), .Z0_f (new_AGEMA_signal_3921), .Z1_t (new_AGEMA_signal_3922), .Z1_f (new_AGEMA_signal_3923) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[30]), .A0_f (new_AGEMA_signal_6506), .A1_t (new_AGEMA_signal_6507), .A1_f (new_AGEMA_signal_6508), .B0_t (Midori_add_Result_Start[30]), .B0_f (new_AGEMA_signal_3430), .B1_t (new_AGEMA_signal_3431), .B1_f (new_AGEMA_signal_3432), .Z0_t (Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6599), .Z1_t (new_AGEMA_signal_6600), .Z1_f (new_AGEMA_signal_6601) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6599), .B1_t (new_AGEMA_signal_6600), .B1_f (new_AGEMA_signal_6601), .Z0_t (Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6728), .Z1_t (new_AGEMA_signal_6729), .Z1_f (new_AGEMA_signal_6730) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6728), .A1_t (new_AGEMA_signal_6729), .A1_f (new_AGEMA_signal_6730), .B0_t (Midori_rounds_round_Result[30]), .B0_f (new_AGEMA_signal_6506), .B1_t (new_AGEMA_signal_6507), .B1_f (new_AGEMA_signal_6508), .Z0_t (Midori_rounds_roundReg_out[30]), .Z0_f (new_AGEMA_signal_2985), .Z1_t (new_AGEMA_signal_2986), .Z1_f (new_AGEMA_signal_2987) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[31]), .A0_f (new_AGEMA_signal_6278), .A1_t (new_AGEMA_signal_6279), .A1_f (new_AGEMA_signal_6280), .B0_t (Midori_add_Result_Start[31]), .B0_f (new_AGEMA_signal_3424), .B1_t (new_AGEMA_signal_3425), .B1_f (new_AGEMA_signal_3426), .Z0_t (Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6398), .Z1_t (new_AGEMA_signal_6399), .Z1_f (new_AGEMA_signal_6400) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6398), .B1_t (new_AGEMA_signal_6399), .B1_f (new_AGEMA_signal_6400), .Z0_t (Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6602), .Z1_t (new_AGEMA_signal_6603), .Z1_f (new_AGEMA_signal_6604) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6602), .A1_t (new_AGEMA_signal_6603), .A1_f (new_AGEMA_signal_6604), .B0_t (Midori_rounds_round_Result[31]), .B0_f (new_AGEMA_signal_6278), .B1_t (new_AGEMA_signal_6279), .B1_f (new_AGEMA_signal_6280), .Z0_t (Midori_rounds_roundReg_out[31]), .Z0_f (new_AGEMA_signal_2982), .Z1_t (new_AGEMA_signal_2983), .Z1_f (new_AGEMA_signal_2984) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[32]), .A0_f (new_AGEMA_signal_6995), .A1_t (new_AGEMA_signal_6996), .A1_f (new_AGEMA_signal_6997), .B0_t (Midori_add_Result_Start[32]), .B0_f (new_AGEMA_signal_3418), .B1_t (new_AGEMA_signal_3419), .B1_f (new_AGEMA_signal_3420), .Z0_t (Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_7028), .Z1_t (new_AGEMA_signal_7029), .Z1_f (new_AGEMA_signal_7030) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_X), .B0_f (new_AGEMA_signal_7028), .B1_t (new_AGEMA_signal_7029), .B1_f (new_AGEMA_signal_7030), .Z0_t (Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7073), .Z1_t (new_AGEMA_signal_7074), .Z1_f (new_AGEMA_signal_7075) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7073), .A1_t (new_AGEMA_signal_7074), .A1_f (new_AGEMA_signal_7075), .B0_t (Midori_rounds_round_Result[32]), .B0_f (new_AGEMA_signal_6995), .B1_t (new_AGEMA_signal_6996), .B1_f (new_AGEMA_signal_6997), .Z0_t (Midori_rounds_roundReg_out[32]), .Z0_f (new_AGEMA_signal_3021), .Z1_t (new_AGEMA_signal_3022), .Z1_f (new_AGEMA_signal_3023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[33]), .A0_f (new_AGEMA_signal_6281), .A1_t (new_AGEMA_signal_6282), .A1_f (new_AGEMA_signal_6283), .B0_t (Midori_add_Result_Start[33]), .B0_f (new_AGEMA_signal_3412), .B1_t (new_AGEMA_signal_3413), .B1_f (new_AGEMA_signal_3414), .Z0_t (Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6401), .Z1_t (new_AGEMA_signal_6402), .Z1_f (new_AGEMA_signal_6403) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6401), .B1_t (new_AGEMA_signal_6402), .B1_f (new_AGEMA_signal_6403), .Z0_t (Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6605), .Z1_t (new_AGEMA_signal_6606), .Z1_f (new_AGEMA_signal_6607) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6605), .A1_t (new_AGEMA_signal_6606), .A1_f (new_AGEMA_signal_6607), .B0_t (Midori_rounds_round_Result[33]), .B0_f (new_AGEMA_signal_6281), .B1_t (new_AGEMA_signal_6282), .B1_f (new_AGEMA_signal_6283), .Z0_t (Midori_rounds_roundReg_out[33]), .Z0_f (new_AGEMA_signal_3936), .Z1_t (new_AGEMA_signal_3937), .Z1_f (new_AGEMA_signal_3938) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[34]), .A0_f (new_AGEMA_signal_6509), .A1_t (new_AGEMA_signal_6510), .A1_f (new_AGEMA_signal_6511), .B0_t (Midori_add_Result_Start[34]), .B0_f (new_AGEMA_signal_3406), .B1_t (new_AGEMA_signal_3407), .B1_f (new_AGEMA_signal_3408), .Z0_t (Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6608), .Z1_t (new_AGEMA_signal_6609), .Z1_f (new_AGEMA_signal_6610) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6608), .B1_t (new_AGEMA_signal_6609), .B1_f (new_AGEMA_signal_6610), .Z0_t (Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6731), .Z1_t (new_AGEMA_signal_6732), .Z1_f (new_AGEMA_signal_6733) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6731), .A1_t (new_AGEMA_signal_6732), .A1_f (new_AGEMA_signal_6733), .B0_t (Midori_rounds_round_Result[34]), .B0_f (new_AGEMA_signal_6509), .B1_t (new_AGEMA_signal_6510), .B1_f (new_AGEMA_signal_6511), .Z0_t (Midori_rounds_roundReg_out[34]), .Z0_f (new_AGEMA_signal_3012), .Z1_t (new_AGEMA_signal_3013), .Z1_f (new_AGEMA_signal_3014) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[35]), .A0_f (new_AGEMA_signal_6287), .A1_t (new_AGEMA_signal_6288), .A1_f (new_AGEMA_signal_6289), .B0_t (Midori_add_Result_Start[35]), .B0_f (new_AGEMA_signal_3400), .B1_t (new_AGEMA_signal_3401), .B1_f (new_AGEMA_signal_3402), .Z0_t (Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6404), .Z1_t (new_AGEMA_signal_6405), .Z1_f (new_AGEMA_signal_6406) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6404), .B1_t (new_AGEMA_signal_6405), .B1_f (new_AGEMA_signal_6406), .Z0_t (Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6611), .Z1_t (new_AGEMA_signal_6612), .Z1_f (new_AGEMA_signal_6613) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6611), .A1_t (new_AGEMA_signal_6612), .A1_f (new_AGEMA_signal_6613), .B0_t (Midori_rounds_round_Result[35]), .B0_f (new_AGEMA_signal_6287), .B1_t (new_AGEMA_signal_6288), .B1_f (new_AGEMA_signal_6289), .Z0_t (Midori_rounds_roundReg_out[35]), .Z0_f (new_AGEMA_signal_3009), .Z1_t (new_AGEMA_signal_3010), .Z1_f (new_AGEMA_signal_3011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[36]), .A0_f (new_AGEMA_signal_6941), .A1_t (new_AGEMA_signal_6942), .A1_f (new_AGEMA_signal_6943), .B0_t (Midori_add_Result_Start[36]), .B0_f (new_AGEMA_signal_3394), .B1_t (new_AGEMA_signal_3395), .B1_f (new_AGEMA_signal_3396), .Z0_t (Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6971), .Z1_t (new_AGEMA_signal_6972), .Z1_f (new_AGEMA_signal_6973) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6971), .B1_t (new_AGEMA_signal_6972), .B1_f (new_AGEMA_signal_6973), .Z0_t (Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7031), .Z1_t (new_AGEMA_signal_7032), .Z1_f (new_AGEMA_signal_7033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7031), .A1_t (new_AGEMA_signal_7032), .A1_f (new_AGEMA_signal_7033), .B0_t (Midori_rounds_round_Result[36]), .B0_f (new_AGEMA_signal_6941), .B1_t (new_AGEMA_signal_6942), .B1_f (new_AGEMA_signal_6943), .Z0_t (Midori_rounds_roundReg_out[36]), .Z0_f (new_AGEMA_signal_3048), .Z1_t (new_AGEMA_signal_3049), .Z1_f (new_AGEMA_signal_3050) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[37]), .A0_f (new_AGEMA_signal_6290), .A1_t (new_AGEMA_signal_6291), .A1_f (new_AGEMA_signal_6292), .B0_t (Midori_add_Result_Start[37]), .B0_f (new_AGEMA_signal_3388), .B1_t (new_AGEMA_signal_3389), .B1_f (new_AGEMA_signal_3390), .Z0_t (Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6407), .Z1_t (new_AGEMA_signal_6408), .Z1_f (new_AGEMA_signal_6409) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6407), .B1_t (new_AGEMA_signal_6408), .B1_f (new_AGEMA_signal_6409), .Z0_t (Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6614), .Z1_t (new_AGEMA_signal_6615), .Z1_f (new_AGEMA_signal_6616) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6614), .A1_t (new_AGEMA_signal_6615), .A1_f (new_AGEMA_signal_6616), .B0_t (Midori_rounds_round_Result[37]), .B0_f (new_AGEMA_signal_6290), .B1_t (new_AGEMA_signal_6291), .B1_f (new_AGEMA_signal_6292), .Z0_t (Midori_rounds_roundReg_out[37]), .Z0_f (new_AGEMA_signal_3951), .Z1_t (new_AGEMA_signal_3952), .Z1_f (new_AGEMA_signal_3953) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[38]), .A0_f (new_AGEMA_signal_6512), .A1_t (new_AGEMA_signal_6513), .A1_f (new_AGEMA_signal_6514), .B0_t (Midori_add_Result_Start[38]), .B0_f (new_AGEMA_signal_3382), .B1_t (new_AGEMA_signal_3383), .B1_f (new_AGEMA_signal_3384), .Z0_t (Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6617), .Z1_t (new_AGEMA_signal_6618), .Z1_f (new_AGEMA_signal_6619) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6617), .B1_t (new_AGEMA_signal_6618), .B1_f (new_AGEMA_signal_6619), .Z0_t (Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6734), .Z1_t (new_AGEMA_signal_6735), .Z1_f (new_AGEMA_signal_6736) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6734), .A1_t (new_AGEMA_signal_6735), .A1_f (new_AGEMA_signal_6736), .B0_t (Midori_rounds_round_Result[38]), .B0_f (new_AGEMA_signal_6512), .B1_t (new_AGEMA_signal_6513), .B1_f (new_AGEMA_signal_6514), .Z0_t (Midori_rounds_roundReg_out[38]), .Z0_f (new_AGEMA_signal_3039), .Z1_t (new_AGEMA_signal_3040), .Z1_f (new_AGEMA_signal_3041) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[39]), .A0_f (new_AGEMA_signal_6296), .A1_t (new_AGEMA_signal_6297), .A1_f (new_AGEMA_signal_6298), .B0_t (Midori_add_Result_Start[39]), .B0_f (new_AGEMA_signal_3376), .B1_t (new_AGEMA_signal_3377), .B1_f (new_AGEMA_signal_3378), .Z0_t (Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6410), .Z1_t (new_AGEMA_signal_6411), .Z1_f (new_AGEMA_signal_6412) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6410), .B1_t (new_AGEMA_signal_6411), .B1_f (new_AGEMA_signal_6412), .Z0_t (Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6620), .Z1_t (new_AGEMA_signal_6621), .Z1_f (new_AGEMA_signal_6622) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6620), .A1_t (new_AGEMA_signal_6621), .A1_f (new_AGEMA_signal_6622), .B0_t (Midori_rounds_round_Result[39]), .B0_f (new_AGEMA_signal_6296), .B1_t (new_AGEMA_signal_6297), .B1_f (new_AGEMA_signal_6298), .Z0_t (Midori_rounds_roundReg_out[39]), .Z0_f (new_AGEMA_signal_3036), .Z1_t (new_AGEMA_signal_3037), .Z1_f (new_AGEMA_signal_3038) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[40]), .A0_f (new_AGEMA_signal_6998), .A1_t (new_AGEMA_signal_6999), .A1_f (new_AGEMA_signal_7000), .B0_t (Midori_add_Result_Start[40]), .B0_f (new_AGEMA_signal_3370), .B1_t (new_AGEMA_signal_3371), .B1_f (new_AGEMA_signal_3372), .Z0_t (Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_7034), .Z1_t (new_AGEMA_signal_7035), .Z1_f (new_AGEMA_signal_7036) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_X), .B0_f (new_AGEMA_signal_7034), .B1_t (new_AGEMA_signal_7035), .B1_f (new_AGEMA_signal_7036), .Z0_t (Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7076), .Z1_t (new_AGEMA_signal_7077), .Z1_f (new_AGEMA_signal_7078) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7076), .A1_t (new_AGEMA_signal_7077), .A1_f (new_AGEMA_signal_7078), .B0_t (Midori_rounds_round_Result[40]), .B0_f (new_AGEMA_signal_6998), .B1_t (new_AGEMA_signal_6999), .B1_f (new_AGEMA_signal_7000), .Z0_t (Midori_rounds_roundReg_out[40]), .Z0_f (new_AGEMA_signal_3072), .Z1_t (new_AGEMA_signal_3073), .Z1_f (new_AGEMA_signal_3074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[41]), .A0_f (new_AGEMA_signal_6299), .A1_t (new_AGEMA_signal_6300), .A1_f (new_AGEMA_signal_6301), .B0_t (Midori_add_Result_Start[41]), .B0_f (new_AGEMA_signal_3364), .B1_t (new_AGEMA_signal_3365), .B1_f (new_AGEMA_signal_3366), .Z0_t (Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6413), .Z1_t (new_AGEMA_signal_6414), .Z1_f (new_AGEMA_signal_6415) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6413), .B1_t (new_AGEMA_signal_6414), .B1_f (new_AGEMA_signal_6415), .Z0_t (Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6623), .Z1_t (new_AGEMA_signal_6624), .Z1_f (new_AGEMA_signal_6625) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6623), .A1_t (new_AGEMA_signal_6624), .A1_f (new_AGEMA_signal_6625), .B0_t (Midori_rounds_round_Result[41]), .B0_f (new_AGEMA_signal_6299), .B1_t (new_AGEMA_signal_6300), .B1_f (new_AGEMA_signal_6301), .Z0_t (Midori_rounds_roundReg_out[41]), .Z0_f (new_AGEMA_signal_3972), .Z1_t (new_AGEMA_signal_3973), .Z1_f (new_AGEMA_signal_3974) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[42]), .A0_f (new_AGEMA_signal_6515), .A1_t (new_AGEMA_signal_6516), .A1_f (new_AGEMA_signal_6517), .B0_t (Midori_add_Result_Start[42]), .B0_f (new_AGEMA_signal_3358), .B1_t (new_AGEMA_signal_3359), .B1_f (new_AGEMA_signal_3360), .Z0_t (Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6626), .Z1_t (new_AGEMA_signal_6627), .Z1_f (new_AGEMA_signal_6628) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6626), .B1_t (new_AGEMA_signal_6627), .B1_f (new_AGEMA_signal_6628), .Z0_t (Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6737), .Z1_t (new_AGEMA_signal_6738), .Z1_f (new_AGEMA_signal_6739) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6737), .A1_t (new_AGEMA_signal_6738), .A1_f (new_AGEMA_signal_6739), .B0_t (Midori_rounds_round_Result[42]), .B0_f (new_AGEMA_signal_6515), .B1_t (new_AGEMA_signal_6516), .B1_f (new_AGEMA_signal_6517), .Z0_t (Midori_rounds_roundReg_out[42]), .Z0_f (new_AGEMA_signal_3063), .Z1_t (new_AGEMA_signal_3064), .Z1_f (new_AGEMA_signal_3065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[43]), .A0_f (new_AGEMA_signal_6305), .A1_t (new_AGEMA_signal_6306), .A1_f (new_AGEMA_signal_6307), .B0_t (Midori_add_Result_Start[43]), .B0_f (new_AGEMA_signal_3352), .B1_t (new_AGEMA_signal_3353), .B1_f (new_AGEMA_signal_3354), .Z0_t (Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6416), .Z1_t (new_AGEMA_signal_6417), .Z1_f (new_AGEMA_signal_6418) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6416), .B1_t (new_AGEMA_signal_6417), .B1_f (new_AGEMA_signal_6418), .Z0_t (Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6629), .Z1_t (new_AGEMA_signal_6630), .Z1_f (new_AGEMA_signal_6631) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6629), .A1_t (new_AGEMA_signal_6630), .A1_f (new_AGEMA_signal_6631), .B0_t (Midori_rounds_round_Result[43]), .B0_f (new_AGEMA_signal_6305), .B1_t (new_AGEMA_signal_6306), .B1_f (new_AGEMA_signal_6307), .Z0_t (Midori_rounds_roundReg_out[43]), .Z0_f (new_AGEMA_signal_3066), .Z1_t (new_AGEMA_signal_3067), .Z1_f (new_AGEMA_signal_3068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[44]), .A0_f (new_AGEMA_signal_7001), .A1_t (new_AGEMA_signal_7002), .A1_f (new_AGEMA_signal_7003), .B0_t (Midori_add_Result_Start[44]), .B0_f (new_AGEMA_signal_3346), .B1_t (new_AGEMA_signal_3347), .B1_f (new_AGEMA_signal_3348), .Z0_t (Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_7037), .Z1_t (new_AGEMA_signal_7038), .Z1_f (new_AGEMA_signal_7039) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_X), .B0_f (new_AGEMA_signal_7037), .B1_t (new_AGEMA_signal_7038), .B1_f (new_AGEMA_signal_7039), .Z0_t (Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7079), .Z1_t (new_AGEMA_signal_7080), .Z1_f (new_AGEMA_signal_7081) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7079), .A1_t (new_AGEMA_signal_7080), .A1_f (new_AGEMA_signal_7081), .B0_t (Midori_rounds_round_Result[44]), .B0_f (new_AGEMA_signal_7001), .B1_t (new_AGEMA_signal_7002), .B1_f (new_AGEMA_signal_7003), .Z0_t (Midori_rounds_roundReg_out[44]), .Z0_f (new_AGEMA_signal_3099), .Z1_t (new_AGEMA_signal_3100), .Z1_f (new_AGEMA_signal_3101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[45]), .A0_f (new_AGEMA_signal_6308), .A1_t (new_AGEMA_signal_6309), .A1_f (new_AGEMA_signal_6310), .B0_t (Midori_add_Result_Start[45]), .B0_f (new_AGEMA_signal_3340), .B1_t (new_AGEMA_signal_3341), .B1_f (new_AGEMA_signal_3342), .Z0_t (Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6419), .Z1_t (new_AGEMA_signal_6420), .Z1_f (new_AGEMA_signal_6421) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6419), .B1_t (new_AGEMA_signal_6420), .B1_f (new_AGEMA_signal_6421), .Z0_t (Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6632), .Z1_t (new_AGEMA_signal_6633), .Z1_f (new_AGEMA_signal_6634) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6632), .A1_t (new_AGEMA_signal_6633), .A1_f (new_AGEMA_signal_6634), .B0_t (Midori_rounds_round_Result[45]), .B0_f (new_AGEMA_signal_6308), .B1_t (new_AGEMA_signal_6309), .B1_f (new_AGEMA_signal_6310), .Z0_t (Midori_rounds_roundReg_out[45]), .Z0_f (new_AGEMA_signal_3987), .Z1_t (new_AGEMA_signal_3988), .Z1_f (new_AGEMA_signal_3989) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[46]), .A0_f (new_AGEMA_signal_6518), .A1_t (new_AGEMA_signal_6519), .A1_f (new_AGEMA_signal_6520), .B0_t (Midori_add_Result_Start[46]), .B0_f (new_AGEMA_signal_3334), .B1_t (new_AGEMA_signal_3335), .B1_f (new_AGEMA_signal_3336), .Z0_t (Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6635), .Z1_t (new_AGEMA_signal_6636), .Z1_f (new_AGEMA_signal_6637) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6635), .B1_t (new_AGEMA_signal_6636), .B1_f (new_AGEMA_signal_6637), .Z0_t (Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6740), .Z1_t (new_AGEMA_signal_6741), .Z1_f (new_AGEMA_signal_6742) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6740), .A1_t (new_AGEMA_signal_6741), .A1_f (new_AGEMA_signal_6742), .B0_t (Midori_rounds_round_Result[46]), .B0_f (new_AGEMA_signal_6518), .B1_t (new_AGEMA_signal_6519), .B1_f (new_AGEMA_signal_6520), .Z0_t (Midori_rounds_roundReg_out[46]), .Z0_f (new_AGEMA_signal_3090), .Z1_t (new_AGEMA_signal_3091), .Z1_f (new_AGEMA_signal_3092) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[47]), .A0_f (new_AGEMA_signal_6314), .A1_t (new_AGEMA_signal_6315), .A1_f (new_AGEMA_signal_6316), .B0_t (Midori_add_Result_Start[47]), .B0_f (new_AGEMA_signal_3328), .B1_t (new_AGEMA_signal_3329), .B1_f (new_AGEMA_signal_3330), .Z0_t (Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6422), .Z1_t (new_AGEMA_signal_6423), .Z1_f (new_AGEMA_signal_6424) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6422), .B1_t (new_AGEMA_signal_6423), .B1_f (new_AGEMA_signal_6424), .Z0_t (Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6638), .Z1_t (new_AGEMA_signal_6639), .Z1_f (new_AGEMA_signal_6640) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6638), .A1_t (new_AGEMA_signal_6639), .A1_f (new_AGEMA_signal_6640), .B0_t (Midori_rounds_round_Result[47]), .B0_f (new_AGEMA_signal_6314), .B1_t (new_AGEMA_signal_6315), .B1_f (new_AGEMA_signal_6316), .Z0_t (Midori_rounds_roundReg_out[47]), .Z0_f (new_AGEMA_signal_3093), .Z1_t (new_AGEMA_signal_3094), .Z1_f (new_AGEMA_signal_3095) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[48]), .A0_f (new_AGEMA_signal_6950), .A1_t (new_AGEMA_signal_6951), .A1_f (new_AGEMA_signal_6952), .B0_t (Midori_add_Result_Start[48]), .B0_f (new_AGEMA_signal_3322), .B1_t (new_AGEMA_signal_3323), .B1_f (new_AGEMA_signal_3324), .Z0_t (Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6974), .Z1_t (new_AGEMA_signal_6975), .Z1_f (new_AGEMA_signal_6976) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6974), .B1_t (new_AGEMA_signal_6975), .B1_f (new_AGEMA_signal_6976), .Z0_t (Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7040), .Z1_t (new_AGEMA_signal_7041), .Z1_f (new_AGEMA_signal_7042) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7040), .A1_t (new_AGEMA_signal_7041), .A1_f (new_AGEMA_signal_7042), .B0_t (Midori_rounds_round_Result[48]), .B0_f (new_AGEMA_signal_6950), .B1_t (new_AGEMA_signal_6951), .B1_f (new_AGEMA_signal_6952), .Z0_t (Midori_rounds_roundReg_out[48]), .Z0_f (new_AGEMA_signal_3126), .Z1_t (new_AGEMA_signal_3127), .Z1_f (new_AGEMA_signal_3128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[49]), .A0_f (new_AGEMA_signal_6317), .A1_t (new_AGEMA_signal_6318), .A1_f (new_AGEMA_signal_6319), .B0_t (Midori_add_Result_Start[49]), .B0_f (new_AGEMA_signal_3316), .B1_t (new_AGEMA_signal_3317), .B1_f (new_AGEMA_signal_3318), .Z0_t (Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6425), .Z1_t (new_AGEMA_signal_6426), .Z1_f (new_AGEMA_signal_6427) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6425), .B1_t (new_AGEMA_signal_6426), .B1_f (new_AGEMA_signal_6427), .Z0_t (Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6641), .Z1_t (new_AGEMA_signal_6642), .Z1_f (new_AGEMA_signal_6643) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6641), .A1_t (new_AGEMA_signal_6642), .A1_f (new_AGEMA_signal_6643), .B0_t (Midori_rounds_round_Result[49]), .B0_f (new_AGEMA_signal_6317), .B1_t (new_AGEMA_signal_6318), .B1_f (new_AGEMA_signal_6319), .Z0_t (Midori_rounds_roundReg_out[49]), .Z0_f (new_AGEMA_signal_4002), .Z1_t (new_AGEMA_signal_4003), .Z1_f (new_AGEMA_signal_4004) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[50]), .A0_f (new_AGEMA_signal_6521), .A1_t (new_AGEMA_signal_6522), .A1_f (new_AGEMA_signal_6523), .B0_t (Midori_add_Result_Start[50]), .B0_f (new_AGEMA_signal_3310), .B1_t (new_AGEMA_signal_3311), .B1_f (new_AGEMA_signal_3312), .Z0_t (Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6644), .Z1_t (new_AGEMA_signal_6645), .Z1_f (new_AGEMA_signal_6646) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6644), .B1_t (new_AGEMA_signal_6645), .B1_f (new_AGEMA_signal_6646), .Z0_t (Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6743), .Z1_t (new_AGEMA_signal_6744), .Z1_f (new_AGEMA_signal_6745) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6743), .A1_t (new_AGEMA_signal_6744), .A1_f (new_AGEMA_signal_6745), .B0_t (Midori_rounds_round_Result[50]), .B0_f (new_AGEMA_signal_6521), .B1_t (new_AGEMA_signal_6522), .B1_f (new_AGEMA_signal_6523), .Z0_t (Midori_rounds_roundReg_out[50]), .Z0_f (new_AGEMA_signal_3117), .Z1_t (new_AGEMA_signal_3118), .Z1_f (new_AGEMA_signal_3119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[51]), .A0_f (new_AGEMA_signal_6323), .A1_t (new_AGEMA_signal_6324), .A1_f (new_AGEMA_signal_6325), .B0_t (Midori_add_Result_Start[51]), .B0_f (new_AGEMA_signal_3304), .B1_t (new_AGEMA_signal_3305), .B1_f (new_AGEMA_signal_3306), .Z0_t (Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6428), .Z1_t (new_AGEMA_signal_6429), .Z1_f (new_AGEMA_signal_6430) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6428), .B1_t (new_AGEMA_signal_6429), .B1_f (new_AGEMA_signal_6430), .Z0_t (Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6647), .Z1_t (new_AGEMA_signal_6648), .Z1_f (new_AGEMA_signal_6649) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6647), .A1_t (new_AGEMA_signal_6648), .A1_f (new_AGEMA_signal_6649), .B0_t (Midori_rounds_round_Result[51]), .B0_f (new_AGEMA_signal_6323), .B1_t (new_AGEMA_signal_6324), .B1_f (new_AGEMA_signal_6325), .Z0_t (Midori_rounds_roundReg_out[51]), .Z0_f (new_AGEMA_signal_3120), .Z1_t (new_AGEMA_signal_3121), .Z1_f (new_AGEMA_signal_3122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[52]), .A0_f (new_AGEMA_signal_6953), .A1_t (new_AGEMA_signal_6954), .A1_f (new_AGEMA_signal_6955), .B0_t (Midori_add_Result_Start[52]), .B0_f (new_AGEMA_signal_3298), .B1_t (new_AGEMA_signal_3299), .B1_f (new_AGEMA_signal_3300), .Z0_t (Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6977), .Z1_t (new_AGEMA_signal_6978), .Z1_f (new_AGEMA_signal_6979) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6977), .B1_t (new_AGEMA_signal_6978), .B1_f (new_AGEMA_signal_6979), .Z0_t (Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7043), .Z1_t (new_AGEMA_signal_7044), .Z1_f (new_AGEMA_signal_7045) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7043), .A1_t (new_AGEMA_signal_7044), .A1_f (new_AGEMA_signal_7045), .B0_t (Midori_rounds_round_Result[52]), .B0_f (new_AGEMA_signal_6953), .B1_t (new_AGEMA_signal_6954), .B1_f (new_AGEMA_signal_6955), .Z0_t (Midori_rounds_roundReg_out[52]), .Z0_f (new_AGEMA_signal_3156), .Z1_t (new_AGEMA_signal_3157), .Z1_f (new_AGEMA_signal_3158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[53]), .A0_f (new_AGEMA_signal_6326), .A1_t (new_AGEMA_signal_6327), .A1_f (new_AGEMA_signal_6328), .B0_t (Midori_add_Result_Start[53]), .B0_f (new_AGEMA_signal_3292), .B1_t (new_AGEMA_signal_3293), .B1_f (new_AGEMA_signal_3294), .Z0_t (Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6431), .Z1_t (new_AGEMA_signal_6432), .Z1_f (new_AGEMA_signal_6433) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6431), .B1_t (new_AGEMA_signal_6432), .B1_f (new_AGEMA_signal_6433), .Z0_t (Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6650), .Z1_t (new_AGEMA_signal_6651), .Z1_f (new_AGEMA_signal_6652) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6650), .A1_t (new_AGEMA_signal_6651), .A1_f (new_AGEMA_signal_6652), .B0_t (Midori_rounds_round_Result[53]), .B0_f (new_AGEMA_signal_6326), .B1_t (new_AGEMA_signal_6327), .B1_f (new_AGEMA_signal_6328), .Z0_t (Midori_rounds_roundReg_out[53]), .Z0_f (new_AGEMA_signal_4011), .Z1_t (new_AGEMA_signal_4012), .Z1_f (new_AGEMA_signal_4013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[54]), .A0_f (new_AGEMA_signal_6524), .A1_t (new_AGEMA_signal_6525), .A1_f (new_AGEMA_signal_6526), .B0_t (Midori_add_Result_Start[54]), .B0_f (new_AGEMA_signal_3286), .B1_t (new_AGEMA_signal_3287), .B1_f (new_AGEMA_signal_3288), .Z0_t (Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6653), .Z1_t (new_AGEMA_signal_6654), .Z1_f (new_AGEMA_signal_6655) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6653), .B1_t (new_AGEMA_signal_6654), .B1_f (new_AGEMA_signal_6655), .Z0_t (Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6746), .Z1_t (new_AGEMA_signal_6747), .Z1_f (new_AGEMA_signal_6748) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6746), .A1_t (new_AGEMA_signal_6747), .A1_f (new_AGEMA_signal_6748), .B0_t (Midori_rounds_round_Result[54]), .B0_f (new_AGEMA_signal_6524), .B1_t (new_AGEMA_signal_6525), .B1_f (new_AGEMA_signal_6526), .Z0_t (Midori_rounds_roundReg_out[54]), .Z0_f (new_AGEMA_signal_3147), .Z1_t (new_AGEMA_signal_3148), .Z1_f (new_AGEMA_signal_3149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[55]), .A0_f (new_AGEMA_signal_6332), .A1_t (new_AGEMA_signal_6333), .A1_f (new_AGEMA_signal_6334), .B0_t (Midori_add_Result_Start[55]), .B0_f (new_AGEMA_signal_3280), .B1_t (new_AGEMA_signal_3281), .B1_f (new_AGEMA_signal_3282), .Z0_t (Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6434), .Z1_t (new_AGEMA_signal_6435), .Z1_f (new_AGEMA_signal_6436) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6434), .B1_t (new_AGEMA_signal_6435), .B1_f (new_AGEMA_signal_6436), .Z0_t (Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6656), .Z1_t (new_AGEMA_signal_6657), .Z1_f (new_AGEMA_signal_6658) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6656), .A1_t (new_AGEMA_signal_6657), .A1_f (new_AGEMA_signal_6658), .B0_t (Midori_rounds_round_Result[55]), .B0_f (new_AGEMA_signal_6332), .B1_t (new_AGEMA_signal_6333), .B1_f (new_AGEMA_signal_6334), .Z0_t (Midori_rounds_roundReg_out[55]), .Z0_f (new_AGEMA_signal_3144), .Z1_t (new_AGEMA_signal_3145), .Z1_f (new_AGEMA_signal_3146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[56]), .A0_f (new_AGEMA_signal_7004), .A1_t (new_AGEMA_signal_7005), .A1_f (new_AGEMA_signal_7006), .B0_t (Midori_add_Result_Start[56]), .B0_f (new_AGEMA_signal_3274), .B1_t (new_AGEMA_signal_3275), .B1_f (new_AGEMA_signal_3276), .Z0_t (Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_7046), .Z1_t (new_AGEMA_signal_7047), .Z1_f (new_AGEMA_signal_7048) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_X), .B0_f (new_AGEMA_signal_7046), .B1_t (new_AGEMA_signal_7047), .B1_f (new_AGEMA_signal_7048), .Z0_t (Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7082), .Z1_t (new_AGEMA_signal_7083), .Z1_f (new_AGEMA_signal_7084) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7082), .A1_t (new_AGEMA_signal_7083), .A1_f (new_AGEMA_signal_7084), .B0_t (Midori_rounds_round_Result[56]), .B0_f (new_AGEMA_signal_7004), .B1_t (new_AGEMA_signal_7005), .B1_f (new_AGEMA_signal_7006), .Z0_t (Midori_rounds_roundReg_out[56]), .Z0_f (new_AGEMA_signal_3183), .Z1_t (new_AGEMA_signal_3184), .Z1_f (new_AGEMA_signal_3185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[57]), .A0_f (new_AGEMA_signal_6335), .A1_t (new_AGEMA_signal_6336), .A1_f (new_AGEMA_signal_6337), .B0_t (Midori_add_Result_Start[57]), .B0_f (new_AGEMA_signal_3268), .B1_t (new_AGEMA_signal_3269), .B1_f (new_AGEMA_signal_3270), .Z0_t (Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6437), .Z1_t (new_AGEMA_signal_6438), .Z1_f (new_AGEMA_signal_6439) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6437), .B1_t (new_AGEMA_signal_6438), .B1_f (new_AGEMA_signal_6439), .Z0_t (Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6659), .Z1_t (new_AGEMA_signal_6660), .Z1_f (new_AGEMA_signal_6661) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6659), .A1_t (new_AGEMA_signal_6660), .A1_f (new_AGEMA_signal_6661), .B0_t (Midori_rounds_round_Result[57]), .B0_f (new_AGEMA_signal_6335), .B1_t (new_AGEMA_signal_6336), .B1_f (new_AGEMA_signal_6337), .Z0_t (Midori_rounds_roundReg_out[57]), .Z0_f (new_AGEMA_signal_4026), .Z1_t (new_AGEMA_signal_4027), .Z1_f (new_AGEMA_signal_4028) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[58]), .A0_f (new_AGEMA_signal_6527), .A1_t (new_AGEMA_signal_6528), .A1_f (new_AGEMA_signal_6529), .B0_t (Midori_add_Result_Start[58]), .B0_f (new_AGEMA_signal_3262), .B1_t (new_AGEMA_signal_3263), .B1_f (new_AGEMA_signal_3264), .Z0_t (Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6662), .Z1_t (new_AGEMA_signal_6663), .Z1_f (new_AGEMA_signal_6664) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6662), .B1_t (new_AGEMA_signal_6663), .B1_f (new_AGEMA_signal_6664), .Z0_t (Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6749), .Z1_t (new_AGEMA_signal_6750), .Z1_f (new_AGEMA_signal_6751) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6749), .A1_t (new_AGEMA_signal_6750), .A1_f (new_AGEMA_signal_6751), .B0_t (Midori_rounds_round_Result[58]), .B0_f (new_AGEMA_signal_6527), .B1_t (new_AGEMA_signal_6528), .B1_f (new_AGEMA_signal_6529), .Z0_t (Midori_rounds_roundReg_out[58]), .Z0_f (new_AGEMA_signal_3174), .Z1_t (new_AGEMA_signal_3175), .Z1_f (new_AGEMA_signal_3176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[59]), .A0_f (new_AGEMA_signal_6341), .A1_t (new_AGEMA_signal_6342), .A1_f (new_AGEMA_signal_6343), .B0_t (Midori_add_Result_Start[59]), .B0_f (new_AGEMA_signal_3256), .B1_t (new_AGEMA_signal_3257), .B1_f (new_AGEMA_signal_3258), .Z0_t (Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6440), .Z1_t (new_AGEMA_signal_6441), .Z1_f (new_AGEMA_signal_6442) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6440), .B1_t (new_AGEMA_signal_6441), .B1_f (new_AGEMA_signal_6442), .Z0_t (Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6665), .Z1_t (new_AGEMA_signal_6666), .Z1_f (new_AGEMA_signal_6667) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6665), .A1_t (new_AGEMA_signal_6666), .A1_f (new_AGEMA_signal_6667), .B0_t (Midori_rounds_round_Result[59]), .B0_f (new_AGEMA_signal_6341), .B1_t (new_AGEMA_signal_6342), .B1_f (new_AGEMA_signal_6343), .Z0_t (Midori_rounds_roundReg_out[59]), .Z0_f (new_AGEMA_signal_3171), .Z1_t (new_AGEMA_signal_3172), .Z1_f (new_AGEMA_signal_3173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[60]), .A0_f (new_AGEMA_signal_7007), .A1_t (new_AGEMA_signal_7008), .A1_f (new_AGEMA_signal_7009), .B0_t (Midori_add_Result_Start[60]), .B0_f (new_AGEMA_signal_3250), .B1_t (new_AGEMA_signal_3251), .B1_f (new_AGEMA_signal_3252), .Z0_t (Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_7049), .Z1_t (new_AGEMA_signal_7050), .Z1_f (new_AGEMA_signal_7051) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_X), .B0_f (new_AGEMA_signal_7049), .B1_t (new_AGEMA_signal_7050), .B1_f (new_AGEMA_signal_7051), .Z0_t (Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_7085), .Z1_t (new_AGEMA_signal_7086), .Z1_f (new_AGEMA_signal_7087) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_7085), .A1_t (new_AGEMA_signal_7086), .A1_f (new_AGEMA_signal_7087), .B0_t (Midori_rounds_round_Result[60]), .B0_f (new_AGEMA_signal_7007), .B1_t (new_AGEMA_signal_7008), .B1_f (new_AGEMA_signal_7009), .Z0_t (Midori_rounds_roundReg_out[60]), .Z0_f (new_AGEMA_signal_3207), .Z1_t (new_AGEMA_signal_3208), .Z1_f (new_AGEMA_signal_3209) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[61]), .A0_f (new_AGEMA_signal_6344), .A1_t (new_AGEMA_signal_6345), .A1_f (new_AGEMA_signal_6346), .B0_t (Midori_add_Result_Start[61]), .B0_f (new_AGEMA_signal_3244), .B1_t (new_AGEMA_signal_3245), .B1_f (new_AGEMA_signal_3246), .Z0_t (Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6443), .Z1_t (new_AGEMA_signal_6444), .Z1_f (new_AGEMA_signal_6445) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6443), .B1_t (new_AGEMA_signal_6444), .B1_f (new_AGEMA_signal_6445), .Z0_t (Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6668), .Z1_t (new_AGEMA_signal_6669), .Z1_f (new_AGEMA_signal_6670) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6668), .A1_t (new_AGEMA_signal_6669), .A1_f (new_AGEMA_signal_6670), .B0_t (Midori_rounds_round_Result[61]), .B0_f (new_AGEMA_signal_6344), .B1_t (new_AGEMA_signal_6345), .B1_f (new_AGEMA_signal_6346), .Z0_t (Midori_rounds_roundReg_out[61]), .Z0_f (new_AGEMA_signal_4047), .Z1_t (new_AGEMA_signal_4048), .Z1_f (new_AGEMA_signal_4049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[62]), .A0_f (new_AGEMA_signal_6530), .A1_t (new_AGEMA_signal_6531), .A1_f (new_AGEMA_signal_6532), .B0_t (Midori_add_Result_Start[62]), .B0_f (new_AGEMA_signal_3238), .B1_t (new_AGEMA_signal_3239), .B1_f (new_AGEMA_signal_3240), .Z0_t (Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6671), .Z1_t (new_AGEMA_signal_6672), .Z1_f (new_AGEMA_signal_6673) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6671), .B1_t (new_AGEMA_signal_6672), .B1_f (new_AGEMA_signal_6673), .Z0_t (Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6752), .Z1_t (new_AGEMA_signal_6753), .Z1_f (new_AGEMA_signal_6754) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6752), .A1_t (new_AGEMA_signal_6753), .A1_f (new_AGEMA_signal_6754), .B0_t (Midori_rounds_round_Result[62]), .B0_f (new_AGEMA_signal_6530), .B1_t (new_AGEMA_signal_6531), .B1_f (new_AGEMA_signal_6532), .Z0_t (Midori_rounds_roundReg_out[62]), .Z0_f (new_AGEMA_signal_3198), .Z1_t (new_AGEMA_signal_3199), .Z1_f (new_AGEMA_signal_3200) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[63]), .A0_f (new_AGEMA_signal_6350), .A1_t (new_AGEMA_signal_6351), .A1_f (new_AGEMA_signal_6352), .B0_t (Midori_add_Result_Start[63]), .B0_f (new_AGEMA_signal_3232), .B1_t (new_AGEMA_signal_3233), .B1_f (new_AGEMA_signal_3234), .Z0_t (Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_X), .Z0_f (new_AGEMA_signal_6446), .Z1_t (new_AGEMA_signal_6447), .Z1_f (new_AGEMA_signal_6448) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_X), .B0_f (new_AGEMA_signal_6446), .B1_t (new_AGEMA_signal_6447), .B1_f (new_AGEMA_signal_6448), .Z0_t (Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_Y), .Z0_f (new_AGEMA_signal_6674), .Z1_t (new_AGEMA_signal_6675), .Z1_f (new_AGEMA_signal_6676) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_Y), .A0_f (new_AGEMA_signal_6674), .A1_t (new_AGEMA_signal_6675), .A1_f (new_AGEMA_signal_6676), .B0_t (Midori_rounds_round_Result[63]), .B0_f (new_AGEMA_signal_6350), .B1_t (new_AGEMA_signal_6351), .B1_f (new_AGEMA_signal_6352), .Z0_t (Midori_rounds_roundReg_out[63]), .Z0_f (new_AGEMA_signal_3201), .Z1_t (new_AGEMA_signal_3202), .Z1_f (new_AGEMA_signal_3203) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n15), .A0_f (new_AGEMA_signal_2811), .A1_t (new_AGEMA_signal_2812), .A1_f (new_AGEMA_signal_2813), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n14), .B0_f (new_AGEMA_signal_3819), .B1_t (new_AGEMA_signal_3820), .B1_f (new_AGEMA_signal_3821), .Z0_t (Midori_rounds_SR_Result[51]), .Z0_f (new_AGEMA_signal_4280), .Z1_t (new_AGEMA_signal_4281), .Z1_f (new_AGEMA_signal_4282) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n13), .A0_f (new_AGEMA_signal_2817), .A1_t (new_AGEMA_signal_2818), .A1_f (new_AGEMA_signal_2819), .B0_t (Midori_rounds_roundReg_out[1]), .B0_f (new_AGEMA_signal_3816), .B1_t (new_AGEMA_signal_3817), .B1_f (new_AGEMA_signal_3818), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n14), .Z0_f (new_AGEMA_signal_3819), .Z1_t (new_AGEMA_signal_3820), .Z1_f (new_AGEMA_signal_3821) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n12), .A0_f (new_AGEMA_signal_2802), .A1_t (new_AGEMA_signal_2803), .A1_f (new_AGEMA_signal_2804), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n11), .B0_f (new_AGEMA_signal_3822), .B1_t (new_AGEMA_signal_3823), .B1_f (new_AGEMA_signal_3824), .Z0_t (Midori_rounds_SR_Result[49]), .Z0_f (new_AGEMA_signal_4283), .Z1_t (new_AGEMA_signal_4284), .Z1_f (new_AGEMA_signal_4285) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U16 ( .A0_t (Midori_rounds_roundReg_out[0]), .A0_f (new_AGEMA_signal_2805), .A1_t (new_AGEMA_signal_2806), .A1_f (new_AGEMA_signal_2807), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n10), .B0_f (new_AGEMA_signal_2799), .B1_t (new_AGEMA_signal_2800), .B1_f (new_AGEMA_signal_2801), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n11), .Z0_f (new_AGEMA_signal_3822), .Z1_t (new_AGEMA_signal_3823), .Z1_f (new_AGEMA_signal_3824) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U15 ( .A0_t (Midori_rounds_roundReg_out[3]), .A0_f (new_AGEMA_signal_2793), .A1_t (new_AGEMA_signal_2794), .A1_f (new_AGEMA_signal_2795), .B0_t (Midori_rounds_roundReg_out[2]), .B0_f (new_AGEMA_signal_2796), .B1_t (new_AGEMA_signal_2797), .B1_f (new_AGEMA_signal_2798), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n10), .Z0_f (new_AGEMA_signal_2799), .Z1_t (new_AGEMA_signal_2800), .Z1_f (new_AGEMA_signal_2801) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U14 ( .A0_t (Midori_rounds_roundReg_out[2]), .A0_f (new_AGEMA_signal_2796), .A1_t (new_AGEMA_signal_2797), .A1_f (new_AGEMA_signal_2798), .B0_t (Midori_rounds_roundReg_out[3]), .B0_f (new_AGEMA_signal_2793), .B1_t (new_AGEMA_signal_2794), .B1_f (new_AGEMA_signal_2795), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n12), .Z0_f (new_AGEMA_signal_2802), .Z1_t (new_AGEMA_signal_2803), .Z1_f (new_AGEMA_signal_2804) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n15), .A0_f (new_AGEMA_signal_2811), .A1_t (new_AGEMA_signal_2812), .A1_f (new_AGEMA_signal_2813), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n7), .B0_f (new_AGEMA_signal_4286), .B1_t (new_AGEMA_signal_4287), .B1_f (new_AGEMA_signal_4288), .Z0_t (Midori_rounds_SR_Result[50]), .Z0_f (new_AGEMA_signal_4682), .Z1_t (new_AGEMA_signal_4683), .Z1_f (new_AGEMA_signal_4684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n6), .A0_f (new_AGEMA_signal_3825), .A1_t (new_AGEMA_signal_3826), .A1_f (new_AGEMA_signal_3827), .B0_t (Midori_rounds_roundReg_out[1]), .B0_f (new_AGEMA_signal_3816), .B1_t (new_AGEMA_signal_3817), .B1_f (new_AGEMA_signal_3818), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n7), .Z0_f (new_AGEMA_signal_4286), .Z1_t (new_AGEMA_signal_4287), .Z1_f (new_AGEMA_signal_4288) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n5), .A0_f (new_AGEMA_signal_2808), .A1_t (new_AGEMA_signal_2809), .A1_f (new_AGEMA_signal_2810), .B0_t (Midori_rounds_roundReg_out[2]), .B0_f (new_AGEMA_signal_2796), .B1_t (new_AGEMA_signal_2797), .B1_f (new_AGEMA_signal_2798), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n6), .Z0_f (new_AGEMA_signal_3825), .Z1_t (new_AGEMA_signal_3826), .Z1_f (new_AGEMA_signal_3827) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U10 ( .A0_t (Midori_rounds_roundReg_out[0]), .A0_f (new_AGEMA_signal_2805), .A1_t (new_AGEMA_signal_2806), .A1_f (new_AGEMA_signal_2807), .B0_t (Midori_rounds_roundReg_out[3]), .B0_f (new_AGEMA_signal_2793), .B1_t (new_AGEMA_signal_2794), .B1_f (new_AGEMA_signal_2795), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n5), .Z0_f (new_AGEMA_signal_2808), .Z1_t (new_AGEMA_signal_2809), .Z1_f (new_AGEMA_signal_2810) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U9 ( .A0_t (Midori_rounds_roundReg_out[3]), .A0_f (new_AGEMA_signal_2793), .A1_t (new_AGEMA_signal_2794), .A1_f (new_AGEMA_signal_2795), .B0_t (Midori_rounds_roundReg_out[0]), .B0_f (new_AGEMA_signal_2805), .B1_t (new_AGEMA_signal_2806), .B1_f (new_AGEMA_signal_2807), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n15), .Z0_f (new_AGEMA_signal_2811), .Z1_t (new_AGEMA_signal_2812), .Z1_f (new_AGEMA_signal_2813) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n13), .A0_f (new_AGEMA_signal_2817), .A1_t (new_AGEMA_signal_2818), .A1_f (new_AGEMA_signal_2819), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n3), .B0_f (new_AGEMA_signal_4289), .B1_t (new_AGEMA_signal_4290), .B1_f (new_AGEMA_signal_4291), .Z0_t (Midori_rounds_SR_Result[48]), .Z0_f (new_AGEMA_signal_4685), .Z1_t (new_AGEMA_signal_4686), .Z1_f (new_AGEMA_signal_4687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U7 ( .A0_t (Midori_rounds_roundReg_out[1]), .A0_f (new_AGEMA_signal_3816), .A1_t (new_AGEMA_signal_3817), .A1_f (new_AGEMA_signal_3818), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n2), .B0_f (new_AGEMA_signal_3828), .B1_t (new_AGEMA_signal_3829), .B1_f (new_AGEMA_signal_3830), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n3), .Z0_f (new_AGEMA_signal_4289), .Z1_t (new_AGEMA_signal_4290), .Z1_f (new_AGEMA_signal_4291) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U6 ( .A0_t (Midori_rounds_roundReg_out[0]), .A0_f (new_AGEMA_signal_2805), .A1_t (new_AGEMA_signal_2806), .A1_f (new_AGEMA_signal_2807), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n1), .B0_f (new_AGEMA_signal_2814), .B1_t (new_AGEMA_signal_2815), .B1_f (new_AGEMA_signal_2816), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n2), .Z0_f (new_AGEMA_signal_3828), .Z1_t (new_AGEMA_signal_3829), .Z1_f (new_AGEMA_signal_3830) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U5 ( .A0_t (Midori_rounds_roundReg_out[2]), .A0_f (new_AGEMA_signal_2796), .A1_t (new_AGEMA_signal_2797), .A1_f (new_AGEMA_signal_2798), .B0_t (Midori_rounds_roundReg_out[3]), .B0_f (new_AGEMA_signal_2793), .B1_t (new_AGEMA_signal_2794), .B1_f (new_AGEMA_signal_2795), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n1), .Z0_f (new_AGEMA_signal_2814), .Z1_t (new_AGEMA_signal_2815), .Z1_f (new_AGEMA_signal_2816) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U3 ( .A0_t (Midori_rounds_roundReg_out[2]), .A0_f (new_AGEMA_signal_2796), .A1_t (new_AGEMA_signal_2797), .A1_f (new_AGEMA_signal_2798), .B0_t (Midori_rounds_roundReg_out[3]), .B0_f (new_AGEMA_signal_2793), .B1_t (new_AGEMA_signal_2794), .B1_f (new_AGEMA_signal_2795), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n13), .Z0_f (new_AGEMA_signal_2817), .Z1_t (new_AGEMA_signal_2818), .Z1_f (new_AGEMA_signal_2819) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n15), .A0_f (new_AGEMA_signal_4292), .A1_t (new_AGEMA_signal_4293), .A1_f (new_AGEMA_signal_4294), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n14), .B0_f (new_AGEMA_signal_2835), .B1_t (new_AGEMA_signal_2836), .B1_f (new_AGEMA_signal_2837), .Z0_t (Midori_rounds_SR_Result[44]), .Z0_f (new_AGEMA_signal_4688), .Z1_t (new_AGEMA_signal_4689), .Z1_f (new_AGEMA_signal_4690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U18 ( .A0_t (Midori_rounds_roundReg_out[5]), .A0_f (new_AGEMA_signal_3837), .A1_t (new_AGEMA_signal_3838), .A1_f (new_AGEMA_signal_3839), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n13), .B0_f (new_AGEMA_signal_3831), .B1_t (new_AGEMA_signal_3832), .B1_f (new_AGEMA_signal_3833), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n15), .Z0_f (new_AGEMA_signal_4292), .Z1_t (new_AGEMA_signal_4293), .Z1_f (new_AGEMA_signal_4294) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U17 ( .A0_t (Midori_rounds_roundReg_out[4]), .A0_f (new_AGEMA_signal_2829), .A1_t (new_AGEMA_signal_2830), .A1_f (new_AGEMA_signal_2831), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n11), .B0_f (new_AGEMA_signal_2826), .B1_t (new_AGEMA_signal_2827), .B1_f (new_AGEMA_signal_2828), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n13), .Z0_f (new_AGEMA_signal_3831), .Z1_t (new_AGEMA_signal_3832), .Z1_f (new_AGEMA_signal_3833) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U16 ( .A0_t (Midori_rounds_roundReg_out[6]), .A0_f (new_AGEMA_signal_2820), .A1_t (new_AGEMA_signal_2821), .A1_f (new_AGEMA_signal_2822), .B0_t (Midori_rounds_roundReg_out[7]), .B0_f (new_AGEMA_signal_2823), .B1_t (new_AGEMA_signal_2824), .B1_f (new_AGEMA_signal_2825), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n11), .Z0_f (new_AGEMA_signal_2826), .Z1_t (new_AGEMA_signal_2827), .Z1_f (new_AGEMA_signal_2828) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n10), .A0_f (new_AGEMA_signal_4295), .A1_t (new_AGEMA_signal_4296), .A1_f (new_AGEMA_signal_4297), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n9), .B0_f (new_AGEMA_signal_2838), .B1_t (new_AGEMA_signal_2839), .B1_f (new_AGEMA_signal_2840), .Z0_t (Midori_rounds_SR_Result[46]), .Z0_f (new_AGEMA_signal_4691), .Z1_t (new_AGEMA_signal_4692), .Z1_f (new_AGEMA_signal_4693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n8), .A0_f (new_AGEMA_signal_3834), .A1_t (new_AGEMA_signal_3835), .A1_f (new_AGEMA_signal_3836), .B0_t (Midori_rounds_roundReg_out[5]), .B0_f (new_AGEMA_signal_3837), .B1_t (new_AGEMA_signal_3838), .B1_f (new_AGEMA_signal_3839), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n10), .Z0_f (new_AGEMA_signal_4295), .Z1_t (new_AGEMA_signal_4296), .Z1_f (new_AGEMA_signal_4297) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n7), .A0_f (new_AGEMA_signal_2832), .A1_t (new_AGEMA_signal_2833), .A1_f (new_AGEMA_signal_2834), .B0_t (Midori_rounds_roundReg_out[6]), .B0_f (new_AGEMA_signal_2820), .B1_t (new_AGEMA_signal_2821), .B1_f (new_AGEMA_signal_2822), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n8), .Z0_f (new_AGEMA_signal_3834), .Z1_t (new_AGEMA_signal_3835), .Z1_f (new_AGEMA_signal_3836) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U12 ( .A0_t (Midori_rounds_roundReg_out[4]), .A0_f (new_AGEMA_signal_2829), .A1_t (new_AGEMA_signal_2830), .A1_f (new_AGEMA_signal_2831), .B0_t (Midori_rounds_roundReg_out[7]), .B0_f (new_AGEMA_signal_2823), .B1_t (new_AGEMA_signal_2824), .B1_f (new_AGEMA_signal_2825), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n7), .Z0_f (new_AGEMA_signal_2832), .Z1_t (new_AGEMA_signal_2833), .Z1_f (new_AGEMA_signal_2834) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n9), .A0_f (new_AGEMA_signal_2838), .A1_t (new_AGEMA_signal_2839), .A1_f (new_AGEMA_signal_2840), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n5), .B0_f (new_AGEMA_signal_3840), .B1_t (new_AGEMA_signal_3841), .B1_f (new_AGEMA_signal_3842), .Z0_t (Midori_rounds_SR_Result[47]), .Z0_f (new_AGEMA_signal_4298), .Z1_t (new_AGEMA_signal_4299), .Z1_f (new_AGEMA_signal_4300) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U10 ( .A0_t (Midori_rounds_roundReg_out[5]), .A0_f (new_AGEMA_signal_3837), .A1_t (new_AGEMA_signal_3838), .A1_f (new_AGEMA_signal_3839), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n14), .B0_f (new_AGEMA_signal_2835), .B1_t (new_AGEMA_signal_2836), .B1_f (new_AGEMA_signal_2837), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n5), .Z0_f (new_AGEMA_signal_3840), .Z1_t (new_AGEMA_signal_3841), .Z1_f (new_AGEMA_signal_3842) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U9 ( .A0_t (Midori_rounds_roundReg_out[6]), .A0_f (new_AGEMA_signal_2820), .A1_t (new_AGEMA_signal_2821), .A1_f (new_AGEMA_signal_2822), .B0_t (Midori_rounds_roundReg_out[7]), .B0_f (new_AGEMA_signal_2823), .B1_t (new_AGEMA_signal_2824), .B1_f (new_AGEMA_signal_2825), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n14), .Z0_f (new_AGEMA_signal_2835), .Z1_t (new_AGEMA_signal_2836), .Z1_f (new_AGEMA_signal_2837) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U8 ( .A0_t (Midori_rounds_roundReg_out[7]), .A0_f (new_AGEMA_signal_2823), .A1_t (new_AGEMA_signal_2824), .A1_f (new_AGEMA_signal_2825), .B0_t (Midori_rounds_roundReg_out[4]), .B0_f (new_AGEMA_signal_2829), .B1_t (new_AGEMA_signal_2830), .B1_f (new_AGEMA_signal_2831), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n9), .Z0_f (new_AGEMA_signal_2838), .Z1_t (new_AGEMA_signal_2839), .Z1_f (new_AGEMA_signal_2840) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n3), .A0_f (new_AGEMA_signal_2844), .A1_t (new_AGEMA_signal_2845), .A1_f (new_AGEMA_signal_2846), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n2), .B0_f (new_AGEMA_signal_3843), .B1_t (new_AGEMA_signal_3844), .B1_f (new_AGEMA_signal_3845), .Z0_t (Midori_rounds_SR_Result[45]), .Z0_f (new_AGEMA_signal_4301), .Z1_t (new_AGEMA_signal_4302), .Z1_f (new_AGEMA_signal_4303) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n1), .A0_f (new_AGEMA_signal_2841), .A1_t (new_AGEMA_signal_2842), .A1_f (new_AGEMA_signal_2843), .B0_t (Midori_rounds_roundReg_out[7]), .B0_f (new_AGEMA_signal_2823), .B1_t (new_AGEMA_signal_2824), .B1_f (new_AGEMA_signal_2825), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n2), .Z0_f (new_AGEMA_signal_3843), .Z1_t (new_AGEMA_signal_3844), .Z1_f (new_AGEMA_signal_3845) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U4 ( .A0_t (Midori_rounds_roundReg_out[6]), .A0_f (new_AGEMA_signal_2820), .A1_t (new_AGEMA_signal_2821), .A1_f (new_AGEMA_signal_2822), .B0_t (Midori_rounds_roundReg_out[4]), .B0_f (new_AGEMA_signal_2829), .B1_t (new_AGEMA_signal_2830), .B1_f (new_AGEMA_signal_2831), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n1), .Z0_f (new_AGEMA_signal_2841), .Z1_t (new_AGEMA_signal_2842), .Z1_f (new_AGEMA_signal_2843) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U1 ( .A0_t (Midori_rounds_roundReg_out[6]), .A0_f (new_AGEMA_signal_2820), .A1_t (new_AGEMA_signal_2821), .A1_f (new_AGEMA_signal_2822), .B0_t (Midori_rounds_roundReg_out[4]), .B0_f (new_AGEMA_signal_2829), .B1_t (new_AGEMA_signal_2830), .B1_f (new_AGEMA_signal_2831), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n3), .Z0_f (new_AGEMA_signal_2844), .Z1_t (new_AGEMA_signal_2845), .Z1_f (new_AGEMA_signal_2846) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n15), .A0_f (new_AGEMA_signal_4304), .A1_t (new_AGEMA_signal_4305), .A1_f (new_AGEMA_signal_4306), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n14), .B0_f (new_AGEMA_signal_2862), .B1_t (new_AGEMA_signal_2863), .B1_f (new_AGEMA_signal_2864), .Z0_t (Midori_rounds_SR_Result[8]), .Z0_f (new_AGEMA_signal_4694), .Z1_t (new_AGEMA_signal_4695), .Z1_f (new_AGEMA_signal_4696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U18 ( .A0_t (Midori_rounds_roundReg_out[9]), .A0_f (new_AGEMA_signal_3852), .A1_t (new_AGEMA_signal_3853), .A1_f (new_AGEMA_signal_3854), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n13), .B0_f (new_AGEMA_signal_3846), .B1_t (new_AGEMA_signal_3847), .B1_f (new_AGEMA_signal_3848), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n15), .Z0_f (new_AGEMA_signal_4304), .Z1_t (new_AGEMA_signal_4305), .Z1_f (new_AGEMA_signal_4306) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U17 ( .A0_t (Midori_rounds_roundReg_out[8]), .A0_f (new_AGEMA_signal_2856), .A1_t (new_AGEMA_signal_2857), .A1_f (new_AGEMA_signal_2858), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n11), .B0_f (new_AGEMA_signal_2853), .B1_t (new_AGEMA_signal_2854), .B1_f (new_AGEMA_signal_2855), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n13), .Z0_f (new_AGEMA_signal_3846), .Z1_t (new_AGEMA_signal_3847), .Z1_f (new_AGEMA_signal_3848) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U16 ( .A0_t (Midori_rounds_roundReg_out[10]), .A0_f (new_AGEMA_signal_2847), .A1_t (new_AGEMA_signal_2848), .A1_f (new_AGEMA_signal_2849), .B0_t (Midori_rounds_roundReg_out[11]), .B0_f (new_AGEMA_signal_2850), .B1_t (new_AGEMA_signal_2851), .B1_f (new_AGEMA_signal_2852), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n11), .Z0_f (new_AGEMA_signal_2853), .Z1_t (new_AGEMA_signal_2854), .Z1_f (new_AGEMA_signal_2855) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n10), .A0_f (new_AGEMA_signal_4307), .A1_t (new_AGEMA_signal_4308), .A1_f (new_AGEMA_signal_4309), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n9), .B0_f (new_AGEMA_signal_2865), .B1_t (new_AGEMA_signal_2866), .B1_f (new_AGEMA_signal_2867), .Z0_t (Midori_rounds_SR_Result[10]), .Z0_f (new_AGEMA_signal_4697), .Z1_t (new_AGEMA_signal_4698), .Z1_f (new_AGEMA_signal_4699) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n8), .A0_f (new_AGEMA_signal_3849), .A1_t (new_AGEMA_signal_3850), .A1_f (new_AGEMA_signal_3851), .B0_t (Midori_rounds_roundReg_out[9]), .B0_f (new_AGEMA_signal_3852), .B1_t (new_AGEMA_signal_3853), .B1_f (new_AGEMA_signal_3854), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n10), .Z0_f (new_AGEMA_signal_4307), .Z1_t (new_AGEMA_signal_4308), .Z1_f (new_AGEMA_signal_4309) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n7), .A0_f (new_AGEMA_signal_2859), .A1_t (new_AGEMA_signal_2860), .A1_f (new_AGEMA_signal_2861), .B0_t (Midori_rounds_roundReg_out[10]), .B0_f (new_AGEMA_signal_2847), .B1_t (new_AGEMA_signal_2848), .B1_f (new_AGEMA_signal_2849), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n8), .Z0_f (new_AGEMA_signal_3849), .Z1_t (new_AGEMA_signal_3850), .Z1_f (new_AGEMA_signal_3851) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U12 ( .A0_t (Midori_rounds_roundReg_out[8]), .A0_f (new_AGEMA_signal_2856), .A1_t (new_AGEMA_signal_2857), .A1_f (new_AGEMA_signal_2858), .B0_t (Midori_rounds_roundReg_out[11]), .B0_f (new_AGEMA_signal_2850), .B1_t (new_AGEMA_signal_2851), .B1_f (new_AGEMA_signal_2852), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n7), .Z0_f (new_AGEMA_signal_2859), .Z1_t (new_AGEMA_signal_2860), .Z1_f (new_AGEMA_signal_2861) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n9), .A0_f (new_AGEMA_signal_2865), .A1_t (new_AGEMA_signal_2866), .A1_f (new_AGEMA_signal_2867), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n5), .B0_f (new_AGEMA_signal_3855), .B1_t (new_AGEMA_signal_3856), .B1_f (new_AGEMA_signal_3857), .Z0_t (Midori_rounds_SR_Result[11]), .Z0_f (new_AGEMA_signal_4310), .Z1_t (new_AGEMA_signal_4311), .Z1_f (new_AGEMA_signal_4312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U10 ( .A0_t (Midori_rounds_roundReg_out[9]), .A0_f (new_AGEMA_signal_3852), .A1_t (new_AGEMA_signal_3853), .A1_f (new_AGEMA_signal_3854), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n14), .B0_f (new_AGEMA_signal_2862), .B1_t (new_AGEMA_signal_2863), .B1_f (new_AGEMA_signal_2864), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n5), .Z0_f (new_AGEMA_signal_3855), .Z1_t (new_AGEMA_signal_3856), .Z1_f (new_AGEMA_signal_3857) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U9 ( .A0_t (Midori_rounds_roundReg_out[10]), .A0_f (new_AGEMA_signal_2847), .A1_t (new_AGEMA_signal_2848), .A1_f (new_AGEMA_signal_2849), .B0_t (Midori_rounds_roundReg_out[11]), .B0_f (new_AGEMA_signal_2850), .B1_t (new_AGEMA_signal_2851), .B1_f (new_AGEMA_signal_2852), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n14), .Z0_f (new_AGEMA_signal_2862), .Z1_t (new_AGEMA_signal_2863), .Z1_f (new_AGEMA_signal_2864) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U8 ( .A0_t (Midori_rounds_roundReg_out[11]), .A0_f (new_AGEMA_signal_2850), .A1_t (new_AGEMA_signal_2851), .A1_f (new_AGEMA_signal_2852), .B0_t (Midori_rounds_roundReg_out[8]), .B0_f (new_AGEMA_signal_2856), .B1_t (new_AGEMA_signal_2857), .B1_f (new_AGEMA_signal_2858), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n9), .Z0_f (new_AGEMA_signal_2865), .Z1_t (new_AGEMA_signal_2866), .Z1_f (new_AGEMA_signal_2867) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n3), .A0_f (new_AGEMA_signal_2871), .A1_t (new_AGEMA_signal_2872), .A1_f (new_AGEMA_signal_2873), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n2), .B0_f (new_AGEMA_signal_3858), .B1_t (new_AGEMA_signal_3859), .B1_f (new_AGEMA_signal_3860), .Z0_t (Midori_rounds_SR_Result[9]), .Z0_f (new_AGEMA_signal_4313), .Z1_t (new_AGEMA_signal_4314), .Z1_f (new_AGEMA_signal_4315) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n1), .A0_f (new_AGEMA_signal_2868), .A1_t (new_AGEMA_signal_2869), .A1_f (new_AGEMA_signal_2870), .B0_t (Midori_rounds_roundReg_out[11]), .B0_f (new_AGEMA_signal_2850), .B1_t (new_AGEMA_signal_2851), .B1_f (new_AGEMA_signal_2852), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n2), .Z0_f (new_AGEMA_signal_3858), .Z1_t (new_AGEMA_signal_3859), .Z1_f (new_AGEMA_signal_3860) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U4 ( .A0_t (Midori_rounds_roundReg_out[10]), .A0_f (new_AGEMA_signal_2847), .A1_t (new_AGEMA_signal_2848), .A1_f (new_AGEMA_signal_2849), .B0_t (Midori_rounds_roundReg_out[8]), .B0_f (new_AGEMA_signal_2856), .B1_t (new_AGEMA_signal_2857), .B1_f (new_AGEMA_signal_2858), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n1), .Z0_f (new_AGEMA_signal_2868), .Z1_t (new_AGEMA_signal_2869), .Z1_f (new_AGEMA_signal_2870) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U1 ( .A0_t (Midori_rounds_roundReg_out[10]), .A0_f (new_AGEMA_signal_2847), .A1_t (new_AGEMA_signal_2848), .A1_f (new_AGEMA_signal_2849), .B0_t (Midori_rounds_roundReg_out[8]), .B0_f (new_AGEMA_signal_2856), .B1_t (new_AGEMA_signal_2857), .B1_f (new_AGEMA_signal_2858), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n3), .Z0_f (new_AGEMA_signal_2871), .Z1_t (new_AGEMA_signal_2872), .Z1_f (new_AGEMA_signal_2873) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n15), .A0_f (new_AGEMA_signal_4316), .A1_t (new_AGEMA_signal_4317), .A1_f (new_AGEMA_signal_4318), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n14), .B0_f (new_AGEMA_signal_2889), .B1_t (new_AGEMA_signal_2890), .B1_f (new_AGEMA_signal_2891), .Z0_t (Midori_rounds_SR_Result[20]), .Z0_f (new_AGEMA_signal_4700), .Z1_t (new_AGEMA_signal_4701), .Z1_f (new_AGEMA_signal_4702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U18 ( .A0_t (Midori_rounds_roundReg_out[13]), .A0_f (new_AGEMA_signal_3867), .A1_t (new_AGEMA_signal_3868), .A1_f (new_AGEMA_signal_3869), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n13), .B0_f (new_AGEMA_signal_3861), .B1_t (new_AGEMA_signal_3862), .B1_f (new_AGEMA_signal_3863), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n15), .Z0_f (new_AGEMA_signal_4316), .Z1_t (new_AGEMA_signal_4317), .Z1_f (new_AGEMA_signal_4318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U17 ( .A0_t (Midori_rounds_roundReg_out[12]), .A0_f (new_AGEMA_signal_2883), .A1_t (new_AGEMA_signal_2884), .A1_f (new_AGEMA_signal_2885), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n11), .B0_f (new_AGEMA_signal_2880), .B1_t (new_AGEMA_signal_2881), .B1_f (new_AGEMA_signal_2882), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n13), .Z0_f (new_AGEMA_signal_3861), .Z1_t (new_AGEMA_signal_3862), .Z1_f (new_AGEMA_signal_3863) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U16 ( .A0_t (Midori_rounds_roundReg_out[14]), .A0_f (new_AGEMA_signal_2874), .A1_t (new_AGEMA_signal_2875), .A1_f (new_AGEMA_signal_2876), .B0_t (Midori_rounds_roundReg_out[15]), .B0_f (new_AGEMA_signal_2877), .B1_t (new_AGEMA_signal_2878), .B1_f (new_AGEMA_signal_2879), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n11), .Z0_f (new_AGEMA_signal_2880), .Z1_t (new_AGEMA_signal_2881), .Z1_f (new_AGEMA_signal_2882) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n10), .A0_f (new_AGEMA_signal_4319), .A1_t (new_AGEMA_signal_4320), .A1_f (new_AGEMA_signal_4321), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n9), .B0_f (new_AGEMA_signal_2892), .B1_t (new_AGEMA_signal_2893), .B1_f (new_AGEMA_signal_2894), .Z0_t (Midori_rounds_SR_Result[22]), .Z0_f (new_AGEMA_signal_4703), .Z1_t (new_AGEMA_signal_4704), .Z1_f (new_AGEMA_signal_4705) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n8), .A0_f (new_AGEMA_signal_3864), .A1_t (new_AGEMA_signal_3865), .A1_f (new_AGEMA_signal_3866), .B0_t (Midori_rounds_roundReg_out[13]), .B0_f (new_AGEMA_signal_3867), .B1_t (new_AGEMA_signal_3868), .B1_f (new_AGEMA_signal_3869), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n10), .Z0_f (new_AGEMA_signal_4319), .Z1_t (new_AGEMA_signal_4320), .Z1_f (new_AGEMA_signal_4321) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n7), .A0_f (new_AGEMA_signal_2886), .A1_t (new_AGEMA_signal_2887), .A1_f (new_AGEMA_signal_2888), .B0_t (Midori_rounds_roundReg_out[14]), .B0_f (new_AGEMA_signal_2874), .B1_t (new_AGEMA_signal_2875), .B1_f (new_AGEMA_signal_2876), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n8), .Z0_f (new_AGEMA_signal_3864), .Z1_t (new_AGEMA_signal_3865), .Z1_f (new_AGEMA_signal_3866) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U12 ( .A0_t (Midori_rounds_roundReg_out[12]), .A0_f (new_AGEMA_signal_2883), .A1_t (new_AGEMA_signal_2884), .A1_f (new_AGEMA_signal_2885), .B0_t (Midori_rounds_roundReg_out[15]), .B0_f (new_AGEMA_signal_2877), .B1_t (new_AGEMA_signal_2878), .B1_f (new_AGEMA_signal_2879), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n7), .Z0_f (new_AGEMA_signal_2886), .Z1_t (new_AGEMA_signal_2887), .Z1_f (new_AGEMA_signal_2888) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n9), .A0_f (new_AGEMA_signal_2892), .A1_t (new_AGEMA_signal_2893), .A1_f (new_AGEMA_signal_2894), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n5), .B0_f (new_AGEMA_signal_3870), .B1_t (new_AGEMA_signal_3871), .B1_f (new_AGEMA_signal_3872), .Z0_t (Midori_rounds_SR_Result[23]), .Z0_f (new_AGEMA_signal_4322), .Z1_t (new_AGEMA_signal_4323), .Z1_f (new_AGEMA_signal_4324) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U10 ( .A0_t (Midori_rounds_roundReg_out[13]), .A0_f (new_AGEMA_signal_3867), .A1_t (new_AGEMA_signal_3868), .A1_f (new_AGEMA_signal_3869), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n14), .B0_f (new_AGEMA_signal_2889), .B1_t (new_AGEMA_signal_2890), .B1_f (new_AGEMA_signal_2891), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n5), .Z0_f (new_AGEMA_signal_3870), .Z1_t (new_AGEMA_signal_3871), .Z1_f (new_AGEMA_signal_3872) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U9 ( .A0_t (Midori_rounds_roundReg_out[14]), .A0_f (new_AGEMA_signal_2874), .A1_t (new_AGEMA_signal_2875), .A1_f (new_AGEMA_signal_2876), .B0_t (Midori_rounds_roundReg_out[15]), .B0_f (new_AGEMA_signal_2877), .B1_t (new_AGEMA_signal_2878), .B1_f (new_AGEMA_signal_2879), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n14), .Z0_f (new_AGEMA_signal_2889), .Z1_t (new_AGEMA_signal_2890), .Z1_f (new_AGEMA_signal_2891) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U8 ( .A0_t (Midori_rounds_roundReg_out[15]), .A0_f (new_AGEMA_signal_2877), .A1_t (new_AGEMA_signal_2878), .A1_f (new_AGEMA_signal_2879), .B0_t (Midori_rounds_roundReg_out[12]), .B0_f (new_AGEMA_signal_2883), .B1_t (new_AGEMA_signal_2884), .B1_f (new_AGEMA_signal_2885), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n9), .Z0_f (new_AGEMA_signal_2892), .Z1_t (new_AGEMA_signal_2893), .Z1_f (new_AGEMA_signal_2894) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n3), .A0_f (new_AGEMA_signal_2898), .A1_t (new_AGEMA_signal_2899), .A1_f (new_AGEMA_signal_2900), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n2), .B0_f (new_AGEMA_signal_3873), .B1_t (new_AGEMA_signal_3874), .B1_f (new_AGEMA_signal_3875), .Z0_t (Midori_rounds_SR_Result[21]), .Z0_f (new_AGEMA_signal_4325), .Z1_t (new_AGEMA_signal_4326), .Z1_f (new_AGEMA_signal_4327) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n1), .A0_f (new_AGEMA_signal_2895), .A1_t (new_AGEMA_signal_2896), .A1_f (new_AGEMA_signal_2897), .B0_t (Midori_rounds_roundReg_out[15]), .B0_f (new_AGEMA_signal_2877), .B1_t (new_AGEMA_signal_2878), .B1_f (new_AGEMA_signal_2879), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n2), .Z0_f (new_AGEMA_signal_3873), .Z1_t (new_AGEMA_signal_3874), .Z1_f (new_AGEMA_signal_3875) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U4 ( .A0_t (Midori_rounds_roundReg_out[14]), .A0_f (new_AGEMA_signal_2874), .A1_t (new_AGEMA_signal_2875), .A1_f (new_AGEMA_signal_2876), .B0_t (Midori_rounds_roundReg_out[12]), .B0_f (new_AGEMA_signal_2883), .B1_t (new_AGEMA_signal_2884), .B1_f (new_AGEMA_signal_2885), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n1), .Z0_f (new_AGEMA_signal_2895), .Z1_t (new_AGEMA_signal_2896), .Z1_f (new_AGEMA_signal_2897) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U1 ( .A0_t (Midori_rounds_roundReg_out[14]), .A0_f (new_AGEMA_signal_2874), .A1_t (new_AGEMA_signal_2875), .A1_f (new_AGEMA_signal_2876), .B0_t (Midori_rounds_roundReg_out[12]), .B0_f (new_AGEMA_signal_2883), .B1_t (new_AGEMA_signal_2884), .B1_f (new_AGEMA_signal_2885), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n3), .Z0_f (new_AGEMA_signal_2898), .Z1_t (new_AGEMA_signal_2899), .Z1_f (new_AGEMA_signal_2900) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n15), .A0_f (new_AGEMA_signal_4328), .A1_t (new_AGEMA_signal_4329), .A1_f (new_AGEMA_signal_4330), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n14), .B0_f (new_AGEMA_signal_2916), .B1_t (new_AGEMA_signal_2917), .B1_f (new_AGEMA_signal_2918), .Z0_t (Midori_rounds_SR_Result[36]), .Z0_f (new_AGEMA_signal_4706), .Z1_t (new_AGEMA_signal_4707), .Z1_f (new_AGEMA_signal_4708) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U18 ( .A0_t (Midori_rounds_roundReg_out[17]), .A0_f (new_AGEMA_signal_3882), .A1_t (new_AGEMA_signal_3883), .A1_f (new_AGEMA_signal_3884), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n13), .B0_f (new_AGEMA_signal_3876), .B1_t (new_AGEMA_signal_3877), .B1_f (new_AGEMA_signal_3878), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n15), .Z0_f (new_AGEMA_signal_4328), .Z1_t (new_AGEMA_signal_4329), .Z1_f (new_AGEMA_signal_4330) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U17 ( .A0_t (Midori_rounds_roundReg_out[16]), .A0_f (new_AGEMA_signal_2910), .A1_t (new_AGEMA_signal_2911), .A1_f (new_AGEMA_signal_2912), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n11), .B0_f (new_AGEMA_signal_2907), .B1_t (new_AGEMA_signal_2908), .B1_f (new_AGEMA_signal_2909), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n13), .Z0_f (new_AGEMA_signal_3876), .Z1_t (new_AGEMA_signal_3877), .Z1_f (new_AGEMA_signal_3878) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U16 ( .A0_t (Midori_rounds_roundReg_out[18]), .A0_f (new_AGEMA_signal_2901), .A1_t (new_AGEMA_signal_2902), .A1_f (new_AGEMA_signal_2903), .B0_t (Midori_rounds_roundReg_out[19]), .B0_f (new_AGEMA_signal_2904), .B1_t (new_AGEMA_signal_2905), .B1_f (new_AGEMA_signal_2906), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n11), .Z0_f (new_AGEMA_signal_2907), .Z1_t (new_AGEMA_signal_2908), .Z1_f (new_AGEMA_signal_2909) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n10), .A0_f (new_AGEMA_signal_4331), .A1_t (new_AGEMA_signal_4332), .A1_f (new_AGEMA_signal_4333), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n9), .B0_f (new_AGEMA_signal_2919), .B1_t (new_AGEMA_signal_2920), .B1_f (new_AGEMA_signal_2921), .Z0_t (Midori_rounds_SR_Result[38]), .Z0_f (new_AGEMA_signal_4709), .Z1_t (new_AGEMA_signal_4710), .Z1_f (new_AGEMA_signal_4711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n8), .A0_f (new_AGEMA_signal_3879), .A1_t (new_AGEMA_signal_3880), .A1_f (new_AGEMA_signal_3881), .B0_t (Midori_rounds_roundReg_out[17]), .B0_f (new_AGEMA_signal_3882), .B1_t (new_AGEMA_signal_3883), .B1_f (new_AGEMA_signal_3884), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n10), .Z0_f (new_AGEMA_signal_4331), .Z1_t (new_AGEMA_signal_4332), .Z1_f (new_AGEMA_signal_4333) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n7), .A0_f (new_AGEMA_signal_2913), .A1_t (new_AGEMA_signal_2914), .A1_f (new_AGEMA_signal_2915), .B0_t (Midori_rounds_roundReg_out[18]), .B0_f (new_AGEMA_signal_2901), .B1_t (new_AGEMA_signal_2902), .B1_f (new_AGEMA_signal_2903), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n8), .Z0_f (new_AGEMA_signal_3879), .Z1_t (new_AGEMA_signal_3880), .Z1_f (new_AGEMA_signal_3881) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U12 ( .A0_t (Midori_rounds_roundReg_out[16]), .A0_f (new_AGEMA_signal_2910), .A1_t (new_AGEMA_signal_2911), .A1_f (new_AGEMA_signal_2912), .B0_t (Midori_rounds_roundReg_out[19]), .B0_f (new_AGEMA_signal_2904), .B1_t (new_AGEMA_signal_2905), .B1_f (new_AGEMA_signal_2906), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n7), .Z0_f (new_AGEMA_signal_2913), .Z1_t (new_AGEMA_signal_2914), .Z1_f (new_AGEMA_signal_2915) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n9), .A0_f (new_AGEMA_signal_2919), .A1_t (new_AGEMA_signal_2920), .A1_f (new_AGEMA_signal_2921), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n5), .B0_f (new_AGEMA_signal_3885), .B1_t (new_AGEMA_signal_3886), .B1_f (new_AGEMA_signal_3887), .Z0_t (Midori_rounds_SR_Result[39]), .Z0_f (new_AGEMA_signal_4334), .Z1_t (new_AGEMA_signal_4335), .Z1_f (new_AGEMA_signal_4336) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U10 ( .A0_t (Midori_rounds_roundReg_out[17]), .A0_f (new_AGEMA_signal_3882), .A1_t (new_AGEMA_signal_3883), .A1_f (new_AGEMA_signal_3884), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n14), .B0_f (new_AGEMA_signal_2916), .B1_t (new_AGEMA_signal_2917), .B1_f (new_AGEMA_signal_2918), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n5), .Z0_f (new_AGEMA_signal_3885), .Z1_t (new_AGEMA_signal_3886), .Z1_f (new_AGEMA_signal_3887) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U9 ( .A0_t (Midori_rounds_roundReg_out[18]), .A0_f (new_AGEMA_signal_2901), .A1_t (new_AGEMA_signal_2902), .A1_f (new_AGEMA_signal_2903), .B0_t (Midori_rounds_roundReg_out[19]), .B0_f (new_AGEMA_signal_2904), .B1_t (new_AGEMA_signal_2905), .B1_f (new_AGEMA_signal_2906), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n14), .Z0_f (new_AGEMA_signal_2916), .Z1_t (new_AGEMA_signal_2917), .Z1_f (new_AGEMA_signal_2918) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U8 ( .A0_t (Midori_rounds_roundReg_out[19]), .A0_f (new_AGEMA_signal_2904), .A1_t (new_AGEMA_signal_2905), .A1_f (new_AGEMA_signal_2906), .B0_t (Midori_rounds_roundReg_out[16]), .B0_f (new_AGEMA_signal_2910), .B1_t (new_AGEMA_signal_2911), .B1_f (new_AGEMA_signal_2912), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n9), .Z0_f (new_AGEMA_signal_2919), .Z1_t (new_AGEMA_signal_2920), .Z1_f (new_AGEMA_signal_2921) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n3), .A0_f (new_AGEMA_signal_2925), .A1_t (new_AGEMA_signal_2926), .A1_f (new_AGEMA_signal_2927), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n2), .B0_f (new_AGEMA_signal_3888), .B1_t (new_AGEMA_signal_3889), .B1_f (new_AGEMA_signal_3890), .Z0_t (Midori_rounds_SR_Result[37]), .Z0_f (new_AGEMA_signal_4337), .Z1_t (new_AGEMA_signal_4338), .Z1_f (new_AGEMA_signal_4339) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n1), .A0_f (new_AGEMA_signal_2922), .A1_t (new_AGEMA_signal_2923), .A1_f (new_AGEMA_signal_2924), .B0_t (Midori_rounds_roundReg_out[19]), .B0_f (new_AGEMA_signal_2904), .B1_t (new_AGEMA_signal_2905), .B1_f (new_AGEMA_signal_2906), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n2), .Z0_f (new_AGEMA_signal_3888), .Z1_t (new_AGEMA_signal_3889), .Z1_f (new_AGEMA_signal_3890) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U4 ( .A0_t (Midori_rounds_roundReg_out[18]), .A0_f (new_AGEMA_signal_2901), .A1_t (new_AGEMA_signal_2902), .A1_f (new_AGEMA_signal_2903), .B0_t (Midori_rounds_roundReg_out[16]), .B0_f (new_AGEMA_signal_2910), .B1_t (new_AGEMA_signal_2911), .B1_f (new_AGEMA_signal_2912), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n1), .Z0_f (new_AGEMA_signal_2922), .Z1_t (new_AGEMA_signal_2923), .Z1_f (new_AGEMA_signal_2924) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U1 ( .A0_t (Midori_rounds_roundReg_out[18]), .A0_f (new_AGEMA_signal_2901), .A1_t (new_AGEMA_signal_2902), .A1_f (new_AGEMA_signal_2903), .B0_t (Midori_rounds_roundReg_out[16]), .B0_f (new_AGEMA_signal_2910), .B1_t (new_AGEMA_signal_2911), .B1_f (new_AGEMA_signal_2912), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n3), .Z0_f (new_AGEMA_signal_2925), .Z1_t (new_AGEMA_signal_2926), .Z1_f (new_AGEMA_signal_2927) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n15), .A0_f (new_AGEMA_signal_4340), .A1_t (new_AGEMA_signal_4341), .A1_f (new_AGEMA_signal_4342), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n14), .B0_f (new_AGEMA_signal_2943), .B1_t (new_AGEMA_signal_2944), .B1_f (new_AGEMA_signal_2945), .Z0_t (Midori_rounds_SR_Result[56]), .Z0_f (new_AGEMA_signal_4712), .Z1_t (new_AGEMA_signal_4713), .Z1_f (new_AGEMA_signal_4714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U18 ( .A0_t (Midori_rounds_roundReg_out[21]), .A0_f (new_AGEMA_signal_3897), .A1_t (new_AGEMA_signal_3898), .A1_f (new_AGEMA_signal_3899), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n13), .B0_f (new_AGEMA_signal_3891), .B1_t (new_AGEMA_signal_3892), .B1_f (new_AGEMA_signal_3893), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n15), .Z0_f (new_AGEMA_signal_4340), .Z1_t (new_AGEMA_signal_4341), .Z1_f (new_AGEMA_signal_4342) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U17 ( .A0_t (Midori_rounds_roundReg_out[20]), .A0_f (new_AGEMA_signal_2937), .A1_t (new_AGEMA_signal_2938), .A1_f (new_AGEMA_signal_2939), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n11), .B0_f (new_AGEMA_signal_2934), .B1_t (new_AGEMA_signal_2935), .B1_f (new_AGEMA_signal_2936), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n13), .Z0_f (new_AGEMA_signal_3891), .Z1_t (new_AGEMA_signal_3892), .Z1_f (new_AGEMA_signal_3893) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U16 ( .A0_t (Midori_rounds_roundReg_out[22]), .A0_f (new_AGEMA_signal_2928), .A1_t (new_AGEMA_signal_2929), .A1_f (new_AGEMA_signal_2930), .B0_t (Midori_rounds_roundReg_out[23]), .B0_f (new_AGEMA_signal_2931), .B1_t (new_AGEMA_signal_2932), .B1_f (new_AGEMA_signal_2933), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n11), .Z0_f (new_AGEMA_signal_2934), .Z1_t (new_AGEMA_signal_2935), .Z1_f (new_AGEMA_signal_2936) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n10), .A0_f (new_AGEMA_signal_4343), .A1_t (new_AGEMA_signal_4344), .A1_f (new_AGEMA_signal_4345), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n9), .B0_f (new_AGEMA_signal_2946), .B1_t (new_AGEMA_signal_2947), .B1_f (new_AGEMA_signal_2948), .Z0_t (Midori_rounds_SR_Result[58]), .Z0_f (new_AGEMA_signal_4715), .Z1_t (new_AGEMA_signal_4716), .Z1_f (new_AGEMA_signal_4717) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n8), .A0_f (new_AGEMA_signal_3894), .A1_t (new_AGEMA_signal_3895), .A1_f (new_AGEMA_signal_3896), .B0_t (Midori_rounds_roundReg_out[21]), .B0_f (new_AGEMA_signal_3897), .B1_t (new_AGEMA_signal_3898), .B1_f (new_AGEMA_signal_3899), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n10), .Z0_f (new_AGEMA_signal_4343), .Z1_t (new_AGEMA_signal_4344), .Z1_f (new_AGEMA_signal_4345) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n7), .A0_f (new_AGEMA_signal_2940), .A1_t (new_AGEMA_signal_2941), .A1_f (new_AGEMA_signal_2942), .B0_t (Midori_rounds_roundReg_out[22]), .B0_f (new_AGEMA_signal_2928), .B1_t (new_AGEMA_signal_2929), .B1_f (new_AGEMA_signal_2930), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n8), .Z0_f (new_AGEMA_signal_3894), .Z1_t (new_AGEMA_signal_3895), .Z1_f (new_AGEMA_signal_3896) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U12 ( .A0_t (Midori_rounds_roundReg_out[20]), .A0_f (new_AGEMA_signal_2937), .A1_t (new_AGEMA_signal_2938), .A1_f (new_AGEMA_signal_2939), .B0_t (Midori_rounds_roundReg_out[23]), .B0_f (new_AGEMA_signal_2931), .B1_t (new_AGEMA_signal_2932), .B1_f (new_AGEMA_signal_2933), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n7), .Z0_f (new_AGEMA_signal_2940), .Z1_t (new_AGEMA_signal_2941), .Z1_f (new_AGEMA_signal_2942) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n9), .A0_f (new_AGEMA_signal_2946), .A1_t (new_AGEMA_signal_2947), .A1_f (new_AGEMA_signal_2948), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n5), .B0_f (new_AGEMA_signal_3900), .B1_t (new_AGEMA_signal_3901), .B1_f (new_AGEMA_signal_3902), .Z0_t (Midori_rounds_SR_Result[59]), .Z0_f (new_AGEMA_signal_4346), .Z1_t (new_AGEMA_signal_4347), .Z1_f (new_AGEMA_signal_4348) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U10 ( .A0_t (Midori_rounds_roundReg_out[21]), .A0_f (new_AGEMA_signal_3897), .A1_t (new_AGEMA_signal_3898), .A1_f (new_AGEMA_signal_3899), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n14), .B0_f (new_AGEMA_signal_2943), .B1_t (new_AGEMA_signal_2944), .B1_f (new_AGEMA_signal_2945), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n5), .Z0_f (new_AGEMA_signal_3900), .Z1_t (new_AGEMA_signal_3901), .Z1_f (new_AGEMA_signal_3902) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U9 ( .A0_t (Midori_rounds_roundReg_out[22]), .A0_f (new_AGEMA_signal_2928), .A1_t (new_AGEMA_signal_2929), .A1_f (new_AGEMA_signal_2930), .B0_t (Midori_rounds_roundReg_out[23]), .B0_f (new_AGEMA_signal_2931), .B1_t (new_AGEMA_signal_2932), .B1_f (new_AGEMA_signal_2933), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n14), .Z0_f (new_AGEMA_signal_2943), .Z1_t (new_AGEMA_signal_2944), .Z1_f (new_AGEMA_signal_2945) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U8 ( .A0_t (Midori_rounds_roundReg_out[23]), .A0_f (new_AGEMA_signal_2931), .A1_t (new_AGEMA_signal_2932), .A1_f (new_AGEMA_signal_2933), .B0_t (Midori_rounds_roundReg_out[20]), .B0_f (new_AGEMA_signal_2937), .B1_t (new_AGEMA_signal_2938), .B1_f (new_AGEMA_signal_2939), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n9), .Z0_f (new_AGEMA_signal_2946), .Z1_t (new_AGEMA_signal_2947), .Z1_f (new_AGEMA_signal_2948) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n3), .A0_f (new_AGEMA_signal_2952), .A1_t (new_AGEMA_signal_2953), .A1_f (new_AGEMA_signal_2954), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n2), .B0_f (new_AGEMA_signal_3903), .B1_t (new_AGEMA_signal_3904), .B1_f (new_AGEMA_signal_3905), .Z0_t (Midori_rounds_SR_Result[57]), .Z0_f (new_AGEMA_signal_4349), .Z1_t (new_AGEMA_signal_4350), .Z1_f (new_AGEMA_signal_4351) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n1), .A0_f (new_AGEMA_signal_2949), .A1_t (new_AGEMA_signal_2950), .A1_f (new_AGEMA_signal_2951), .B0_t (Midori_rounds_roundReg_out[23]), .B0_f (new_AGEMA_signal_2931), .B1_t (new_AGEMA_signal_2932), .B1_f (new_AGEMA_signal_2933), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n2), .Z0_f (new_AGEMA_signal_3903), .Z1_t (new_AGEMA_signal_3904), .Z1_f (new_AGEMA_signal_3905) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U4 ( .A0_t (Midori_rounds_roundReg_out[22]), .A0_f (new_AGEMA_signal_2928), .A1_t (new_AGEMA_signal_2929), .A1_f (new_AGEMA_signal_2930), .B0_t (Midori_rounds_roundReg_out[20]), .B0_f (new_AGEMA_signal_2937), .B1_t (new_AGEMA_signal_2938), .B1_f (new_AGEMA_signal_2939), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n1), .Z0_f (new_AGEMA_signal_2949), .Z1_t (new_AGEMA_signal_2950), .Z1_f (new_AGEMA_signal_2951) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U1 ( .A0_t (Midori_rounds_roundReg_out[22]), .A0_f (new_AGEMA_signal_2928), .A1_t (new_AGEMA_signal_2929), .A1_f (new_AGEMA_signal_2930), .B0_t (Midori_rounds_roundReg_out[20]), .B0_f (new_AGEMA_signal_2937), .B1_t (new_AGEMA_signal_2938), .B1_f (new_AGEMA_signal_2939), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n3), .Z0_f (new_AGEMA_signal_2952), .Z1_t (new_AGEMA_signal_2953), .Z1_f (new_AGEMA_signal_2954) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n15), .A0_f (new_AGEMA_signal_4352), .A1_t (new_AGEMA_signal_4353), .A1_f (new_AGEMA_signal_4354), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n14), .B0_f (new_AGEMA_signal_2970), .B1_t (new_AGEMA_signal_2971), .B1_f (new_AGEMA_signal_2972), .Z0_t (Midori_rounds_SR_Result[28]), .Z0_f (new_AGEMA_signal_4718), .Z1_t (new_AGEMA_signal_4719), .Z1_f (new_AGEMA_signal_4720) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U18 ( .A0_t (Midori_rounds_roundReg_out[25]), .A0_f (new_AGEMA_signal_3912), .A1_t (new_AGEMA_signal_3913), .A1_f (new_AGEMA_signal_3914), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n13), .B0_f (new_AGEMA_signal_3906), .B1_t (new_AGEMA_signal_3907), .B1_f (new_AGEMA_signal_3908), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n15), .Z0_f (new_AGEMA_signal_4352), .Z1_t (new_AGEMA_signal_4353), .Z1_f (new_AGEMA_signal_4354) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U17 ( .A0_t (Midori_rounds_roundReg_out[24]), .A0_f (new_AGEMA_signal_2964), .A1_t (new_AGEMA_signal_2965), .A1_f (new_AGEMA_signal_2966), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n11), .B0_f (new_AGEMA_signal_2961), .B1_t (new_AGEMA_signal_2962), .B1_f (new_AGEMA_signal_2963), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n13), .Z0_f (new_AGEMA_signal_3906), .Z1_t (new_AGEMA_signal_3907), .Z1_f (new_AGEMA_signal_3908) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U16 ( .A0_t (Midori_rounds_roundReg_out[26]), .A0_f (new_AGEMA_signal_2955), .A1_t (new_AGEMA_signal_2956), .A1_f (new_AGEMA_signal_2957), .B0_t (Midori_rounds_roundReg_out[27]), .B0_f (new_AGEMA_signal_2958), .B1_t (new_AGEMA_signal_2959), .B1_f (new_AGEMA_signal_2960), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n11), .Z0_f (new_AGEMA_signal_2961), .Z1_t (new_AGEMA_signal_2962), .Z1_f (new_AGEMA_signal_2963) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n10), .A0_f (new_AGEMA_signal_4355), .A1_t (new_AGEMA_signal_4356), .A1_f (new_AGEMA_signal_4357), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n9), .B0_f (new_AGEMA_signal_2973), .B1_t (new_AGEMA_signal_2974), .B1_f (new_AGEMA_signal_2975), .Z0_t (Midori_rounds_SR_Result[30]), .Z0_f (new_AGEMA_signal_4721), .Z1_t (new_AGEMA_signal_4722), .Z1_f (new_AGEMA_signal_4723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n8), .A0_f (new_AGEMA_signal_3909), .A1_t (new_AGEMA_signal_3910), .A1_f (new_AGEMA_signal_3911), .B0_t (Midori_rounds_roundReg_out[25]), .B0_f (new_AGEMA_signal_3912), .B1_t (new_AGEMA_signal_3913), .B1_f (new_AGEMA_signal_3914), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n10), .Z0_f (new_AGEMA_signal_4355), .Z1_t (new_AGEMA_signal_4356), .Z1_f (new_AGEMA_signal_4357) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n7), .A0_f (new_AGEMA_signal_2967), .A1_t (new_AGEMA_signal_2968), .A1_f (new_AGEMA_signal_2969), .B0_t (Midori_rounds_roundReg_out[26]), .B0_f (new_AGEMA_signal_2955), .B1_t (new_AGEMA_signal_2956), .B1_f (new_AGEMA_signal_2957), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n8), .Z0_f (new_AGEMA_signal_3909), .Z1_t (new_AGEMA_signal_3910), .Z1_f (new_AGEMA_signal_3911) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U12 ( .A0_t (Midori_rounds_roundReg_out[24]), .A0_f (new_AGEMA_signal_2964), .A1_t (new_AGEMA_signal_2965), .A1_f (new_AGEMA_signal_2966), .B0_t (Midori_rounds_roundReg_out[27]), .B0_f (new_AGEMA_signal_2958), .B1_t (new_AGEMA_signal_2959), .B1_f (new_AGEMA_signal_2960), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n7), .Z0_f (new_AGEMA_signal_2967), .Z1_t (new_AGEMA_signal_2968), .Z1_f (new_AGEMA_signal_2969) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n9), .A0_f (new_AGEMA_signal_2973), .A1_t (new_AGEMA_signal_2974), .A1_f (new_AGEMA_signal_2975), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n5), .B0_f (new_AGEMA_signal_3915), .B1_t (new_AGEMA_signal_3916), .B1_f (new_AGEMA_signal_3917), .Z0_t (Midori_rounds_SR_Result[31]), .Z0_f (new_AGEMA_signal_4358), .Z1_t (new_AGEMA_signal_4359), .Z1_f (new_AGEMA_signal_4360) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U10 ( .A0_t (Midori_rounds_roundReg_out[25]), .A0_f (new_AGEMA_signal_3912), .A1_t (new_AGEMA_signal_3913), .A1_f (new_AGEMA_signal_3914), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n14), .B0_f (new_AGEMA_signal_2970), .B1_t (new_AGEMA_signal_2971), .B1_f (new_AGEMA_signal_2972), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n5), .Z0_f (new_AGEMA_signal_3915), .Z1_t (new_AGEMA_signal_3916), .Z1_f (new_AGEMA_signal_3917) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U9 ( .A0_t (Midori_rounds_roundReg_out[26]), .A0_f (new_AGEMA_signal_2955), .A1_t (new_AGEMA_signal_2956), .A1_f (new_AGEMA_signal_2957), .B0_t (Midori_rounds_roundReg_out[27]), .B0_f (new_AGEMA_signal_2958), .B1_t (new_AGEMA_signal_2959), .B1_f (new_AGEMA_signal_2960), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n14), .Z0_f (new_AGEMA_signal_2970), .Z1_t (new_AGEMA_signal_2971), .Z1_f (new_AGEMA_signal_2972) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U8 ( .A0_t (Midori_rounds_roundReg_out[27]), .A0_f (new_AGEMA_signal_2958), .A1_t (new_AGEMA_signal_2959), .A1_f (new_AGEMA_signal_2960), .B0_t (Midori_rounds_roundReg_out[24]), .B0_f (new_AGEMA_signal_2964), .B1_t (new_AGEMA_signal_2965), .B1_f (new_AGEMA_signal_2966), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n9), .Z0_f (new_AGEMA_signal_2973), .Z1_t (new_AGEMA_signal_2974), .Z1_f (new_AGEMA_signal_2975) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n3), .A0_f (new_AGEMA_signal_2979), .A1_t (new_AGEMA_signal_2980), .A1_f (new_AGEMA_signal_2981), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n2), .B0_f (new_AGEMA_signal_3918), .B1_t (new_AGEMA_signal_3919), .B1_f (new_AGEMA_signal_3920), .Z0_t (Midori_rounds_SR_Result[29]), .Z0_f (new_AGEMA_signal_4361), .Z1_t (new_AGEMA_signal_4362), .Z1_f (new_AGEMA_signal_4363) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n1), .A0_f (new_AGEMA_signal_2976), .A1_t (new_AGEMA_signal_2977), .A1_f (new_AGEMA_signal_2978), .B0_t (Midori_rounds_roundReg_out[27]), .B0_f (new_AGEMA_signal_2958), .B1_t (new_AGEMA_signal_2959), .B1_f (new_AGEMA_signal_2960), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n2), .Z0_f (new_AGEMA_signal_3918), .Z1_t (new_AGEMA_signal_3919), .Z1_f (new_AGEMA_signal_3920) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U4 ( .A0_t (Midori_rounds_roundReg_out[26]), .A0_f (new_AGEMA_signal_2955), .A1_t (new_AGEMA_signal_2956), .A1_f (new_AGEMA_signal_2957), .B0_t (Midori_rounds_roundReg_out[24]), .B0_f (new_AGEMA_signal_2964), .B1_t (new_AGEMA_signal_2965), .B1_f (new_AGEMA_signal_2966), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n1), .Z0_f (new_AGEMA_signal_2976), .Z1_t (new_AGEMA_signal_2977), .Z1_f (new_AGEMA_signal_2978) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U1 ( .A0_t (Midori_rounds_roundReg_out[26]), .A0_f (new_AGEMA_signal_2955), .A1_t (new_AGEMA_signal_2956), .A1_f (new_AGEMA_signal_2957), .B0_t (Midori_rounds_roundReg_out[24]), .B0_f (new_AGEMA_signal_2964), .B1_t (new_AGEMA_signal_2965), .B1_f (new_AGEMA_signal_2966), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n3), .Z0_f (new_AGEMA_signal_2979), .Z1_t (new_AGEMA_signal_2980), .Z1_f (new_AGEMA_signal_2981) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n15), .A0_f (new_AGEMA_signal_3000), .A1_t (new_AGEMA_signal_3001), .A1_f (new_AGEMA_signal_3002), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n14), .B0_f (new_AGEMA_signal_3924), .B1_t (new_AGEMA_signal_3925), .B1_f (new_AGEMA_signal_3926), .Z0_t (Midori_rounds_SR_Result[3]), .Z0_f (new_AGEMA_signal_4364), .Z1_t (new_AGEMA_signal_4365), .Z1_f (new_AGEMA_signal_4366) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n13), .A0_f (new_AGEMA_signal_3006), .A1_t (new_AGEMA_signal_3007), .A1_f (new_AGEMA_signal_3008), .B0_t (Midori_rounds_roundReg_out[29]), .B0_f (new_AGEMA_signal_3921), .B1_t (new_AGEMA_signal_3922), .B1_f (new_AGEMA_signal_3923), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n14), .Z0_f (new_AGEMA_signal_3924), .Z1_t (new_AGEMA_signal_3925), .Z1_f (new_AGEMA_signal_3926) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n12), .A0_f (new_AGEMA_signal_2991), .A1_t (new_AGEMA_signal_2992), .A1_f (new_AGEMA_signal_2993), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n11), .B0_f (new_AGEMA_signal_3927), .B1_t (new_AGEMA_signal_3928), .B1_f (new_AGEMA_signal_3929), .Z0_t (Midori_rounds_SR_Result[1]), .Z0_f (new_AGEMA_signal_4367), .Z1_t (new_AGEMA_signal_4368), .Z1_f (new_AGEMA_signal_4369) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U16 ( .A0_t (Midori_rounds_roundReg_out[28]), .A0_f (new_AGEMA_signal_2994), .A1_t (new_AGEMA_signal_2995), .A1_f (new_AGEMA_signal_2996), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n10), .B0_f (new_AGEMA_signal_2988), .B1_t (new_AGEMA_signal_2989), .B1_f (new_AGEMA_signal_2990), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n11), .Z0_f (new_AGEMA_signal_3927), .Z1_t (new_AGEMA_signal_3928), .Z1_f (new_AGEMA_signal_3929) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U15 ( .A0_t (Midori_rounds_roundReg_out[31]), .A0_f (new_AGEMA_signal_2982), .A1_t (new_AGEMA_signal_2983), .A1_f (new_AGEMA_signal_2984), .B0_t (Midori_rounds_roundReg_out[30]), .B0_f (new_AGEMA_signal_2985), .B1_t (new_AGEMA_signal_2986), .B1_f (new_AGEMA_signal_2987), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n10), .Z0_f (new_AGEMA_signal_2988), .Z1_t (new_AGEMA_signal_2989), .Z1_f (new_AGEMA_signal_2990) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U14 ( .A0_t (Midori_rounds_roundReg_out[30]), .A0_f (new_AGEMA_signal_2985), .A1_t (new_AGEMA_signal_2986), .A1_f (new_AGEMA_signal_2987), .B0_t (Midori_rounds_roundReg_out[31]), .B0_f (new_AGEMA_signal_2982), .B1_t (new_AGEMA_signal_2983), .B1_f (new_AGEMA_signal_2984), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n12), .Z0_f (new_AGEMA_signal_2991), .Z1_t (new_AGEMA_signal_2992), .Z1_f (new_AGEMA_signal_2993) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n15), .A0_f (new_AGEMA_signal_3000), .A1_t (new_AGEMA_signal_3001), .A1_f (new_AGEMA_signal_3002), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n7), .B0_f (new_AGEMA_signal_4370), .B1_t (new_AGEMA_signal_4371), .B1_f (new_AGEMA_signal_4372), .Z0_t (Midori_rounds_SR_Result[2]), .Z0_f (new_AGEMA_signal_4724), .Z1_t (new_AGEMA_signal_4725), .Z1_f (new_AGEMA_signal_4726) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n6), .A0_f (new_AGEMA_signal_3930), .A1_t (new_AGEMA_signal_3931), .A1_f (new_AGEMA_signal_3932), .B0_t (Midori_rounds_roundReg_out[29]), .B0_f (new_AGEMA_signal_3921), .B1_t (new_AGEMA_signal_3922), .B1_f (new_AGEMA_signal_3923), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n7), .Z0_f (new_AGEMA_signal_4370), .Z1_t (new_AGEMA_signal_4371), .Z1_f (new_AGEMA_signal_4372) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n5), .A0_f (new_AGEMA_signal_2997), .A1_t (new_AGEMA_signal_2998), .A1_f (new_AGEMA_signal_2999), .B0_t (Midori_rounds_roundReg_out[30]), .B0_f (new_AGEMA_signal_2985), .B1_t (new_AGEMA_signal_2986), .B1_f (new_AGEMA_signal_2987), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n6), .Z0_f (new_AGEMA_signal_3930), .Z1_t (new_AGEMA_signal_3931), .Z1_f (new_AGEMA_signal_3932) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U10 ( .A0_t (Midori_rounds_roundReg_out[28]), .A0_f (new_AGEMA_signal_2994), .A1_t (new_AGEMA_signal_2995), .A1_f (new_AGEMA_signal_2996), .B0_t (Midori_rounds_roundReg_out[31]), .B0_f (new_AGEMA_signal_2982), .B1_t (new_AGEMA_signal_2983), .B1_f (new_AGEMA_signal_2984), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n5), .Z0_f (new_AGEMA_signal_2997), .Z1_t (new_AGEMA_signal_2998), .Z1_f (new_AGEMA_signal_2999) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U9 ( .A0_t (Midori_rounds_roundReg_out[31]), .A0_f (new_AGEMA_signal_2982), .A1_t (new_AGEMA_signal_2983), .A1_f (new_AGEMA_signal_2984), .B0_t (Midori_rounds_roundReg_out[28]), .B0_f (new_AGEMA_signal_2994), .B1_t (new_AGEMA_signal_2995), .B1_f (new_AGEMA_signal_2996), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n15), .Z0_f (new_AGEMA_signal_3000), .Z1_t (new_AGEMA_signal_3001), .Z1_f (new_AGEMA_signal_3002) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n13), .A0_f (new_AGEMA_signal_3006), .A1_t (new_AGEMA_signal_3007), .A1_f (new_AGEMA_signal_3008), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n3), .B0_f (new_AGEMA_signal_4373), .B1_t (new_AGEMA_signal_4374), .B1_f (new_AGEMA_signal_4375), .Z0_t (Midori_rounds_SR_Result[0]), .Z0_f (new_AGEMA_signal_4727), .Z1_t (new_AGEMA_signal_4728), .Z1_f (new_AGEMA_signal_4729) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U7 ( .A0_t (Midori_rounds_roundReg_out[29]), .A0_f (new_AGEMA_signal_3921), .A1_t (new_AGEMA_signal_3922), .A1_f (new_AGEMA_signal_3923), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n2), .B0_f (new_AGEMA_signal_3933), .B1_t (new_AGEMA_signal_3934), .B1_f (new_AGEMA_signal_3935), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n3), .Z0_f (new_AGEMA_signal_4373), .Z1_t (new_AGEMA_signal_4374), .Z1_f (new_AGEMA_signal_4375) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U6 ( .A0_t (Midori_rounds_roundReg_out[28]), .A0_f (new_AGEMA_signal_2994), .A1_t (new_AGEMA_signal_2995), .A1_f (new_AGEMA_signal_2996), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n1), .B0_f (new_AGEMA_signal_3003), .B1_t (new_AGEMA_signal_3004), .B1_f (new_AGEMA_signal_3005), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n2), .Z0_f (new_AGEMA_signal_3933), .Z1_t (new_AGEMA_signal_3934), .Z1_f (new_AGEMA_signal_3935) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U5 ( .A0_t (Midori_rounds_roundReg_out[30]), .A0_f (new_AGEMA_signal_2985), .A1_t (new_AGEMA_signal_2986), .A1_f (new_AGEMA_signal_2987), .B0_t (Midori_rounds_roundReg_out[31]), .B0_f (new_AGEMA_signal_2982), .B1_t (new_AGEMA_signal_2983), .B1_f (new_AGEMA_signal_2984), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n1), .Z0_f (new_AGEMA_signal_3003), .Z1_t (new_AGEMA_signal_3004), .Z1_f (new_AGEMA_signal_3005) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U3 ( .A0_t (Midori_rounds_roundReg_out[30]), .A0_f (new_AGEMA_signal_2985), .A1_t (new_AGEMA_signal_2986), .A1_f (new_AGEMA_signal_2987), .B0_t (Midori_rounds_roundReg_out[31]), .B0_f (new_AGEMA_signal_2982), .B1_t (new_AGEMA_signal_2983), .B1_f (new_AGEMA_signal_2984), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n13), .Z0_f (new_AGEMA_signal_3006), .Z1_t (new_AGEMA_signal_3007), .Z1_f (new_AGEMA_signal_3008) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n15), .A0_f (new_AGEMA_signal_3027), .A1_t (new_AGEMA_signal_3028), .A1_f (new_AGEMA_signal_3029), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n14), .B0_f (new_AGEMA_signal_3939), .B1_t (new_AGEMA_signal_3940), .B1_f (new_AGEMA_signal_3941), .Z0_t (Midori_rounds_SR_Result[15]), .Z0_f (new_AGEMA_signal_4376), .Z1_t (new_AGEMA_signal_4377), .Z1_f (new_AGEMA_signal_4378) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n13), .A0_f (new_AGEMA_signal_3033), .A1_t (new_AGEMA_signal_3034), .A1_f (new_AGEMA_signal_3035), .B0_t (Midori_rounds_roundReg_out[33]), .B0_f (new_AGEMA_signal_3936), .B1_t (new_AGEMA_signal_3937), .B1_f (new_AGEMA_signal_3938), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n14), .Z0_f (new_AGEMA_signal_3939), .Z1_t (new_AGEMA_signal_3940), .Z1_f (new_AGEMA_signal_3941) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n12), .A0_f (new_AGEMA_signal_3018), .A1_t (new_AGEMA_signal_3019), .A1_f (new_AGEMA_signal_3020), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n11), .B0_f (new_AGEMA_signal_3942), .B1_t (new_AGEMA_signal_3943), .B1_f (new_AGEMA_signal_3944), .Z0_t (Midori_rounds_SR_Result[13]), .Z0_f (new_AGEMA_signal_4379), .Z1_t (new_AGEMA_signal_4380), .Z1_f (new_AGEMA_signal_4381) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U16 ( .A0_t (Midori_rounds_roundReg_out[32]), .A0_f (new_AGEMA_signal_3021), .A1_t (new_AGEMA_signal_3022), .A1_f (new_AGEMA_signal_3023), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n10), .B0_f (new_AGEMA_signal_3015), .B1_t (new_AGEMA_signal_3016), .B1_f (new_AGEMA_signal_3017), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n11), .Z0_f (new_AGEMA_signal_3942), .Z1_t (new_AGEMA_signal_3943), .Z1_f (new_AGEMA_signal_3944) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U15 ( .A0_t (Midori_rounds_roundReg_out[35]), .A0_f (new_AGEMA_signal_3009), .A1_t (new_AGEMA_signal_3010), .A1_f (new_AGEMA_signal_3011), .B0_t (Midori_rounds_roundReg_out[34]), .B0_f (new_AGEMA_signal_3012), .B1_t (new_AGEMA_signal_3013), .B1_f (new_AGEMA_signal_3014), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n10), .Z0_f (new_AGEMA_signal_3015), .Z1_t (new_AGEMA_signal_3016), .Z1_f (new_AGEMA_signal_3017) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U14 ( .A0_t (Midori_rounds_roundReg_out[34]), .A0_f (new_AGEMA_signal_3012), .A1_t (new_AGEMA_signal_3013), .A1_f (new_AGEMA_signal_3014), .B0_t (Midori_rounds_roundReg_out[35]), .B0_f (new_AGEMA_signal_3009), .B1_t (new_AGEMA_signal_3010), .B1_f (new_AGEMA_signal_3011), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n12), .Z0_f (new_AGEMA_signal_3018), .Z1_t (new_AGEMA_signal_3019), .Z1_f (new_AGEMA_signal_3020) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n15), .A0_f (new_AGEMA_signal_3027), .A1_t (new_AGEMA_signal_3028), .A1_f (new_AGEMA_signal_3029), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n7), .B0_f (new_AGEMA_signal_4382), .B1_t (new_AGEMA_signal_4383), .B1_f (new_AGEMA_signal_4384), .Z0_t (Midori_rounds_SR_Result[14]), .Z0_f (new_AGEMA_signal_4730), .Z1_t (new_AGEMA_signal_4731), .Z1_f (new_AGEMA_signal_4732) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n6), .A0_f (new_AGEMA_signal_3945), .A1_t (new_AGEMA_signal_3946), .A1_f (new_AGEMA_signal_3947), .B0_t (Midori_rounds_roundReg_out[33]), .B0_f (new_AGEMA_signal_3936), .B1_t (new_AGEMA_signal_3937), .B1_f (new_AGEMA_signal_3938), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n7), .Z0_f (new_AGEMA_signal_4382), .Z1_t (new_AGEMA_signal_4383), .Z1_f (new_AGEMA_signal_4384) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n5), .A0_f (new_AGEMA_signal_3024), .A1_t (new_AGEMA_signal_3025), .A1_f (new_AGEMA_signal_3026), .B0_t (Midori_rounds_roundReg_out[34]), .B0_f (new_AGEMA_signal_3012), .B1_t (new_AGEMA_signal_3013), .B1_f (new_AGEMA_signal_3014), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n6), .Z0_f (new_AGEMA_signal_3945), .Z1_t (new_AGEMA_signal_3946), .Z1_f (new_AGEMA_signal_3947) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U10 ( .A0_t (Midori_rounds_roundReg_out[32]), .A0_f (new_AGEMA_signal_3021), .A1_t (new_AGEMA_signal_3022), .A1_f (new_AGEMA_signal_3023), .B0_t (Midori_rounds_roundReg_out[35]), .B0_f (new_AGEMA_signal_3009), .B1_t (new_AGEMA_signal_3010), .B1_f (new_AGEMA_signal_3011), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n5), .Z0_f (new_AGEMA_signal_3024), .Z1_t (new_AGEMA_signal_3025), .Z1_f (new_AGEMA_signal_3026) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U9 ( .A0_t (Midori_rounds_roundReg_out[35]), .A0_f (new_AGEMA_signal_3009), .A1_t (new_AGEMA_signal_3010), .A1_f (new_AGEMA_signal_3011), .B0_t (Midori_rounds_roundReg_out[32]), .B0_f (new_AGEMA_signal_3021), .B1_t (new_AGEMA_signal_3022), .B1_f (new_AGEMA_signal_3023), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n15), .Z0_f (new_AGEMA_signal_3027), .Z1_t (new_AGEMA_signal_3028), .Z1_f (new_AGEMA_signal_3029) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n13), .A0_f (new_AGEMA_signal_3033), .A1_t (new_AGEMA_signal_3034), .A1_f (new_AGEMA_signal_3035), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n3), .B0_f (new_AGEMA_signal_4385), .B1_t (new_AGEMA_signal_4386), .B1_f (new_AGEMA_signal_4387), .Z0_t (Midori_rounds_SR_Result[12]), .Z0_f (new_AGEMA_signal_4733), .Z1_t (new_AGEMA_signal_4734), .Z1_f (new_AGEMA_signal_4735) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U7 ( .A0_t (Midori_rounds_roundReg_out[33]), .A0_f (new_AGEMA_signal_3936), .A1_t (new_AGEMA_signal_3937), .A1_f (new_AGEMA_signal_3938), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n2), .B0_f (new_AGEMA_signal_3948), .B1_t (new_AGEMA_signal_3949), .B1_f (new_AGEMA_signal_3950), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n3), .Z0_f (new_AGEMA_signal_4385), .Z1_t (new_AGEMA_signal_4386), .Z1_f (new_AGEMA_signal_4387) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U6 ( .A0_t (Midori_rounds_roundReg_out[32]), .A0_f (new_AGEMA_signal_3021), .A1_t (new_AGEMA_signal_3022), .A1_f (new_AGEMA_signal_3023), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n1), .B0_f (new_AGEMA_signal_3030), .B1_t (new_AGEMA_signal_3031), .B1_f (new_AGEMA_signal_3032), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n2), .Z0_f (new_AGEMA_signal_3948), .Z1_t (new_AGEMA_signal_3949), .Z1_f (new_AGEMA_signal_3950) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U5 ( .A0_t (Midori_rounds_roundReg_out[34]), .A0_f (new_AGEMA_signal_3012), .A1_t (new_AGEMA_signal_3013), .A1_f (new_AGEMA_signal_3014), .B0_t (Midori_rounds_roundReg_out[35]), .B0_f (new_AGEMA_signal_3009), .B1_t (new_AGEMA_signal_3010), .B1_f (new_AGEMA_signal_3011), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n1), .Z0_f (new_AGEMA_signal_3030), .Z1_t (new_AGEMA_signal_3031), .Z1_f (new_AGEMA_signal_3032) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U3 ( .A0_t (Midori_rounds_roundReg_out[34]), .A0_f (new_AGEMA_signal_3012), .A1_t (new_AGEMA_signal_3013), .A1_f (new_AGEMA_signal_3014), .B0_t (Midori_rounds_roundReg_out[35]), .B0_f (new_AGEMA_signal_3009), .B1_t (new_AGEMA_signal_3010), .B1_f (new_AGEMA_signal_3011), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n13), .Z0_f (new_AGEMA_signal_3033), .Z1_t (new_AGEMA_signal_3034), .Z1_f (new_AGEMA_signal_3035) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n15), .A0_f (new_AGEMA_signal_3054), .A1_t (new_AGEMA_signal_3055), .A1_f (new_AGEMA_signal_3056), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n14), .B0_f (new_AGEMA_signal_3954), .B1_t (new_AGEMA_signal_3955), .B1_f (new_AGEMA_signal_3956), .Z0_t (Midori_rounds_SR_Result[19]), .Z0_f (new_AGEMA_signal_4388), .Z1_t (new_AGEMA_signal_4389), .Z1_f (new_AGEMA_signal_4390) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n13), .A0_f (new_AGEMA_signal_3060), .A1_t (new_AGEMA_signal_3061), .A1_f (new_AGEMA_signal_3062), .B0_t (Midori_rounds_roundReg_out[37]), .B0_f (new_AGEMA_signal_3951), .B1_t (new_AGEMA_signal_3952), .B1_f (new_AGEMA_signal_3953), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n14), .Z0_f (new_AGEMA_signal_3954), .Z1_t (new_AGEMA_signal_3955), .Z1_f (new_AGEMA_signal_3956) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n12), .A0_f (new_AGEMA_signal_3045), .A1_t (new_AGEMA_signal_3046), .A1_f (new_AGEMA_signal_3047), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n11), .B0_f (new_AGEMA_signal_3957), .B1_t (new_AGEMA_signal_3958), .B1_f (new_AGEMA_signal_3959), .Z0_t (Midori_rounds_SR_Result[17]), .Z0_f (new_AGEMA_signal_4391), .Z1_t (new_AGEMA_signal_4392), .Z1_f (new_AGEMA_signal_4393) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U16 ( .A0_t (Midori_rounds_roundReg_out[36]), .A0_f (new_AGEMA_signal_3048), .A1_t (new_AGEMA_signal_3049), .A1_f (new_AGEMA_signal_3050), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n10), .B0_f (new_AGEMA_signal_3042), .B1_t (new_AGEMA_signal_3043), .B1_f (new_AGEMA_signal_3044), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n11), .Z0_f (new_AGEMA_signal_3957), .Z1_t (new_AGEMA_signal_3958), .Z1_f (new_AGEMA_signal_3959) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U15 ( .A0_t (Midori_rounds_roundReg_out[39]), .A0_f (new_AGEMA_signal_3036), .A1_t (new_AGEMA_signal_3037), .A1_f (new_AGEMA_signal_3038), .B0_t (Midori_rounds_roundReg_out[38]), .B0_f (new_AGEMA_signal_3039), .B1_t (new_AGEMA_signal_3040), .B1_f (new_AGEMA_signal_3041), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n10), .Z0_f (new_AGEMA_signal_3042), .Z1_t (new_AGEMA_signal_3043), .Z1_f (new_AGEMA_signal_3044) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U14 ( .A0_t (Midori_rounds_roundReg_out[38]), .A0_f (new_AGEMA_signal_3039), .A1_t (new_AGEMA_signal_3040), .A1_f (new_AGEMA_signal_3041), .B0_t (Midori_rounds_roundReg_out[39]), .B0_f (new_AGEMA_signal_3036), .B1_t (new_AGEMA_signal_3037), .B1_f (new_AGEMA_signal_3038), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n12), .Z0_f (new_AGEMA_signal_3045), .Z1_t (new_AGEMA_signal_3046), .Z1_f (new_AGEMA_signal_3047) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n15), .A0_f (new_AGEMA_signal_3054), .A1_t (new_AGEMA_signal_3055), .A1_f (new_AGEMA_signal_3056), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n7), .B0_f (new_AGEMA_signal_4394), .B1_t (new_AGEMA_signal_4395), .B1_f (new_AGEMA_signal_4396), .Z0_t (Midori_rounds_SR_Result[18]), .Z0_f (new_AGEMA_signal_4736), .Z1_t (new_AGEMA_signal_4737), .Z1_f (new_AGEMA_signal_4738) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n6), .A0_f (new_AGEMA_signal_3960), .A1_t (new_AGEMA_signal_3961), .A1_f (new_AGEMA_signal_3962), .B0_t (Midori_rounds_roundReg_out[37]), .B0_f (new_AGEMA_signal_3951), .B1_t (new_AGEMA_signal_3952), .B1_f (new_AGEMA_signal_3953), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n7), .Z0_f (new_AGEMA_signal_4394), .Z1_t (new_AGEMA_signal_4395), .Z1_f (new_AGEMA_signal_4396) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n5), .A0_f (new_AGEMA_signal_3051), .A1_t (new_AGEMA_signal_3052), .A1_f (new_AGEMA_signal_3053), .B0_t (Midori_rounds_roundReg_out[38]), .B0_f (new_AGEMA_signal_3039), .B1_t (new_AGEMA_signal_3040), .B1_f (new_AGEMA_signal_3041), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n6), .Z0_f (new_AGEMA_signal_3960), .Z1_t (new_AGEMA_signal_3961), .Z1_f (new_AGEMA_signal_3962) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U10 ( .A0_t (Midori_rounds_roundReg_out[36]), .A0_f (new_AGEMA_signal_3048), .A1_t (new_AGEMA_signal_3049), .A1_f (new_AGEMA_signal_3050), .B0_t (Midori_rounds_roundReg_out[39]), .B0_f (new_AGEMA_signal_3036), .B1_t (new_AGEMA_signal_3037), .B1_f (new_AGEMA_signal_3038), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n5), .Z0_f (new_AGEMA_signal_3051), .Z1_t (new_AGEMA_signal_3052), .Z1_f (new_AGEMA_signal_3053) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U9 ( .A0_t (Midori_rounds_roundReg_out[39]), .A0_f (new_AGEMA_signal_3036), .A1_t (new_AGEMA_signal_3037), .A1_f (new_AGEMA_signal_3038), .B0_t (Midori_rounds_roundReg_out[36]), .B0_f (new_AGEMA_signal_3048), .B1_t (new_AGEMA_signal_3049), .B1_f (new_AGEMA_signal_3050), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n15), .Z0_f (new_AGEMA_signal_3054), .Z1_t (new_AGEMA_signal_3055), .Z1_f (new_AGEMA_signal_3056) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n13), .A0_f (new_AGEMA_signal_3060), .A1_t (new_AGEMA_signal_3061), .A1_f (new_AGEMA_signal_3062), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n3), .B0_f (new_AGEMA_signal_4397), .B1_t (new_AGEMA_signal_4398), .B1_f (new_AGEMA_signal_4399), .Z0_t (Midori_rounds_SR_Result[16]), .Z0_f (new_AGEMA_signal_4739), .Z1_t (new_AGEMA_signal_4740), .Z1_f (new_AGEMA_signal_4741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U7 ( .A0_t (Midori_rounds_roundReg_out[37]), .A0_f (new_AGEMA_signal_3951), .A1_t (new_AGEMA_signal_3952), .A1_f (new_AGEMA_signal_3953), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n2), .B0_f (new_AGEMA_signal_3963), .B1_t (new_AGEMA_signal_3964), .B1_f (new_AGEMA_signal_3965), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n3), .Z0_f (new_AGEMA_signal_4397), .Z1_t (new_AGEMA_signal_4398), .Z1_f (new_AGEMA_signal_4399) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U6 ( .A0_t (Midori_rounds_roundReg_out[36]), .A0_f (new_AGEMA_signal_3048), .A1_t (new_AGEMA_signal_3049), .A1_f (new_AGEMA_signal_3050), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n1), .B0_f (new_AGEMA_signal_3057), .B1_t (new_AGEMA_signal_3058), .B1_f (new_AGEMA_signal_3059), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n2), .Z0_f (new_AGEMA_signal_3963), .Z1_t (new_AGEMA_signal_3964), .Z1_f (new_AGEMA_signal_3965) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U5 ( .A0_t (Midori_rounds_roundReg_out[38]), .A0_f (new_AGEMA_signal_3039), .A1_t (new_AGEMA_signal_3040), .A1_f (new_AGEMA_signal_3041), .B0_t (Midori_rounds_roundReg_out[39]), .B0_f (new_AGEMA_signal_3036), .B1_t (new_AGEMA_signal_3037), .B1_f (new_AGEMA_signal_3038), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n1), .Z0_f (new_AGEMA_signal_3057), .Z1_t (new_AGEMA_signal_3058), .Z1_f (new_AGEMA_signal_3059) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U3 ( .A0_t (Midori_rounds_roundReg_out[38]), .A0_f (new_AGEMA_signal_3039), .A1_t (new_AGEMA_signal_3040), .A1_f (new_AGEMA_signal_3041), .B0_t (Midori_rounds_roundReg_out[39]), .B0_f (new_AGEMA_signal_3036), .B1_t (new_AGEMA_signal_3037), .B1_f (new_AGEMA_signal_3038), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n13), .Z0_f (new_AGEMA_signal_3060), .Z1_t (new_AGEMA_signal_3061), .Z1_f (new_AGEMA_signal_3062) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n15), .A0_f (new_AGEMA_signal_4400), .A1_t (new_AGEMA_signal_4401), .A1_f (new_AGEMA_signal_4402), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n14), .B0_f (new_AGEMA_signal_3078), .B1_t (new_AGEMA_signal_3079), .B1_f (new_AGEMA_signal_3080), .Z0_t (Midori_rounds_SR_Result[52]), .Z0_f (new_AGEMA_signal_4742), .Z1_t (new_AGEMA_signal_4743), .Z1_f (new_AGEMA_signal_4744) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U18 ( .A0_t (Midori_rounds_roundReg_out[41]), .A0_f (new_AGEMA_signal_3972), .A1_t (new_AGEMA_signal_3973), .A1_f (new_AGEMA_signal_3974), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n13), .B0_f (new_AGEMA_signal_3966), .B1_t (new_AGEMA_signal_3967), .B1_f (new_AGEMA_signal_3968), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n15), .Z0_f (new_AGEMA_signal_4400), .Z1_t (new_AGEMA_signal_4401), .Z1_f (new_AGEMA_signal_4402) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U17 ( .A0_t (Midori_rounds_roundReg_out[40]), .A0_f (new_AGEMA_signal_3072), .A1_t (new_AGEMA_signal_3073), .A1_f (new_AGEMA_signal_3074), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n11), .B0_f (new_AGEMA_signal_3069), .B1_t (new_AGEMA_signal_3070), .B1_f (new_AGEMA_signal_3071), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n13), .Z0_f (new_AGEMA_signal_3966), .Z1_t (new_AGEMA_signal_3967), .Z1_f (new_AGEMA_signal_3968) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U16 ( .A0_t (Midori_rounds_roundReg_out[42]), .A0_f (new_AGEMA_signal_3063), .A1_t (new_AGEMA_signal_3064), .A1_f (new_AGEMA_signal_3065), .B0_t (Midori_rounds_roundReg_out[43]), .B0_f (new_AGEMA_signal_3066), .B1_t (new_AGEMA_signal_3067), .B1_f (new_AGEMA_signal_3068), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n11), .Z0_f (new_AGEMA_signal_3069), .Z1_t (new_AGEMA_signal_3070), .Z1_f (new_AGEMA_signal_3071) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n10), .A0_f (new_AGEMA_signal_4403), .A1_t (new_AGEMA_signal_4404), .A1_f (new_AGEMA_signal_4405), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n9), .B0_f (new_AGEMA_signal_3081), .B1_t (new_AGEMA_signal_3082), .B1_f (new_AGEMA_signal_3083), .Z0_t (Midori_rounds_SR_Result[54]), .Z0_f (new_AGEMA_signal_4745), .Z1_t (new_AGEMA_signal_4746), .Z1_f (new_AGEMA_signal_4747) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n8), .A0_f (new_AGEMA_signal_3969), .A1_t (new_AGEMA_signal_3970), .A1_f (new_AGEMA_signal_3971), .B0_t (Midori_rounds_roundReg_out[41]), .B0_f (new_AGEMA_signal_3972), .B1_t (new_AGEMA_signal_3973), .B1_f (new_AGEMA_signal_3974), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n10), .Z0_f (new_AGEMA_signal_4403), .Z1_t (new_AGEMA_signal_4404), .Z1_f (new_AGEMA_signal_4405) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n7), .A0_f (new_AGEMA_signal_3075), .A1_t (new_AGEMA_signal_3076), .A1_f (new_AGEMA_signal_3077), .B0_t (Midori_rounds_roundReg_out[42]), .B0_f (new_AGEMA_signal_3063), .B1_t (new_AGEMA_signal_3064), .B1_f (new_AGEMA_signal_3065), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n8), .Z0_f (new_AGEMA_signal_3969), .Z1_t (new_AGEMA_signal_3970), .Z1_f (new_AGEMA_signal_3971) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U12 ( .A0_t (Midori_rounds_roundReg_out[40]), .A0_f (new_AGEMA_signal_3072), .A1_t (new_AGEMA_signal_3073), .A1_f (new_AGEMA_signal_3074), .B0_t (Midori_rounds_roundReg_out[43]), .B0_f (new_AGEMA_signal_3066), .B1_t (new_AGEMA_signal_3067), .B1_f (new_AGEMA_signal_3068), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n7), .Z0_f (new_AGEMA_signal_3075), .Z1_t (new_AGEMA_signal_3076), .Z1_f (new_AGEMA_signal_3077) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n9), .A0_f (new_AGEMA_signal_3081), .A1_t (new_AGEMA_signal_3082), .A1_f (new_AGEMA_signal_3083), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n5), .B0_f (new_AGEMA_signal_3975), .B1_t (new_AGEMA_signal_3976), .B1_f (new_AGEMA_signal_3977), .Z0_t (Midori_rounds_SR_Result[55]), .Z0_f (new_AGEMA_signal_4406), .Z1_t (new_AGEMA_signal_4407), .Z1_f (new_AGEMA_signal_4408) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U10 ( .A0_t (Midori_rounds_roundReg_out[41]), .A0_f (new_AGEMA_signal_3972), .A1_t (new_AGEMA_signal_3973), .A1_f (new_AGEMA_signal_3974), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n14), .B0_f (new_AGEMA_signal_3078), .B1_t (new_AGEMA_signal_3079), .B1_f (new_AGEMA_signal_3080), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n5), .Z0_f (new_AGEMA_signal_3975), .Z1_t (new_AGEMA_signal_3976), .Z1_f (new_AGEMA_signal_3977) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U9 ( .A0_t (Midori_rounds_roundReg_out[42]), .A0_f (new_AGEMA_signal_3063), .A1_t (new_AGEMA_signal_3064), .A1_f (new_AGEMA_signal_3065), .B0_t (Midori_rounds_roundReg_out[43]), .B0_f (new_AGEMA_signal_3066), .B1_t (new_AGEMA_signal_3067), .B1_f (new_AGEMA_signal_3068), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n14), .Z0_f (new_AGEMA_signal_3078), .Z1_t (new_AGEMA_signal_3079), .Z1_f (new_AGEMA_signal_3080) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U8 ( .A0_t (Midori_rounds_roundReg_out[43]), .A0_f (new_AGEMA_signal_3066), .A1_t (new_AGEMA_signal_3067), .A1_f (new_AGEMA_signal_3068), .B0_t (Midori_rounds_roundReg_out[40]), .B0_f (new_AGEMA_signal_3072), .B1_t (new_AGEMA_signal_3073), .B1_f (new_AGEMA_signal_3074), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n9), .Z0_f (new_AGEMA_signal_3081), .Z1_t (new_AGEMA_signal_3082), .Z1_f (new_AGEMA_signal_3083) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n3), .A0_f (new_AGEMA_signal_3087), .A1_t (new_AGEMA_signal_3088), .A1_f (new_AGEMA_signal_3089), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n2), .B0_f (new_AGEMA_signal_3978), .B1_t (new_AGEMA_signal_3979), .B1_f (new_AGEMA_signal_3980), .Z0_t (Midori_rounds_SR_Result[53]), .Z0_f (new_AGEMA_signal_4409), .Z1_t (new_AGEMA_signal_4410), .Z1_f (new_AGEMA_signal_4411) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n1), .A0_f (new_AGEMA_signal_3084), .A1_t (new_AGEMA_signal_3085), .A1_f (new_AGEMA_signal_3086), .B0_t (Midori_rounds_roundReg_out[43]), .B0_f (new_AGEMA_signal_3066), .B1_t (new_AGEMA_signal_3067), .B1_f (new_AGEMA_signal_3068), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n2), .Z0_f (new_AGEMA_signal_3978), .Z1_t (new_AGEMA_signal_3979), .Z1_f (new_AGEMA_signal_3980) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U4 ( .A0_t (Midori_rounds_roundReg_out[42]), .A0_f (new_AGEMA_signal_3063), .A1_t (new_AGEMA_signal_3064), .A1_f (new_AGEMA_signal_3065), .B0_t (Midori_rounds_roundReg_out[40]), .B0_f (new_AGEMA_signal_3072), .B1_t (new_AGEMA_signal_3073), .B1_f (new_AGEMA_signal_3074), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n1), .Z0_f (new_AGEMA_signal_3084), .Z1_t (new_AGEMA_signal_3085), .Z1_f (new_AGEMA_signal_3086) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U1 ( .A0_t (Midori_rounds_roundReg_out[42]), .A0_f (new_AGEMA_signal_3063), .A1_t (new_AGEMA_signal_3064), .A1_f (new_AGEMA_signal_3065), .B0_t (Midori_rounds_roundReg_out[40]), .B0_f (new_AGEMA_signal_3072), .B1_t (new_AGEMA_signal_3073), .B1_f (new_AGEMA_signal_3074), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n3), .Z0_f (new_AGEMA_signal_3087), .Z1_t (new_AGEMA_signal_3088), .Z1_f (new_AGEMA_signal_3089) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n15), .A0_f (new_AGEMA_signal_4412), .A1_t (new_AGEMA_signal_4413), .A1_f (new_AGEMA_signal_4414), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n14), .B0_f (new_AGEMA_signal_3105), .B1_t (new_AGEMA_signal_3106), .B1_f (new_AGEMA_signal_3107), .Z0_t (Midori_rounds_SR_Result[40]), .Z0_f (new_AGEMA_signal_4748), .Z1_t (new_AGEMA_signal_4749), .Z1_f (new_AGEMA_signal_4750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U18 ( .A0_t (Midori_rounds_roundReg_out[45]), .A0_f (new_AGEMA_signal_3987), .A1_t (new_AGEMA_signal_3988), .A1_f (new_AGEMA_signal_3989), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n13), .B0_f (new_AGEMA_signal_3981), .B1_t (new_AGEMA_signal_3982), .B1_f (new_AGEMA_signal_3983), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n15), .Z0_f (new_AGEMA_signal_4412), .Z1_t (new_AGEMA_signal_4413), .Z1_f (new_AGEMA_signal_4414) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U17 ( .A0_t (Midori_rounds_roundReg_out[44]), .A0_f (new_AGEMA_signal_3099), .A1_t (new_AGEMA_signal_3100), .A1_f (new_AGEMA_signal_3101), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n11), .B0_f (new_AGEMA_signal_3096), .B1_t (new_AGEMA_signal_3097), .B1_f (new_AGEMA_signal_3098), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n13), .Z0_f (new_AGEMA_signal_3981), .Z1_t (new_AGEMA_signal_3982), .Z1_f (new_AGEMA_signal_3983) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U16 ( .A0_t (Midori_rounds_roundReg_out[46]), .A0_f (new_AGEMA_signal_3090), .A1_t (new_AGEMA_signal_3091), .A1_f (new_AGEMA_signal_3092), .B0_t (Midori_rounds_roundReg_out[47]), .B0_f (new_AGEMA_signal_3093), .B1_t (new_AGEMA_signal_3094), .B1_f (new_AGEMA_signal_3095), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n11), .Z0_f (new_AGEMA_signal_3096), .Z1_t (new_AGEMA_signal_3097), .Z1_f (new_AGEMA_signal_3098) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n10), .A0_f (new_AGEMA_signal_4415), .A1_t (new_AGEMA_signal_4416), .A1_f (new_AGEMA_signal_4417), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n9), .B0_f (new_AGEMA_signal_3108), .B1_t (new_AGEMA_signal_3109), .B1_f (new_AGEMA_signal_3110), .Z0_t (Midori_rounds_SR_Result[42]), .Z0_f (new_AGEMA_signal_4751), .Z1_t (new_AGEMA_signal_4752), .Z1_f (new_AGEMA_signal_4753) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n8), .A0_f (new_AGEMA_signal_3984), .A1_t (new_AGEMA_signal_3985), .A1_f (new_AGEMA_signal_3986), .B0_t (Midori_rounds_roundReg_out[45]), .B0_f (new_AGEMA_signal_3987), .B1_t (new_AGEMA_signal_3988), .B1_f (new_AGEMA_signal_3989), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n10), .Z0_f (new_AGEMA_signal_4415), .Z1_t (new_AGEMA_signal_4416), .Z1_f (new_AGEMA_signal_4417) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n7), .A0_f (new_AGEMA_signal_3102), .A1_t (new_AGEMA_signal_3103), .A1_f (new_AGEMA_signal_3104), .B0_t (Midori_rounds_roundReg_out[46]), .B0_f (new_AGEMA_signal_3090), .B1_t (new_AGEMA_signal_3091), .B1_f (new_AGEMA_signal_3092), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n8), .Z0_f (new_AGEMA_signal_3984), .Z1_t (new_AGEMA_signal_3985), .Z1_f (new_AGEMA_signal_3986) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U12 ( .A0_t (Midori_rounds_roundReg_out[44]), .A0_f (new_AGEMA_signal_3099), .A1_t (new_AGEMA_signal_3100), .A1_f (new_AGEMA_signal_3101), .B0_t (Midori_rounds_roundReg_out[47]), .B0_f (new_AGEMA_signal_3093), .B1_t (new_AGEMA_signal_3094), .B1_f (new_AGEMA_signal_3095), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n7), .Z0_f (new_AGEMA_signal_3102), .Z1_t (new_AGEMA_signal_3103), .Z1_f (new_AGEMA_signal_3104) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n9), .A0_f (new_AGEMA_signal_3108), .A1_t (new_AGEMA_signal_3109), .A1_f (new_AGEMA_signal_3110), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n5), .B0_f (new_AGEMA_signal_3990), .B1_t (new_AGEMA_signal_3991), .B1_f (new_AGEMA_signal_3992), .Z0_t (Midori_rounds_SR_Result[43]), .Z0_f (new_AGEMA_signal_4418), .Z1_t (new_AGEMA_signal_4419), .Z1_f (new_AGEMA_signal_4420) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U10 ( .A0_t (Midori_rounds_roundReg_out[45]), .A0_f (new_AGEMA_signal_3987), .A1_t (new_AGEMA_signal_3988), .A1_f (new_AGEMA_signal_3989), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n14), .B0_f (new_AGEMA_signal_3105), .B1_t (new_AGEMA_signal_3106), .B1_f (new_AGEMA_signal_3107), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n5), .Z0_f (new_AGEMA_signal_3990), .Z1_t (new_AGEMA_signal_3991), .Z1_f (new_AGEMA_signal_3992) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U9 ( .A0_t (Midori_rounds_roundReg_out[46]), .A0_f (new_AGEMA_signal_3090), .A1_t (new_AGEMA_signal_3091), .A1_f (new_AGEMA_signal_3092), .B0_t (Midori_rounds_roundReg_out[47]), .B0_f (new_AGEMA_signal_3093), .B1_t (new_AGEMA_signal_3094), .B1_f (new_AGEMA_signal_3095), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n14), .Z0_f (new_AGEMA_signal_3105), .Z1_t (new_AGEMA_signal_3106), .Z1_f (new_AGEMA_signal_3107) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U8 ( .A0_t (Midori_rounds_roundReg_out[47]), .A0_f (new_AGEMA_signal_3093), .A1_t (new_AGEMA_signal_3094), .A1_f (new_AGEMA_signal_3095), .B0_t (Midori_rounds_roundReg_out[44]), .B0_f (new_AGEMA_signal_3099), .B1_t (new_AGEMA_signal_3100), .B1_f (new_AGEMA_signal_3101), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n9), .Z0_f (new_AGEMA_signal_3108), .Z1_t (new_AGEMA_signal_3109), .Z1_f (new_AGEMA_signal_3110) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n3), .A0_f (new_AGEMA_signal_3114), .A1_t (new_AGEMA_signal_3115), .A1_f (new_AGEMA_signal_3116), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n2), .B0_f (new_AGEMA_signal_3993), .B1_t (new_AGEMA_signal_3994), .B1_f (new_AGEMA_signal_3995), .Z0_t (Midori_rounds_SR_Result[41]), .Z0_f (new_AGEMA_signal_4421), .Z1_t (new_AGEMA_signal_4422), .Z1_f (new_AGEMA_signal_4423) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n1), .A0_f (new_AGEMA_signal_3111), .A1_t (new_AGEMA_signal_3112), .A1_f (new_AGEMA_signal_3113), .B0_t (Midori_rounds_roundReg_out[47]), .B0_f (new_AGEMA_signal_3093), .B1_t (new_AGEMA_signal_3094), .B1_f (new_AGEMA_signal_3095), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n2), .Z0_f (new_AGEMA_signal_3993), .Z1_t (new_AGEMA_signal_3994), .Z1_f (new_AGEMA_signal_3995) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U4 ( .A0_t (Midori_rounds_roundReg_out[46]), .A0_f (new_AGEMA_signal_3090), .A1_t (new_AGEMA_signal_3091), .A1_f (new_AGEMA_signal_3092), .B0_t (Midori_rounds_roundReg_out[44]), .B0_f (new_AGEMA_signal_3099), .B1_t (new_AGEMA_signal_3100), .B1_f (new_AGEMA_signal_3101), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n1), .Z0_f (new_AGEMA_signal_3111), .Z1_t (new_AGEMA_signal_3112), .Z1_f (new_AGEMA_signal_3113) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U1 ( .A0_t (Midori_rounds_roundReg_out[46]), .A0_f (new_AGEMA_signal_3090), .A1_t (new_AGEMA_signal_3091), .A1_f (new_AGEMA_signal_3092), .B0_t (Midori_rounds_roundReg_out[44]), .B0_f (new_AGEMA_signal_3099), .B1_t (new_AGEMA_signal_3100), .B1_f (new_AGEMA_signal_3101), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n3), .Z0_f (new_AGEMA_signal_3114), .Z1_t (new_AGEMA_signal_3115), .Z1_f (new_AGEMA_signal_3116) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n15), .A0_f (new_AGEMA_signal_4424), .A1_t (new_AGEMA_signal_4425), .A1_f (new_AGEMA_signal_4426), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n14), .B0_f (new_AGEMA_signal_3132), .B1_t (new_AGEMA_signal_3133), .B1_f (new_AGEMA_signal_3134), .Z0_t (Midori_rounds_SR_Result[24]), .Z0_f (new_AGEMA_signal_4754), .Z1_t (new_AGEMA_signal_4755), .Z1_f (new_AGEMA_signal_4756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U18 ( .A0_t (Midori_rounds_roundReg_out[49]), .A0_f (new_AGEMA_signal_4002), .A1_t (new_AGEMA_signal_4003), .A1_f (new_AGEMA_signal_4004), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n13), .B0_f (new_AGEMA_signal_3996), .B1_t (new_AGEMA_signal_3997), .B1_f (new_AGEMA_signal_3998), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n15), .Z0_f (new_AGEMA_signal_4424), .Z1_t (new_AGEMA_signal_4425), .Z1_f (new_AGEMA_signal_4426) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U17 ( .A0_t (Midori_rounds_roundReg_out[48]), .A0_f (new_AGEMA_signal_3126), .A1_t (new_AGEMA_signal_3127), .A1_f (new_AGEMA_signal_3128), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n11), .B0_f (new_AGEMA_signal_3123), .B1_t (new_AGEMA_signal_3124), .B1_f (new_AGEMA_signal_3125), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n13), .Z0_f (new_AGEMA_signal_3996), .Z1_t (new_AGEMA_signal_3997), .Z1_f (new_AGEMA_signal_3998) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U16 ( .A0_t (Midori_rounds_roundReg_out[50]), .A0_f (new_AGEMA_signal_3117), .A1_t (new_AGEMA_signal_3118), .A1_f (new_AGEMA_signal_3119), .B0_t (Midori_rounds_roundReg_out[51]), .B0_f (new_AGEMA_signal_3120), .B1_t (new_AGEMA_signal_3121), .B1_f (new_AGEMA_signal_3122), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n11), .Z0_f (new_AGEMA_signal_3123), .Z1_t (new_AGEMA_signal_3124), .Z1_f (new_AGEMA_signal_3125) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n10), .A0_f (new_AGEMA_signal_4427), .A1_t (new_AGEMA_signal_4428), .A1_f (new_AGEMA_signal_4429), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n9), .B0_f (new_AGEMA_signal_3135), .B1_t (new_AGEMA_signal_3136), .B1_f (new_AGEMA_signal_3137), .Z0_t (Midori_rounds_SR_Result[26]), .Z0_f (new_AGEMA_signal_4757), .Z1_t (new_AGEMA_signal_4758), .Z1_f (new_AGEMA_signal_4759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n8), .A0_f (new_AGEMA_signal_3999), .A1_t (new_AGEMA_signal_4000), .A1_f (new_AGEMA_signal_4001), .B0_t (Midori_rounds_roundReg_out[49]), .B0_f (new_AGEMA_signal_4002), .B1_t (new_AGEMA_signal_4003), .B1_f (new_AGEMA_signal_4004), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n10), .Z0_f (new_AGEMA_signal_4427), .Z1_t (new_AGEMA_signal_4428), .Z1_f (new_AGEMA_signal_4429) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n7), .A0_f (new_AGEMA_signal_3129), .A1_t (new_AGEMA_signal_3130), .A1_f (new_AGEMA_signal_3131), .B0_t (Midori_rounds_roundReg_out[50]), .B0_f (new_AGEMA_signal_3117), .B1_t (new_AGEMA_signal_3118), .B1_f (new_AGEMA_signal_3119), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n8), .Z0_f (new_AGEMA_signal_3999), .Z1_t (new_AGEMA_signal_4000), .Z1_f (new_AGEMA_signal_4001) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U12 ( .A0_t (Midori_rounds_roundReg_out[48]), .A0_f (new_AGEMA_signal_3126), .A1_t (new_AGEMA_signal_3127), .A1_f (new_AGEMA_signal_3128), .B0_t (Midori_rounds_roundReg_out[51]), .B0_f (new_AGEMA_signal_3120), .B1_t (new_AGEMA_signal_3121), .B1_f (new_AGEMA_signal_3122), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n7), .Z0_f (new_AGEMA_signal_3129), .Z1_t (new_AGEMA_signal_3130), .Z1_f (new_AGEMA_signal_3131) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n9), .A0_f (new_AGEMA_signal_3135), .A1_t (new_AGEMA_signal_3136), .A1_f (new_AGEMA_signal_3137), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n5), .B0_f (new_AGEMA_signal_4005), .B1_t (new_AGEMA_signal_4006), .B1_f (new_AGEMA_signal_4007), .Z0_t (Midori_rounds_SR_Result[27]), .Z0_f (new_AGEMA_signal_4430), .Z1_t (new_AGEMA_signal_4431), .Z1_f (new_AGEMA_signal_4432) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U10 ( .A0_t (Midori_rounds_roundReg_out[49]), .A0_f (new_AGEMA_signal_4002), .A1_t (new_AGEMA_signal_4003), .A1_f (new_AGEMA_signal_4004), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n14), .B0_f (new_AGEMA_signal_3132), .B1_t (new_AGEMA_signal_3133), .B1_f (new_AGEMA_signal_3134), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n5), .Z0_f (new_AGEMA_signal_4005), .Z1_t (new_AGEMA_signal_4006), .Z1_f (new_AGEMA_signal_4007) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U9 ( .A0_t (Midori_rounds_roundReg_out[50]), .A0_f (new_AGEMA_signal_3117), .A1_t (new_AGEMA_signal_3118), .A1_f (new_AGEMA_signal_3119), .B0_t (Midori_rounds_roundReg_out[51]), .B0_f (new_AGEMA_signal_3120), .B1_t (new_AGEMA_signal_3121), .B1_f (new_AGEMA_signal_3122), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n14), .Z0_f (new_AGEMA_signal_3132), .Z1_t (new_AGEMA_signal_3133), .Z1_f (new_AGEMA_signal_3134) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U8 ( .A0_t (Midori_rounds_roundReg_out[51]), .A0_f (new_AGEMA_signal_3120), .A1_t (new_AGEMA_signal_3121), .A1_f (new_AGEMA_signal_3122), .B0_t (Midori_rounds_roundReg_out[48]), .B0_f (new_AGEMA_signal_3126), .B1_t (new_AGEMA_signal_3127), .B1_f (new_AGEMA_signal_3128), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n9), .Z0_f (new_AGEMA_signal_3135), .Z1_t (new_AGEMA_signal_3136), .Z1_f (new_AGEMA_signal_3137) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n3), .A0_f (new_AGEMA_signal_3141), .A1_t (new_AGEMA_signal_3142), .A1_f (new_AGEMA_signal_3143), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n2), .B0_f (new_AGEMA_signal_4008), .B1_t (new_AGEMA_signal_4009), .B1_f (new_AGEMA_signal_4010), .Z0_t (Midori_rounds_SR_Result[25]), .Z0_f (new_AGEMA_signal_4433), .Z1_t (new_AGEMA_signal_4434), .Z1_f (new_AGEMA_signal_4435) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n1), .A0_f (new_AGEMA_signal_3138), .A1_t (new_AGEMA_signal_3139), .A1_f (new_AGEMA_signal_3140), .B0_t (Midori_rounds_roundReg_out[51]), .B0_f (new_AGEMA_signal_3120), .B1_t (new_AGEMA_signal_3121), .B1_f (new_AGEMA_signal_3122), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n2), .Z0_f (new_AGEMA_signal_4008), .Z1_t (new_AGEMA_signal_4009), .Z1_f (new_AGEMA_signal_4010) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U4 ( .A0_t (Midori_rounds_roundReg_out[50]), .A0_f (new_AGEMA_signal_3117), .A1_t (new_AGEMA_signal_3118), .A1_f (new_AGEMA_signal_3119), .B0_t (Midori_rounds_roundReg_out[48]), .B0_f (new_AGEMA_signal_3126), .B1_t (new_AGEMA_signal_3127), .B1_f (new_AGEMA_signal_3128), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n1), .Z0_f (new_AGEMA_signal_3138), .Z1_t (new_AGEMA_signal_3139), .Z1_f (new_AGEMA_signal_3140) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U1 ( .A0_t (Midori_rounds_roundReg_out[50]), .A0_f (new_AGEMA_signal_3117), .A1_t (new_AGEMA_signal_3118), .A1_f (new_AGEMA_signal_3119), .B0_t (Midori_rounds_roundReg_out[48]), .B0_f (new_AGEMA_signal_3126), .B1_t (new_AGEMA_signal_3127), .B1_f (new_AGEMA_signal_3128), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n3), .Z0_f (new_AGEMA_signal_3141), .Z1_t (new_AGEMA_signal_3142), .Z1_f (new_AGEMA_signal_3143) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n15), .A0_f (new_AGEMA_signal_3162), .A1_t (new_AGEMA_signal_3163), .A1_f (new_AGEMA_signal_3164), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n14), .B0_f (new_AGEMA_signal_4014), .B1_t (new_AGEMA_signal_4015), .B1_f (new_AGEMA_signal_4016), .Z0_t (Midori_rounds_SR_Result[7]), .Z0_f (new_AGEMA_signal_4436), .Z1_t (new_AGEMA_signal_4437), .Z1_f (new_AGEMA_signal_4438) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n13), .A0_f (new_AGEMA_signal_3168), .A1_t (new_AGEMA_signal_3169), .A1_f (new_AGEMA_signal_3170), .B0_t (Midori_rounds_roundReg_out[53]), .B0_f (new_AGEMA_signal_4011), .B1_t (new_AGEMA_signal_4012), .B1_f (new_AGEMA_signal_4013), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n14), .Z0_f (new_AGEMA_signal_4014), .Z1_t (new_AGEMA_signal_4015), .Z1_f (new_AGEMA_signal_4016) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n12), .A0_f (new_AGEMA_signal_3153), .A1_t (new_AGEMA_signal_3154), .A1_f (new_AGEMA_signal_3155), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n11), .B0_f (new_AGEMA_signal_4017), .B1_t (new_AGEMA_signal_4018), .B1_f (new_AGEMA_signal_4019), .Z0_t (Midori_rounds_SR_Result[5]), .Z0_f (new_AGEMA_signal_4439), .Z1_t (new_AGEMA_signal_4440), .Z1_f (new_AGEMA_signal_4441) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U16 ( .A0_t (Midori_rounds_roundReg_out[52]), .A0_f (new_AGEMA_signal_3156), .A1_t (new_AGEMA_signal_3157), .A1_f (new_AGEMA_signal_3158), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n10), .B0_f (new_AGEMA_signal_3150), .B1_t (new_AGEMA_signal_3151), .B1_f (new_AGEMA_signal_3152), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n11), .Z0_f (new_AGEMA_signal_4017), .Z1_t (new_AGEMA_signal_4018), .Z1_f (new_AGEMA_signal_4019) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U15 ( .A0_t (Midori_rounds_roundReg_out[55]), .A0_f (new_AGEMA_signal_3144), .A1_t (new_AGEMA_signal_3145), .A1_f (new_AGEMA_signal_3146), .B0_t (Midori_rounds_roundReg_out[54]), .B0_f (new_AGEMA_signal_3147), .B1_t (new_AGEMA_signal_3148), .B1_f (new_AGEMA_signal_3149), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n10), .Z0_f (new_AGEMA_signal_3150), .Z1_t (new_AGEMA_signal_3151), .Z1_f (new_AGEMA_signal_3152) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U14 ( .A0_t (Midori_rounds_roundReg_out[54]), .A0_f (new_AGEMA_signal_3147), .A1_t (new_AGEMA_signal_3148), .A1_f (new_AGEMA_signal_3149), .B0_t (Midori_rounds_roundReg_out[55]), .B0_f (new_AGEMA_signal_3144), .B1_t (new_AGEMA_signal_3145), .B1_f (new_AGEMA_signal_3146), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n12), .Z0_f (new_AGEMA_signal_3153), .Z1_t (new_AGEMA_signal_3154), .Z1_f (new_AGEMA_signal_3155) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n15), .A0_f (new_AGEMA_signal_3162), .A1_t (new_AGEMA_signal_3163), .A1_f (new_AGEMA_signal_3164), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n7), .B0_f (new_AGEMA_signal_4442), .B1_t (new_AGEMA_signal_4443), .B1_f (new_AGEMA_signal_4444), .Z0_t (Midori_rounds_SR_Result[6]), .Z0_f (new_AGEMA_signal_4760), .Z1_t (new_AGEMA_signal_4761), .Z1_f (new_AGEMA_signal_4762) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n6), .A0_f (new_AGEMA_signal_4020), .A1_t (new_AGEMA_signal_4021), .A1_f (new_AGEMA_signal_4022), .B0_t (Midori_rounds_roundReg_out[53]), .B0_f (new_AGEMA_signal_4011), .B1_t (new_AGEMA_signal_4012), .B1_f (new_AGEMA_signal_4013), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n7), .Z0_f (new_AGEMA_signal_4442), .Z1_t (new_AGEMA_signal_4443), .Z1_f (new_AGEMA_signal_4444) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n5), .A0_f (new_AGEMA_signal_3159), .A1_t (new_AGEMA_signal_3160), .A1_f (new_AGEMA_signal_3161), .B0_t (Midori_rounds_roundReg_out[54]), .B0_f (new_AGEMA_signal_3147), .B1_t (new_AGEMA_signal_3148), .B1_f (new_AGEMA_signal_3149), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n6), .Z0_f (new_AGEMA_signal_4020), .Z1_t (new_AGEMA_signal_4021), .Z1_f (new_AGEMA_signal_4022) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U10 ( .A0_t (Midori_rounds_roundReg_out[52]), .A0_f (new_AGEMA_signal_3156), .A1_t (new_AGEMA_signal_3157), .A1_f (new_AGEMA_signal_3158), .B0_t (Midori_rounds_roundReg_out[55]), .B0_f (new_AGEMA_signal_3144), .B1_t (new_AGEMA_signal_3145), .B1_f (new_AGEMA_signal_3146), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n5), .Z0_f (new_AGEMA_signal_3159), .Z1_t (new_AGEMA_signal_3160), .Z1_f (new_AGEMA_signal_3161) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U9 ( .A0_t (Midori_rounds_roundReg_out[55]), .A0_f (new_AGEMA_signal_3144), .A1_t (new_AGEMA_signal_3145), .A1_f (new_AGEMA_signal_3146), .B0_t (Midori_rounds_roundReg_out[52]), .B0_f (new_AGEMA_signal_3156), .B1_t (new_AGEMA_signal_3157), .B1_f (new_AGEMA_signal_3158), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n15), .Z0_f (new_AGEMA_signal_3162), .Z1_t (new_AGEMA_signal_3163), .Z1_f (new_AGEMA_signal_3164) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n13), .A0_f (new_AGEMA_signal_3168), .A1_t (new_AGEMA_signal_3169), .A1_f (new_AGEMA_signal_3170), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n3), .B0_f (new_AGEMA_signal_4445), .B1_t (new_AGEMA_signal_4446), .B1_f (new_AGEMA_signal_4447), .Z0_t (Midori_rounds_SR_Result[4]), .Z0_f (new_AGEMA_signal_4763), .Z1_t (new_AGEMA_signal_4764), .Z1_f (new_AGEMA_signal_4765) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U7 ( .A0_t (Midori_rounds_roundReg_out[53]), .A0_f (new_AGEMA_signal_4011), .A1_t (new_AGEMA_signal_4012), .A1_f (new_AGEMA_signal_4013), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n2), .B0_f (new_AGEMA_signal_4023), .B1_t (new_AGEMA_signal_4024), .B1_f (new_AGEMA_signal_4025), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n3), .Z0_f (new_AGEMA_signal_4445), .Z1_t (new_AGEMA_signal_4446), .Z1_f (new_AGEMA_signal_4447) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U6 ( .A0_t (Midori_rounds_roundReg_out[52]), .A0_f (new_AGEMA_signal_3156), .A1_t (new_AGEMA_signal_3157), .A1_f (new_AGEMA_signal_3158), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n1), .B0_f (new_AGEMA_signal_3165), .B1_t (new_AGEMA_signal_3166), .B1_f (new_AGEMA_signal_3167), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n2), .Z0_f (new_AGEMA_signal_4023), .Z1_t (new_AGEMA_signal_4024), .Z1_f (new_AGEMA_signal_4025) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U5 ( .A0_t (Midori_rounds_roundReg_out[54]), .A0_f (new_AGEMA_signal_3147), .A1_t (new_AGEMA_signal_3148), .A1_f (new_AGEMA_signal_3149), .B0_t (Midori_rounds_roundReg_out[55]), .B0_f (new_AGEMA_signal_3144), .B1_t (new_AGEMA_signal_3145), .B1_f (new_AGEMA_signal_3146), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n1), .Z0_f (new_AGEMA_signal_3165), .Z1_t (new_AGEMA_signal_3166), .Z1_f (new_AGEMA_signal_3167) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U3 ( .A0_t (Midori_rounds_roundReg_out[54]), .A0_f (new_AGEMA_signal_3147), .A1_t (new_AGEMA_signal_3148), .A1_f (new_AGEMA_signal_3149), .B0_t (Midori_rounds_roundReg_out[55]), .B0_f (new_AGEMA_signal_3144), .B1_t (new_AGEMA_signal_3145), .B1_f (new_AGEMA_signal_3146), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n13), .Z0_f (new_AGEMA_signal_3168), .Z1_t (new_AGEMA_signal_3169), .Z1_f (new_AGEMA_signal_3170) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n15), .A0_f (new_AGEMA_signal_3189), .A1_t (new_AGEMA_signal_3190), .A1_f (new_AGEMA_signal_3191), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n14), .B0_f (new_AGEMA_signal_4029), .B1_t (new_AGEMA_signal_4030), .B1_f (new_AGEMA_signal_4031), .Z0_t (Midori_rounds_SR_Result[35]), .Z0_f (new_AGEMA_signal_4448), .Z1_t (new_AGEMA_signal_4449), .Z1_f (new_AGEMA_signal_4450) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n13), .A0_f (new_AGEMA_signal_3195), .A1_t (new_AGEMA_signal_3196), .A1_f (new_AGEMA_signal_3197), .B0_t (Midori_rounds_roundReg_out[57]), .B0_f (new_AGEMA_signal_4026), .B1_t (new_AGEMA_signal_4027), .B1_f (new_AGEMA_signal_4028), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n14), .Z0_f (new_AGEMA_signal_4029), .Z1_t (new_AGEMA_signal_4030), .Z1_f (new_AGEMA_signal_4031) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n12), .A0_f (new_AGEMA_signal_3180), .A1_t (new_AGEMA_signal_3181), .A1_f (new_AGEMA_signal_3182), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n11), .B0_f (new_AGEMA_signal_4032), .B1_t (new_AGEMA_signal_4033), .B1_f (new_AGEMA_signal_4034), .Z0_t (Midori_rounds_SR_Result[33]), .Z0_f (new_AGEMA_signal_4451), .Z1_t (new_AGEMA_signal_4452), .Z1_f (new_AGEMA_signal_4453) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U16 ( .A0_t (Midori_rounds_roundReg_out[56]), .A0_f (new_AGEMA_signal_3183), .A1_t (new_AGEMA_signal_3184), .A1_f (new_AGEMA_signal_3185), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n10), .B0_f (new_AGEMA_signal_3177), .B1_t (new_AGEMA_signal_3178), .B1_f (new_AGEMA_signal_3179), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n11), .Z0_f (new_AGEMA_signal_4032), .Z1_t (new_AGEMA_signal_4033), .Z1_f (new_AGEMA_signal_4034) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U15 ( .A0_t (Midori_rounds_roundReg_out[59]), .A0_f (new_AGEMA_signal_3171), .A1_t (new_AGEMA_signal_3172), .A1_f (new_AGEMA_signal_3173), .B0_t (Midori_rounds_roundReg_out[58]), .B0_f (new_AGEMA_signal_3174), .B1_t (new_AGEMA_signal_3175), .B1_f (new_AGEMA_signal_3176), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n10), .Z0_f (new_AGEMA_signal_3177), .Z1_t (new_AGEMA_signal_3178), .Z1_f (new_AGEMA_signal_3179) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U14 ( .A0_t (Midori_rounds_roundReg_out[58]), .A0_f (new_AGEMA_signal_3174), .A1_t (new_AGEMA_signal_3175), .A1_f (new_AGEMA_signal_3176), .B0_t (Midori_rounds_roundReg_out[59]), .B0_f (new_AGEMA_signal_3171), .B1_t (new_AGEMA_signal_3172), .B1_f (new_AGEMA_signal_3173), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n12), .Z0_f (new_AGEMA_signal_3180), .Z1_t (new_AGEMA_signal_3181), .Z1_f (new_AGEMA_signal_3182) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n15), .A0_f (new_AGEMA_signal_3189), .A1_t (new_AGEMA_signal_3190), .A1_f (new_AGEMA_signal_3191), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n7), .B0_f (new_AGEMA_signal_4454), .B1_t (new_AGEMA_signal_4455), .B1_f (new_AGEMA_signal_4456), .Z0_t (Midori_rounds_SR_Result[34]), .Z0_f (new_AGEMA_signal_4766), .Z1_t (new_AGEMA_signal_4767), .Z1_f (new_AGEMA_signal_4768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n6), .A0_f (new_AGEMA_signal_4035), .A1_t (new_AGEMA_signal_4036), .A1_f (new_AGEMA_signal_4037), .B0_t (Midori_rounds_roundReg_out[57]), .B0_f (new_AGEMA_signal_4026), .B1_t (new_AGEMA_signal_4027), .B1_f (new_AGEMA_signal_4028), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n7), .Z0_f (new_AGEMA_signal_4454), .Z1_t (new_AGEMA_signal_4455), .Z1_f (new_AGEMA_signal_4456) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n5), .A0_f (new_AGEMA_signal_3186), .A1_t (new_AGEMA_signal_3187), .A1_f (new_AGEMA_signal_3188), .B0_t (Midori_rounds_roundReg_out[58]), .B0_f (new_AGEMA_signal_3174), .B1_t (new_AGEMA_signal_3175), .B1_f (new_AGEMA_signal_3176), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n6), .Z0_f (new_AGEMA_signal_4035), .Z1_t (new_AGEMA_signal_4036), .Z1_f (new_AGEMA_signal_4037) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U10 ( .A0_t (Midori_rounds_roundReg_out[56]), .A0_f (new_AGEMA_signal_3183), .A1_t (new_AGEMA_signal_3184), .A1_f (new_AGEMA_signal_3185), .B0_t (Midori_rounds_roundReg_out[59]), .B0_f (new_AGEMA_signal_3171), .B1_t (new_AGEMA_signal_3172), .B1_f (new_AGEMA_signal_3173), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n5), .Z0_f (new_AGEMA_signal_3186), .Z1_t (new_AGEMA_signal_3187), .Z1_f (new_AGEMA_signal_3188) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U9 ( .A0_t (Midori_rounds_roundReg_out[59]), .A0_f (new_AGEMA_signal_3171), .A1_t (new_AGEMA_signal_3172), .A1_f (new_AGEMA_signal_3173), .B0_t (Midori_rounds_roundReg_out[56]), .B0_f (new_AGEMA_signal_3183), .B1_t (new_AGEMA_signal_3184), .B1_f (new_AGEMA_signal_3185), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n15), .Z0_f (new_AGEMA_signal_3189), .Z1_t (new_AGEMA_signal_3190), .Z1_f (new_AGEMA_signal_3191) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n13), .A0_f (new_AGEMA_signal_3195), .A1_t (new_AGEMA_signal_3196), .A1_f (new_AGEMA_signal_3197), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n3), .B0_f (new_AGEMA_signal_4457), .B1_t (new_AGEMA_signal_4458), .B1_f (new_AGEMA_signal_4459), .Z0_t (Midori_rounds_SR_Result[32]), .Z0_f (new_AGEMA_signal_4769), .Z1_t (new_AGEMA_signal_4770), .Z1_f (new_AGEMA_signal_4771) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U7 ( .A0_t (Midori_rounds_roundReg_out[57]), .A0_f (new_AGEMA_signal_4026), .A1_t (new_AGEMA_signal_4027), .A1_f (new_AGEMA_signal_4028), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n2), .B0_f (new_AGEMA_signal_4038), .B1_t (new_AGEMA_signal_4039), .B1_f (new_AGEMA_signal_4040), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n3), .Z0_f (new_AGEMA_signal_4457), .Z1_t (new_AGEMA_signal_4458), .Z1_f (new_AGEMA_signal_4459) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U6 ( .A0_t (Midori_rounds_roundReg_out[56]), .A0_f (new_AGEMA_signal_3183), .A1_t (new_AGEMA_signal_3184), .A1_f (new_AGEMA_signal_3185), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n1), .B0_f (new_AGEMA_signal_3192), .B1_t (new_AGEMA_signal_3193), .B1_f (new_AGEMA_signal_3194), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n2), .Z0_f (new_AGEMA_signal_4038), .Z1_t (new_AGEMA_signal_4039), .Z1_f (new_AGEMA_signal_4040) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U5 ( .A0_t (Midori_rounds_roundReg_out[58]), .A0_f (new_AGEMA_signal_3174), .A1_t (new_AGEMA_signal_3175), .A1_f (new_AGEMA_signal_3176), .B0_t (Midori_rounds_roundReg_out[59]), .B0_f (new_AGEMA_signal_3171), .B1_t (new_AGEMA_signal_3172), .B1_f (new_AGEMA_signal_3173), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n1), .Z0_f (new_AGEMA_signal_3192), .Z1_t (new_AGEMA_signal_3193), .Z1_f (new_AGEMA_signal_3194) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U3 ( .A0_t (Midori_rounds_roundReg_out[58]), .A0_f (new_AGEMA_signal_3174), .A1_t (new_AGEMA_signal_3175), .A1_f (new_AGEMA_signal_3176), .B0_t (Midori_rounds_roundReg_out[59]), .B0_f (new_AGEMA_signal_3171), .B1_t (new_AGEMA_signal_3172), .B1_f (new_AGEMA_signal_3173), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n13), .Z0_f (new_AGEMA_signal_3195), .Z1_t (new_AGEMA_signal_3196), .Z1_f (new_AGEMA_signal_3197) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n15), .A0_f (new_AGEMA_signal_4460), .A1_t (new_AGEMA_signal_4461), .A1_f (new_AGEMA_signal_4462), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n14), .B0_f (new_AGEMA_signal_3213), .B1_t (new_AGEMA_signal_3214), .B1_f (new_AGEMA_signal_3215), .Z0_t (Midori_rounds_SR_Result[60]), .Z0_f (new_AGEMA_signal_4772), .Z1_t (new_AGEMA_signal_4773), .Z1_f (new_AGEMA_signal_4774) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U18 ( .A0_t (Midori_rounds_roundReg_out[61]), .A0_f (new_AGEMA_signal_4047), .A1_t (new_AGEMA_signal_4048), .A1_f (new_AGEMA_signal_4049), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n13), .B0_f (new_AGEMA_signal_4041), .B1_t (new_AGEMA_signal_4042), .B1_f (new_AGEMA_signal_4043), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n15), .Z0_f (new_AGEMA_signal_4460), .Z1_t (new_AGEMA_signal_4461), .Z1_f (new_AGEMA_signal_4462) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U17 ( .A0_t (Midori_rounds_roundReg_out[60]), .A0_f (new_AGEMA_signal_3207), .A1_t (new_AGEMA_signal_3208), .A1_f (new_AGEMA_signal_3209), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n11), .B0_f (new_AGEMA_signal_3204), .B1_t (new_AGEMA_signal_3205), .B1_f (new_AGEMA_signal_3206), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n13), .Z0_f (new_AGEMA_signal_4041), .Z1_t (new_AGEMA_signal_4042), .Z1_f (new_AGEMA_signal_4043) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U16 ( .A0_t (Midori_rounds_roundReg_out[62]), .A0_f (new_AGEMA_signal_3198), .A1_t (new_AGEMA_signal_3199), .A1_f (new_AGEMA_signal_3200), .B0_t (Midori_rounds_roundReg_out[63]), .B0_f (new_AGEMA_signal_3201), .B1_t (new_AGEMA_signal_3202), .B1_f (new_AGEMA_signal_3203), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n11), .Z0_f (new_AGEMA_signal_3204), .Z1_t (new_AGEMA_signal_3205), .Z1_f (new_AGEMA_signal_3206) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n10), .A0_f (new_AGEMA_signal_4463), .A1_t (new_AGEMA_signal_4464), .A1_f (new_AGEMA_signal_4465), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n9), .B0_f (new_AGEMA_signal_3216), .B1_t (new_AGEMA_signal_3217), .B1_f (new_AGEMA_signal_3218), .Z0_t (Midori_rounds_SR_Result[62]), .Z0_f (new_AGEMA_signal_4775), .Z1_t (new_AGEMA_signal_4776), .Z1_f (new_AGEMA_signal_4777) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n8), .A0_f (new_AGEMA_signal_4044), .A1_t (new_AGEMA_signal_4045), .A1_f (new_AGEMA_signal_4046), .B0_t (Midori_rounds_roundReg_out[61]), .B0_f (new_AGEMA_signal_4047), .B1_t (new_AGEMA_signal_4048), .B1_f (new_AGEMA_signal_4049), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n10), .Z0_f (new_AGEMA_signal_4463), .Z1_t (new_AGEMA_signal_4464), .Z1_f (new_AGEMA_signal_4465) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n7), .A0_f (new_AGEMA_signal_3210), .A1_t (new_AGEMA_signal_3211), .A1_f (new_AGEMA_signal_3212), .B0_t (Midori_rounds_roundReg_out[62]), .B0_f (new_AGEMA_signal_3198), .B1_t (new_AGEMA_signal_3199), .B1_f (new_AGEMA_signal_3200), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n8), .Z0_f (new_AGEMA_signal_4044), .Z1_t (new_AGEMA_signal_4045), .Z1_f (new_AGEMA_signal_4046) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U12 ( .A0_t (Midori_rounds_roundReg_out[60]), .A0_f (new_AGEMA_signal_3207), .A1_t (new_AGEMA_signal_3208), .A1_f (new_AGEMA_signal_3209), .B0_t (Midori_rounds_roundReg_out[63]), .B0_f (new_AGEMA_signal_3201), .B1_t (new_AGEMA_signal_3202), .B1_f (new_AGEMA_signal_3203), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n7), .Z0_f (new_AGEMA_signal_3210), .Z1_t (new_AGEMA_signal_3211), .Z1_f (new_AGEMA_signal_3212) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n9), .A0_f (new_AGEMA_signal_3216), .A1_t (new_AGEMA_signal_3217), .A1_f (new_AGEMA_signal_3218), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n5), .B0_f (new_AGEMA_signal_4050), .B1_t (new_AGEMA_signal_4051), .B1_f (new_AGEMA_signal_4052), .Z0_t (Midori_rounds_SR_Result[63]), .Z0_f (new_AGEMA_signal_4466), .Z1_t (new_AGEMA_signal_4467), .Z1_f (new_AGEMA_signal_4468) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U10 ( .A0_t (Midori_rounds_roundReg_out[61]), .A0_f (new_AGEMA_signal_4047), .A1_t (new_AGEMA_signal_4048), .A1_f (new_AGEMA_signal_4049), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n14), .B0_f (new_AGEMA_signal_3213), .B1_t (new_AGEMA_signal_3214), .B1_f (new_AGEMA_signal_3215), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n5), .Z0_f (new_AGEMA_signal_4050), .Z1_t (new_AGEMA_signal_4051), .Z1_f (new_AGEMA_signal_4052) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U9 ( .A0_t (Midori_rounds_roundReg_out[62]), .A0_f (new_AGEMA_signal_3198), .A1_t (new_AGEMA_signal_3199), .A1_f (new_AGEMA_signal_3200), .B0_t (Midori_rounds_roundReg_out[63]), .B0_f (new_AGEMA_signal_3201), .B1_t (new_AGEMA_signal_3202), .B1_f (new_AGEMA_signal_3203), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n14), .Z0_f (new_AGEMA_signal_3213), .Z1_t (new_AGEMA_signal_3214), .Z1_f (new_AGEMA_signal_3215) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U8 ( .A0_t (Midori_rounds_roundReg_out[63]), .A0_f (new_AGEMA_signal_3201), .A1_t (new_AGEMA_signal_3202), .A1_f (new_AGEMA_signal_3203), .B0_t (Midori_rounds_roundReg_out[60]), .B0_f (new_AGEMA_signal_3207), .B1_t (new_AGEMA_signal_3208), .B1_f (new_AGEMA_signal_3209), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n9), .Z0_f (new_AGEMA_signal_3216), .Z1_t (new_AGEMA_signal_3217), .Z1_f (new_AGEMA_signal_3218) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n3), .A0_f (new_AGEMA_signal_3222), .A1_t (new_AGEMA_signal_3223), .A1_f (new_AGEMA_signal_3224), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n2), .B0_f (new_AGEMA_signal_4053), .B1_t (new_AGEMA_signal_4054), .B1_f (new_AGEMA_signal_4055), .Z0_t (Midori_rounds_SR_Result[61]), .Z0_f (new_AGEMA_signal_4469), .Z1_t (new_AGEMA_signal_4470), .Z1_f (new_AGEMA_signal_4471) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n1), .A0_f (new_AGEMA_signal_3219), .A1_t (new_AGEMA_signal_3220), .A1_f (new_AGEMA_signal_3221), .B0_t (Midori_rounds_roundReg_out[63]), .B0_f (new_AGEMA_signal_3201), .B1_t (new_AGEMA_signal_3202), .B1_f (new_AGEMA_signal_3203), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n2), .Z0_f (new_AGEMA_signal_4053), .Z1_t (new_AGEMA_signal_4054), .Z1_f (new_AGEMA_signal_4055) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U4 ( .A0_t (Midori_rounds_roundReg_out[62]), .A0_f (new_AGEMA_signal_3198), .A1_t (new_AGEMA_signal_3199), .A1_f (new_AGEMA_signal_3200), .B0_t (Midori_rounds_roundReg_out[60]), .B0_f (new_AGEMA_signal_3207), .B1_t (new_AGEMA_signal_3208), .B1_f (new_AGEMA_signal_3209), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n1), .Z0_f (new_AGEMA_signal_3219), .Z1_t (new_AGEMA_signal_3220), .Z1_f (new_AGEMA_signal_3221) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U1 ( .A0_t (Midori_rounds_roundReg_out[62]), .A0_f (new_AGEMA_signal_3198), .A1_t (new_AGEMA_signal_3199), .A1_f (new_AGEMA_signal_3200), .B0_t (Midori_rounds_roundReg_out[60]), .B0_f (new_AGEMA_signal_3207), .B1_t (new_AGEMA_signal_3208), .B1_f (new_AGEMA_signal_3209), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n3), .Z0_f (new_AGEMA_signal_3222), .Z1_t (new_AGEMA_signal_3223), .Z1_f (new_AGEMA_signal_3224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_0_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[0]), .A0_f (new_AGEMA_signal_4727), .A1_t (new_AGEMA_signal_4728), .A1_f (new_AGEMA_signal_4729), .B0_t (Midori_rounds_sub_ResultXORkey[0]), .B0_f (new_AGEMA_signal_5809), .B1_t (new_AGEMA_signal_5810), .B1_f (new_AGEMA_signal_5811), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_5990), .Z1_t (new_AGEMA_signal_5991), .Z1_f (new_AGEMA_signal_5992) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_5990), .B1_t (new_AGEMA_signal_5991), .B1_f (new_AGEMA_signal_5992), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_6170), .Z1_t (new_AGEMA_signal_6171), .Z1_f (new_AGEMA_signal_6172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_0_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_6170), .A1_t (new_AGEMA_signal_6171), .A1_f (new_AGEMA_signal_6172), .B0_t (Midori_rounds_SR_Result[0]), .B0_f (new_AGEMA_signal_4727), .B1_t (new_AGEMA_signal_4728), .B1_f (new_AGEMA_signal_4729), .Z0_t (Midori_rounds_mul_input[0]), .Z0_f (new_AGEMA_signal_6449), .Z1_t (new_AGEMA_signal_6450), .Z1_f (new_AGEMA_signal_6451) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_1_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[1]), .A0_f (new_AGEMA_signal_4367), .A1_t (new_AGEMA_signal_4368), .A1_f (new_AGEMA_signal_4369), .B0_t (Midori_rounds_sub_ResultXORkey[1]), .B0_f (new_AGEMA_signal_4615), .B1_t (new_AGEMA_signal_4616), .B1_f (new_AGEMA_signal_4617), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_4936), .Z1_t (new_AGEMA_signal_4937), .Z1_f (new_AGEMA_signal_4938) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_4936), .B1_t (new_AGEMA_signal_4937), .B1_f (new_AGEMA_signal_4938), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_5044), .Z1_t (new_AGEMA_signal_5045), .Z1_f (new_AGEMA_signal_5046) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_1_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_5044), .A1_t (new_AGEMA_signal_5045), .A1_f (new_AGEMA_signal_5046), .B0_t (Midori_rounds_SR_Result[1]), .B0_f (new_AGEMA_signal_4367), .B1_t (new_AGEMA_signal_4368), .B1_f (new_AGEMA_signal_4369), .Z0_t (Midori_rounds_mul_input[1]), .Z0_f (new_AGEMA_signal_5201), .Z1_t (new_AGEMA_signal_5202), .Z1_f (new_AGEMA_signal_5203) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_2_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[2]), .A0_f (new_AGEMA_signal_4724), .A1_t (new_AGEMA_signal_4725), .A1_f (new_AGEMA_signal_4726), .B0_t (Midori_rounds_sub_ResultXORkey[2]), .B0_f (new_AGEMA_signal_4893), .B1_t (new_AGEMA_signal_4894), .B1_f (new_AGEMA_signal_4895), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_5047), .Z1_t (new_AGEMA_signal_5048), .Z1_f (new_AGEMA_signal_5049) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_5047), .B1_t (new_AGEMA_signal_5048), .B1_f (new_AGEMA_signal_5049), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_5204), .Z1_t (new_AGEMA_signal_5205), .Z1_f (new_AGEMA_signal_5206) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_2_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_5204), .A1_t (new_AGEMA_signal_5205), .A1_f (new_AGEMA_signal_5206), .B0_t (Midori_rounds_SR_Result[2]), .B0_f (new_AGEMA_signal_4724), .B1_t (new_AGEMA_signal_4725), .B1_f (new_AGEMA_signal_4726), .Z0_t (Midori_rounds_mul_input[2]), .Z0_f (new_AGEMA_signal_5362), .Z1_t (new_AGEMA_signal_5363), .Z1_f (new_AGEMA_signal_5364) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_3_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[3]), .A0_f (new_AGEMA_signal_4364), .A1_t (new_AGEMA_signal_4365), .A1_f (new_AGEMA_signal_4366), .B0_t (Midori_rounds_sub_ResultXORkey[3]), .B0_f (new_AGEMA_signal_4612), .B1_t (new_AGEMA_signal_4613), .B1_f (new_AGEMA_signal_4614), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_4939), .Z1_t (new_AGEMA_signal_4940), .Z1_f (new_AGEMA_signal_4941) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_4939), .B1_t (new_AGEMA_signal_4940), .B1_f (new_AGEMA_signal_4941), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_5050), .Z1_t (new_AGEMA_signal_5051), .Z1_f (new_AGEMA_signal_5052) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_3_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_5050), .A1_t (new_AGEMA_signal_5051), .A1_f (new_AGEMA_signal_5052), .B0_t (Midori_rounds_SR_Result[3]), .B0_f (new_AGEMA_signal_4364), .B1_t (new_AGEMA_signal_4365), .B1_f (new_AGEMA_signal_4366), .Z0_t (Midori_rounds_mul_input[3]), .Z0_f (new_AGEMA_signal_5207), .Z1_t (new_AGEMA_signal_5208), .Z1_f (new_AGEMA_signal_5209) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_4_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[4]), .A0_f (new_AGEMA_signal_4763), .A1_t (new_AGEMA_signal_4764), .A1_f (new_AGEMA_signal_4765), .B0_t (Midori_rounds_sub_ResultXORkey[4]), .B0_f (new_AGEMA_signal_6167), .B1_t (new_AGEMA_signal_6168), .B1_f (new_AGEMA_signal_6169), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_4_U1_X), .Z0_f (new_AGEMA_signal_6452), .Z1_t (new_AGEMA_signal_6453), .Z1_f (new_AGEMA_signal_6454) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_4_U1_X), .B0_f (new_AGEMA_signal_6452), .B1_t (new_AGEMA_signal_6453), .B1_f (new_AGEMA_signal_6454), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_4_U1_Y), .Z0_f (new_AGEMA_signal_6677), .Z1_t (new_AGEMA_signal_6678), .Z1_f (new_AGEMA_signal_6679) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_4_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_4_U1_Y), .A0_f (new_AGEMA_signal_6677), .A1_t (new_AGEMA_signal_6678), .A1_f (new_AGEMA_signal_6679), .B0_t (Midori_rounds_SR_Result[4]), .B0_f (new_AGEMA_signal_4763), .B1_t (new_AGEMA_signal_4764), .B1_f (new_AGEMA_signal_4765), .Z0_t (Midori_rounds_mul_input[4]), .Z0_f (new_AGEMA_signal_6755), .Z1_t (new_AGEMA_signal_6756), .Z1_f (new_AGEMA_signal_6757) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_5_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[5]), .A0_f (new_AGEMA_signal_4439), .A1_t (new_AGEMA_signal_4440), .A1_f (new_AGEMA_signal_4441), .B0_t (Midori_rounds_sub_ResultXORkey[5]), .B0_f (new_AGEMA_signal_4609), .B1_t (new_AGEMA_signal_4610), .B1_f (new_AGEMA_signal_4611), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_5_U1_X), .Z0_f (new_AGEMA_signal_4942), .Z1_t (new_AGEMA_signal_4943), .Z1_f (new_AGEMA_signal_4944) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_5_U1_X), .B0_f (new_AGEMA_signal_4942), .B1_t (new_AGEMA_signal_4943), .B1_f (new_AGEMA_signal_4944), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_5_U1_Y), .Z0_f (new_AGEMA_signal_5053), .Z1_t (new_AGEMA_signal_5054), .Z1_f (new_AGEMA_signal_5055) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_5_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_5_U1_Y), .A0_f (new_AGEMA_signal_5053), .A1_t (new_AGEMA_signal_5054), .A1_f (new_AGEMA_signal_5055), .B0_t (Midori_rounds_SR_Result[5]), .B0_f (new_AGEMA_signal_4439), .B1_t (new_AGEMA_signal_4440), .B1_f (new_AGEMA_signal_4441), .Z0_t (Midori_rounds_mul_input[5]), .Z0_f (new_AGEMA_signal_5210), .Z1_t (new_AGEMA_signal_5211), .Z1_f (new_AGEMA_signal_5212) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_6_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[6]), .A0_f (new_AGEMA_signal_4760), .A1_t (new_AGEMA_signal_4761), .A1_f (new_AGEMA_signal_4762), .B0_t (Midori_rounds_sub_ResultXORkey[6]), .B0_f (new_AGEMA_signal_4896), .B1_t (new_AGEMA_signal_4897), .B1_f (new_AGEMA_signal_4898), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_6_U1_X), .Z0_f (new_AGEMA_signal_5056), .Z1_t (new_AGEMA_signal_5057), .Z1_f (new_AGEMA_signal_5058) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_6_U1_X), .B0_f (new_AGEMA_signal_5056), .B1_t (new_AGEMA_signal_5057), .B1_f (new_AGEMA_signal_5058), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_6_U1_Y), .Z0_f (new_AGEMA_signal_5213), .Z1_t (new_AGEMA_signal_5214), .Z1_f (new_AGEMA_signal_5215) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_6_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_6_U1_Y), .A0_f (new_AGEMA_signal_5213), .A1_t (new_AGEMA_signal_5214), .A1_f (new_AGEMA_signal_5215), .B0_t (Midori_rounds_SR_Result[6]), .B0_f (new_AGEMA_signal_4760), .B1_t (new_AGEMA_signal_4761), .B1_f (new_AGEMA_signal_4762), .Z0_t (Midori_rounds_mul_input[6]), .Z0_f (new_AGEMA_signal_5365), .Z1_t (new_AGEMA_signal_5366), .Z1_f (new_AGEMA_signal_5367) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_7_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[7]), .A0_f (new_AGEMA_signal_4436), .A1_t (new_AGEMA_signal_4437), .A1_f (new_AGEMA_signal_4438), .B0_t (Midori_rounds_sub_ResultXORkey[7]), .B0_f (new_AGEMA_signal_4606), .B1_t (new_AGEMA_signal_4607), .B1_f (new_AGEMA_signal_4608), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_7_U1_X), .Z0_f (new_AGEMA_signal_4945), .Z1_t (new_AGEMA_signal_4946), .Z1_f (new_AGEMA_signal_4947) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_7_U1_X), .B0_f (new_AGEMA_signal_4945), .B1_t (new_AGEMA_signal_4946), .B1_f (new_AGEMA_signal_4947), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_7_U1_Y), .Z0_f (new_AGEMA_signal_5059), .Z1_t (new_AGEMA_signal_5060), .Z1_f (new_AGEMA_signal_5061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_7_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_7_U1_Y), .A0_f (new_AGEMA_signal_5059), .A1_t (new_AGEMA_signal_5060), .A1_f (new_AGEMA_signal_5061), .B0_t (Midori_rounds_SR_Result[7]), .B0_f (new_AGEMA_signal_4436), .B1_t (new_AGEMA_signal_4437), .B1_f (new_AGEMA_signal_4438), .Z0_t (Midori_rounds_mul_input[7]), .Z0_f (new_AGEMA_signal_5216), .Z1_t (new_AGEMA_signal_5217), .Z1_f (new_AGEMA_signal_5218) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_8_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[8]), .A0_f (new_AGEMA_signal_4694), .A1_t (new_AGEMA_signal_4695), .A1_f (new_AGEMA_signal_4696), .B0_t (Midori_rounds_sub_ResultXORkey[8]), .B0_f (new_AGEMA_signal_5806), .B1_t (new_AGEMA_signal_5807), .B1_f (new_AGEMA_signal_5808), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_8_U1_X), .Z0_f (new_AGEMA_signal_5993), .Z1_t (new_AGEMA_signal_5994), .Z1_f (new_AGEMA_signal_5995) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_8_U1_X), .B0_f (new_AGEMA_signal_5993), .B1_t (new_AGEMA_signal_5994), .B1_f (new_AGEMA_signal_5995), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_8_U1_Y), .Z0_f (new_AGEMA_signal_6173), .Z1_t (new_AGEMA_signal_6174), .Z1_f (new_AGEMA_signal_6175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_8_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_8_U1_Y), .A0_f (new_AGEMA_signal_6173), .A1_t (new_AGEMA_signal_6174), .A1_f (new_AGEMA_signal_6175), .B0_t (Midori_rounds_SR_Result[8]), .B0_f (new_AGEMA_signal_4694), .B1_t (new_AGEMA_signal_4695), .B1_f (new_AGEMA_signal_4696), .Z0_t (Midori_rounds_mul_input[8]), .Z0_f (new_AGEMA_signal_6455), .Z1_t (new_AGEMA_signal_6456), .Z1_f (new_AGEMA_signal_6457) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_9_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[9]), .A0_f (new_AGEMA_signal_4313), .A1_t (new_AGEMA_signal_4314), .A1_f (new_AGEMA_signal_4315), .B0_t (Midori_rounds_sub_ResultXORkey[9]), .B0_f (new_AGEMA_signal_4657), .B1_t (new_AGEMA_signal_4658), .B1_f (new_AGEMA_signal_4659), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_9_U1_X), .Z0_f (new_AGEMA_signal_4948), .Z1_t (new_AGEMA_signal_4949), .Z1_f (new_AGEMA_signal_4950) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_9_U1_X), .B0_f (new_AGEMA_signal_4948), .B1_t (new_AGEMA_signal_4949), .B1_f (new_AGEMA_signal_4950), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_9_U1_Y), .Z0_f (new_AGEMA_signal_5062), .Z1_t (new_AGEMA_signal_5063), .Z1_f (new_AGEMA_signal_5064) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_9_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_9_U1_Y), .A0_f (new_AGEMA_signal_5062), .A1_t (new_AGEMA_signal_5063), .A1_f (new_AGEMA_signal_5064), .B0_t (Midori_rounds_SR_Result[9]), .B0_f (new_AGEMA_signal_4313), .B1_t (new_AGEMA_signal_4314), .B1_f (new_AGEMA_signal_4315), .Z0_t (Midori_rounds_mul_input[9]), .Z0_f (new_AGEMA_signal_5219), .Z1_t (new_AGEMA_signal_5220), .Z1_f (new_AGEMA_signal_5221) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_10_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[10]), .A0_f (new_AGEMA_signal_4697), .A1_t (new_AGEMA_signal_4698), .A1_f (new_AGEMA_signal_4699), .B0_t (Midori_rounds_sub_ResultXORkey[10]), .B0_f (new_AGEMA_signal_4917), .B1_t (new_AGEMA_signal_4918), .B1_f (new_AGEMA_signal_4919), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_10_U1_X), .Z0_f (new_AGEMA_signal_5065), .Z1_t (new_AGEMA_signal_5066), .Z1_f (new_AGEMA_signal_5067) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_10_U1_X), .B0_f (new_AGEMA_signal_5065), .B1_t (new_AGEMA_signal_5066), .B1_f (new_AGEMA_signal_5067), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_10_U1_Y), .Z0_f (new_AGEMA_signal_5222), .Z1_t (new_AGEMA_signal_5223), .Z1_f (new_AGEMA_signal_5224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_10_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_10_U1_Y), .A0_f (new_AGEMA_signal_5222), .A1_t (new_AGEMA_signal_5223), .A1_f (new_AGEMA_signal_5224), .B0_t (Midori_rounds_SR_Result[10]), .B0_f (new_AGEMA_signal_4697), .B1_t (new_AGEMA_signal_4698), .B1_f (new_AGEMA_signal_4699), .Z0_t (Midori_rounds_mul_input[10]), .Z0_f (new_AGEMA_signal_5368), .Z1_t (new_AGEMA_signal_5369), .Z1_f (new_AGEMA_signal_5370) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_11_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[11]), .A0_f (new_AGEMA_signal_4310), .A1_t (new_AGEMA_signal_4311), .A1_f (new_AGEMA_signal_4312), .B0_t (Midori_rounds_sub_ResultXORkey[11]), .B0_f (new_AGEMA_signal_4654), .B1_t (new_AGEMA_signal_4655), .B1_f (new_AGEMA_signal_4656), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_11_U1_X), .Z0_f (new_AGEMA_signal_4951), .Z1_t (new_AGEMA_signal_4952), .Z1_f (new_AGEMA_signal_4953) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_11_U1_X), .B0_f (new_AGEMA_signal_4951), .B1_t (new_AGEMA_signal_4952), .B1_f (new_AGEMA_signal_4953), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_11_U1_Y), .Z0_f (new_AGEMA_signal_5068), .Z1_t (new_AGEMA_signal_5069), .Z1_f (new_AGEMA_signal_5070) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_11_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_11_U1_Y), .A0_f (new_AGEMA_signal_5068), .A1_t (new_AGEMA_signal_5069), .A1_f (new_AGEMA_signal_5070), .B0_t (Midori_rounds_SR_Result[11]), .B0_f (new_AGEMA_signal_4310), .B1_t (new_AGEMA_signal_4311), .B1_f (new_AGEMA_signal_4312), .Z0_t (Midori_rounds_mul_input[11]), .Z0_f (new_AGEMA_signal_5225), .Z1_t (new_AGEMA_signal_5226), .Z1_f (new_AGEMA_signal_5227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_12_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[12]), .A0_f (new_AGEMA_signal_4733), .A1_t (new_AGEMA_signal_4734), .A1_f (new_AGEMA_signal_4735), .B0_t (Midori_rounds_sub_ResultXORkey[12]), .B0_f (new_AGEMA_signal_5791), .B1_t (new_AGEMA_signal_5792), .B1_f (new_AGEMA_signal_5793), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_12_U1_X), .Z0_f (new_AGEMA_signal_5996), .Z1_t (new_AGEMA_signal_5997), .Z1_f (new_AGEMA_signal_5998) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_12_U1_X), .B0_f (new_AGEMA_signal_5996), .B1_t (new_AGEMA_signal_5997), .B1_f (new_AGEMA_signal_5998), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_12_U1_Y), .Z0_f (new_AGEMA_signal_6176), .Z1_t (new_AGEMA_signal_6177), .Z1_f (new_AGEMA_signal_6178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_12_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_12_U1_Y), .A0_f (new_AGEMA_signal_6176), .A1_t (new_AGEMA_signal_6177), .A1_f (new_AGEMA_signal_6178), .B0_t (Midori_rounds_SR_Result[12]), .B0_f (new_AGEMA_signal_4733), .B1_t (new_AGEMA_signal_4734), .B1_f (new_AGEMA_signal_4735), .Z0_t (Midori_rounds_mul_input[12]), .Z0_f (new_AGEMA_signal_6458), .Z1_t (new_AGEMA_signal_6459), .Z1_f (new_AGEMA_signal_6460) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_13_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[13]), .A0_f (new_AGEMA_signal_4379), .A1_t (new_AGEMA_signal_4380), .A1_f (new_AGEMA_signal_4381), .B0_t (Midori_rounds_sub_ResultXORkey[13]), .B0_f (new_AGEMA_signal_4663), .B1_t (new_AGEMA_signal_4664), .B1_f (new_AGEMA_signal_4665), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_13_U1_X), .Z0_f (new_AGEMA_signal_4954), .Z1_t (new_AGEMA_signal_4955), .Z1_f (new_AGEMA_signal_4956) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_13_U1_X), .B0_f (new_AGEMA_signal_4954), .B1_t (new_AGEMA_signal_4955), .B1_f (new_AGEMA_signal_4956), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_13_U1_Y), .Z0_f (new_AGEMA_signal_5071), .Z1_t (new_AGEMA_signal_5072), .Z1_f (new_AGEMA_signal_5073) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_13_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_13_U1_Y), .A0_f (new_AGEMA_signal_5071), .A1_t (new_AGEMA_signal_5072), .A1_f (new_AGEMA_signal_5073), .B0_t (Midori_rounds_SR_Result[13]), .B0_f (new_AGEMA_signal_4379), .B1_t (new_AGEMA_signal_4380), .B1_f (new_AGEMA_signal_4381), .Z0_t (Midori_rounds_mul_input[13]), .Z0_f (new_AGEMA_signal_5228), .Z1_t (new_AGEMA_signal_5229), .Z1_f (new_AGEMA_signal_5230) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_14_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[14]), .A0_f (new_AGEMA_signal_4730), .A1_t (new_AGEMA_signal_4731), .A1_f (new_AGEMA_signal_4732), .B0_t (Midori_rounds_sub_ResultXORkey[14]), .B0_f (new_AGEMA_signal_4920), .B1_t (new_AGEMA_signal_4921), .B1_f (new_AGEMA_signal_4922), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_14_U1_X), .Z0_f (new_AGEMA_signal_5074), .Z1_t (new_AGEMA_signal_5075), .Z1_f (new_AGEMA_signal_5076) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_14_U1_X), .B0_f (new_AGEMA_signal_5074), .B1_t (new_AGEMA_signal_5075), .B1_f (new_AGEMA_signal_5076), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_14_U1_Y), .Z0_f (new_AGEMA_signal_5231), .Z1_t (new_AGEMA_signal_5232), .Z1_f (new_AGEMA_signal_5233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_14_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_14_U1_Y), .A0_f (new_AGEMA_signal_5231), .A1_t (new_AGEMA_signal_5232), .A1_f (new_AGEMA_signal_5233), .B0_t (Midori_rounds_SR_Result[14]), .B0_f (new_AGEMA_signal_4730), .B1_t (new_AGEMA_signal_4731), .B1_f (new_AGEMA_signal_4732), .Z0_t (Midori_rounds_mul_input[14]), .Z0_f (new_AGEMA_signal_5371), .Z1_t (new_AGEMA_signal_5372), .Z1_f (new_AGEMA_signal_5373) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_15_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[15]), .A0_f (new_AGEMA_signal_4376), .A1_t (new_AGEMA_signal_4377), .A1_f (new_AGEMA_signal_4378), .B0_t (Midori_rounds_sub_ResultXORkey[15]), .B0_f (new_AGEMA_signal_4660), .B1_t (new_AGEMA_signal_4661), .B1_f (new_AGEMA_signal_4662), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_15_U1_X), .Z0_f (new_AGEMA_signal_4957), .Z1_t (new_AGEMA_signal_4958), .Z1_f (new_AGEMA_signal_4959) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_15_U1_X), .B0_f (new_AGEMA_signal_4957), .B1_t (new_AGEMA_signal_4958), .B1_f (new_AGEMA_signal_4959), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_15_U1_Y), .Z0_f (new_AGEMA_signal_5077), .Z1_t (new_AGEMA_signal_5078), .Z1_f (new_AGEMA_signal_5079) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_15_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_15_U1_Y), .A0_f (new_AGEMA_signal_5077), .A1_t (new_AGEMA_signal_5078), .A1_f (new_AGEMA_signal_5079), .B0_t (Midori_rounds_SR_Result[15]), .B0_f (new_AGEMA_signal_4376), .B1_t (new_AGEMA_signal_4377), .B1_f (new_AGEMA_signal_4378), .Z0_t (Midori_rounds_mul_input[15]), .Z0_f (new_AGEMA_signal_5234), .Z1_t (new_AGEMA_signal_5235), .Z1_f (new_AGEMA_signal_5236) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_16_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[16]), .A0_f (new_AGEMA_signal_4739), .A1_t (new_AGEMA_signal_4740), .A1_f (new_AGEMA_signal_4741), .B0_t (Midori_rounds_sub_ResultXORkey[16]), .B0_f (new_AGEMA_signal_5987), .B1_t (new_AGEMA_signal_5988), .B1_f (new_AGEMA_signal_5989), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_16_U1_X), .Z0_f (new_AGEMA_signal_6179), .Z1_t (new_AGEMA_signal_6180), .Z1_f (new_AGEMA_signal_6181) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_16_U1_X), .B0_f (new_AGEMA_signal_6179), .B1_t (new_AGEMA_signal_6180), .B1_f (new_AGEMA_signal_6181), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_16_U1_Y), .Z0_f (new_AGEMA_signal_6461), .Z1_t (new_AGEMA_signal_6462), .Z1_f (new_AGEMA_signal_6463) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_16_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_16_U1_Y), .A0_f (new_AGEMA_signal_6461), .A1_t (new_AGEMA_signal_6462), .A1_f (new_AGEMA_signal_6463), .B0_t (Midori_rounds_SR_Result[16]), .B0_f (new_AGEMA_signal_4739), .B1_t (new_AGEMA_signal_4740), .B1_f (new_AGEMA_signal_4741), .Z0_t (Midori_rounds_mul_input[16]), .Z0_f (new_AGEMA_signal_6680), .Z1_t (new_AGEMA_signal_6681), .Z1_f (new_AGEMA_signal_6682) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_17_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[17]), .A0_f (new_AGEMA_signal_4391), .A1_t (new_AGEMA_signal_4392), .A1_f (new_AGEMA_signal_4393), .B0_t (Midori_rounds_sub_ResultXORkey[17]), .B0_f (new_AGEMA_signal_4585), .B1_t (new_AGEMA_signal_4586), .B1_f (new_AGEMA_signal_4587), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_17_U1_X), .Z0_f (new_AGEMA_signal_4960), .Z1_t (new_AGEMA_signal_4961), .Z1_f (new_AGEMA_signal_4962) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_17_U1_X), .B0_f (new_AGEMA_signal_4960), .B1_t (new_AGEMA_signal_4961), .B1_f (new_AGEMA_signal_4962), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_17_U1_Y), .Z0_f (new_AGEMA_signal_5080), .Z1_t (new_AGEMA_signal_5081), .Z1_f (new_AGEMA_signal_5082) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_17_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_17_U1_Y), .A0_f (new_AGEMA_signal_5080), .A1_t (new_AGEMA_signal_5081), .A1_f (new_AGEMA_signal_5082), .B0_t (Midori_rounds_SR_Result[17]), .B0_f (new_AGEMA_signal_4391), .B1_t (new_AGEMA_signal_4392), .B1_f (new_AGEMA_signal_4393), .Z0_t (Midori_rounds_mul_input[17]), .Z0_f (new_AGEMA_signal_5237), .Z1_t (new_AGEMA_signal_5238), .Z1_f (new_AGEMA_signal_5239) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_18_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[18]), .A0_f (new_AGEMA_signal_4736), .A1_t (new_AGEMA_signal_4737), .A1_f (new_AGEMA_signal_4738), .B0_t (Midori_rounds_sub_ResultXORkey[18]), .B0_f (new_AGEMA_signal_4881), .B1_t (new_AGEMA_signal_4882), .B1_f (new_AGEMA_signal_4883), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_18_U1_X), .Z0_f (new_AGEMA_signal_5083), .Z1_t (new_AGEMA_signal_5084), .Z1_f (new_AGEMA_signal_5085) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_18_U1_X), .B0_f (new_AGEMA_signal_5083), .B1_t (new_AGEMA_signal_5084), .B1_f (new_AGEMA_signal_5085), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_18_U1_Y), .Z0_f (new_AGEMA_signal_5240), .Z1_t (new_AGEMA_signal_5241), .Z1_f (new_AGEMA_signal_5242) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_18_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_18_U1_Y), .A0_f (new_AGEMA_signal_5240), .A1_t (new_AGEMA_signal_5241), .A1_f (new_AGEMA_signal_5242), .B0_t (Midori_rounds_SR_Result[18]), .B0_f (new_AGEMA_signal_4736), .B1_t (new_AGEMA_signal_4737), .B1_f (new_AGEMA_signal_4738), .Z0_t (Midori_rounds_mul_input[18]), .Z0_f (new_AGEMA_signal_5374), .Z1_t (new_AGEMA_signal_5375), .Z1_f (new_AGEMA_signal_5376) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_19_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[19]), .A0_f (new_AGEMA_signal_4388), .A1_t (new_AGEMA_signal_4389), .A1_f (new_AGEMA_signal_4390), .B0_t (Midori_rounds_sub_ResultXORkey[19]), .B0_f (new_AGEMA_signal_4582), .B1_t (new_AGEMA_signal_4583), .B1_f (new_AGEMA_signal_4584), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_19_U1_X), .Z0_f (new_AGEMA_signal_4963), .Z1_t (new_AGEMA_signal_4964), .Z1_f (new_AGEMA_signal_4965) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_19_U1_X), .B0_f (new_AGEMA_signal_4963), .B1_t (new_AGEMA_signal_4964), .B1_f (new_AGEMA_signal_4965), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_19_U1_Y), .Z0_f (new_AGEMA_signal_5086), .Z1_t (new_AGEMA_signal_5087), .Z1_f (new_AGEMA_signal_5088) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_19_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_19_U1_Y), .A0_f (new_AGEMA_signal_5086), .A1_t (new_AGEMA_signal_5087), .A1_f (new_AGEMA_signal_5088), .B0_t (Midori_rounds_SR_Result[19]), .B0_f (new_AGEMA_signal_4388), .B1_t (new_AGEMA_signal_4389), .B1_f (new_AGEMA_signal_4390), .Z0_t (Midori_rounds_mul_input[19]), .Z0_f (new_AGEMA_signal_5243), .Z1_t (new_AGEMA_signal_5244), .Z1_f (new_AGEMA_signal_5245) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_20_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[20]), .A0_f (new_AGEMA_signal_4700), .A1_t (new_AGEMA_signal_4701), .A1_f (new_AGEMA_signal_4702), .B0_t (Midori_rounds_sub_ResultXORkey[20]), .B0_f (new_AGEMA_signal_5631), .B1_t (new_AGEMA_signal_5632), .B1_f (new_AGEMA_signal_5633), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_20_U1_X), .Z0_f (new_AGEMA_signal_5864), .Z1_t (new_AGEMA_signal_5865), .Z1_f (new_AGEMA_signal_5866) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_20_U1_X), .B0_f (new_AGEMA_signal_5864), .B1_t (new_AGEMA_signal_5865), .B1_f (new_AGEMA_signal_5866), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_20_U1_Y), .Z0_f (new_AGEMA_signal_5999), .Z1_t (new_AGEMA_signal_6000), .Z1_f (new_AGEMA_signal_6001) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_20_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_20_U1_Y), .A0_f (new_AGEMA_signal_5999), .A1_t (new_AGEMA_signal_6000), .A1_f (new_AGEMA_signal_6001), .B0_t (Midori_rounds_SR_Result[20]), .B0_f (new_AGEMA_signal_4700), .B1_t (new_AGEMA_signal_4701), .B1_f (new_AGEMA_signal_4702), .Z0_t (Midori_rounds_mul_input[20]), .Z0_f (new_AGEMA_signal_6182), .Z1_t (new_AGEMA_signal_6183), .Z1_f (new_AGEMA_signal_6184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_21_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[21]), .A0_f (new_AGEMA_signal_4325), .A1_t (new_AGEMA_signal_4326), .A1_f (new_AGEMA_signal_4327), .B0_t (Midori_rounds_sub_ResultXORkey[21]), .B0_f (new_AGEMA_signal_4603), .B1_t (new_AGEMA_signal_4604), .B1_f (new_AGEMA_signal_4605), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_21_U1_X), .Z0_f (new_AGEMA_signal_4966), .Z1_t (new_AGEMA_signal_4967), .Z1_f (new_AGEMA_signal_4968) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_21_U1_X), .B0_f (new_AGEMA_signal_4966), .B1_t (new_AGEMA_signal_4967), .B1_f (new_AGEMA_signal_4968), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_21_U1_Y), .Z0_f (new_AGEMA_signal_5089), .Z1_t (new_AGEMA_signal_5090), .Z1_f (new_AGEMA_signal_5091) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_21_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_21_U1_Y), .A0_f (new_AGEMA_signal_5089), .A1_t (new_AGEMA_signal_5090), .A1_f (new_AGEMA_signal_5091), .B0_t (Midori_rounds_SR_Result[21]), .B0_f (new_AGEMA_signal_4325), .B1_t (new_AGEMA_signal_4326), .B1_f (new_AGEMA_signal_4327), .Z0_t (Midori_rounds_mul_input[21]), .Z0_f (new_AGEMA_signal_5246), .Z1_t (new_AGEMA_signal_5247), .Z1_f (new_AGEMA_signal_5248) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_22_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[22]), .A0_f (new_AGEMA_signal_4703), .A1_t (new_AGEMA_signal_4704), .A1_f (new_AGEMA_signal_4705), .B0_t (Midori_rounds_sub_ResultXORkey[22]), .B0_f (new_AGEMA_signal_4890), .B1_t (new_AGEMA_signal_4891), .B1_f (new_AGEMA_signal_4892), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_22_U1_X), .Z0_f (new_AGEMA_signal_5092), .Z1_t (new_AGEMA_signal_5093), .Z1_f (new_AGEMA_signal_5094) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_22_U1_X), .B0_f (new_AGEMA_signal_5092), .B1_t (new_AGEMA_signal_5093), .B1_f (new_AGEMA_signal_5094), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_22_U1_Y), .Z0_f (new_AGEMA_signal_5249), .Z1_t (new_AGEMA_signal_5250), .Z1_f (new_AGEMA_signal_5251) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_22_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_22_U1_Y), .A0_f (new_AGEMA_signal_5249), .A1_t (new_AGEMA_signal_5250), .A1_f (new_AGEMA_signal_5251), .B0_t (Midori_rounds_SR_Result[22]), .B0_f (new_AGEMA_signal_4703), .B1_t (new_AGEMA_signal_4704), .B1_f (new_AGEMA_signal_4705), .Z0_t (Midori_rounds_mul_input[22]), .Z0_f (new_AGEMA_signal_5377), .Z1_t (new_AGEMA_signal_5378), .Z1_f (new_AGEMA_signal_5379) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_23_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[23]), .A0_f (new_AGEMA_signal_4322), .A1_t (new_AGEMA_signal_4323), .A1_f (new_AGEMA_signal_4324), .B0_t (Midori_rounds_sub_ResultXORkey[23]), .B0_f (new_AGEMA_signal_4600), .B1_t (new_AGEMA_signal_4601), .B1_f (new_AGEMA_signal_4602), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_23_U1_X), .Z0_f (new_AGEMA_signal_4969), .Z1_t (new_AGEMA_signal_4970), .Z1_f (new_AGEMA_signal_4971) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_23_U1_X), .B0_f (new_AGEMA_signal_4969), .B1_t (new_AGEMA_signal_4970), .B1_f (new_AGEMA_signal_4971), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_23_U1_Y), .Z0_f (new_AGEMA_signal_5095), .Z1_t (new_AGEMA_signal_5096), .Z1_f (new_AGEMA_signal_5097) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_23_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_23_U1_Y), .A0_f (new_AGEMA_signal_5095), .A1_t (new_AGEMA_signal_5096), .A1_f (new_AGEMA_signal_5097), .B0_t (Midori_rounds_SR_Result[23]), .B0_f (new_AGEMA_signal_4322), .B1_t (new_AGEMA_signal_4323), .B1_f (new_AGEMA_signal_4324), .Z0_t (Midori_rounds_mul_input[23]), .Z0_f (new_AGEMA_signal_5252), .Z1_t (new_AGEMA_signal_5253), .Z1_f (new_AGEMA_signal_5254) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_24_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[24]), .A0_f (new_AGEMA_signal_4754), .A1_t (new_AGEMA_signal_4755), .A1_f (new_AGEMA_signal_4756), .B0_t (Midori_rounds_sub_ResultXORkey[24]), .B0_f (new_AGEMA_signal_5464), .B1_t (new_AGEMA_signal_5465), .B1_f (new_AGEMA_signal_5466), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_24_U1_X), .Z0_f (new_AGEMA_signal_5734), .Z1_t (new_AGEMA_signal_5735), .Z1_f (new_AGEMA_signal_5736) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_24_U1_X), .B0_f (new_AGEMA_signal_5734), .B1_t (new_AGEMA_signal_5735), .B1_f (new_AGEMA_signal_5736), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_24_U1_Y), .Z0_f (new_AGEMA_signal_5867), .Z1_t (new_AGEMA_signal_5868), .Z1_f (new_AGEMA_signal_5869) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_24_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_24_U1_Y), .A0_f (new_AGEMA_signal_5867), .A1_t (new_AGEMA_signal_5868), .A1_f (new_AGEMA_signal_5869), .B0_t (Midori_rounds_SR_Result[24]), .B0_f (new_AGEMA_signal_4754), .B1_t (new_AGEMA_signal_4755), .B1_f (new_AGEMA_signal_4756), .Z0_t (Midori_rounds_mul_input[24]), .Z0_f (new_AGEMA_signal_6002), .Z1_t (new_AGEMA_signal_6003), .Z1_f (new_AGEMA_signal_6004) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_25_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[25]), .A0_f (new_AGEMA_signal_4433), .A1_t (new_AGEMA_signal_4434), .A1_f (new_AGEMA_signal_4435), .B0_t (Midori_rounds_sub_ResultXORkey[25]), .B0_f (new_AGEMA_signal_4651), .B1_t (new_AGEMA_signal_4652), .B1_f (new_AGEMA_signal_4653), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_25_U1_X), .Z0_f (new_AGEMA_signal_4972), .Z1_t (new_AGEMA_signal_4973), .Z1_f (new_AGEMA_signal_4974) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_25_U1_X), .B0_f (new_AGEMA_signal_4972), .B1_t (new_AGEMA_signal_4973), .B1_f (new_AGEMA_signal_4974), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_25_U1_Y), .Z0_f (new_AGEMA_signal_5098), .Z1_t (new_AGEMA_signal_5099), .Z1_f (new_AGEMA_signal_5100) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_25_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_25_U1_Y), .A0_f (new_AGEMA_signal_5098), .A1_t (new_AGEMA_signal_5099), .A1_f (new_AGEMA_signal_5100), .B0_t (Midori_rounds_SR_Result[25]), .B0_f (new_AGEMA_signal_4433), .B1_t (new_AGEMA_signal_4434), .B1_f (new_AGEMA_signal_4435), .Z0_t (Midori_rounds_mul_input[25]), .Z0_f (new_AGEMA_signal_5255), .Z1_t (new_AGEMA_signal_5256), .Z1_f (new_AGEMA_signal_5257) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_26_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[26]), .A0_f (new_AGEMA_signal_4757), .A1_t (new_AGEMA_signal_4758), .A1_f (new_AGEMA_signal_4759), .B0_t (Midori_rounds_sub_ResultXORkey[26]), .B0_f (new_AGEMA_signal_4899), .B1_t (new_AGEMA_signal_4900), .B1_f (new_AGEMA_signal_4901), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_26_U1_X), .Z0_f (new_AGEMA_signal_5101), .Z1_t (new_AGEMA_signal_5102), .Z1_f (new_AGEMA_signal_5103) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_26_U1_X), .B0_f (new_AGEMA_signal_5101), .B1_t (new_AGEMA_signal_5102), .B1_f (new_AGEMA_signal_5103), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_26_U1_Y), .Z0_f (new_AGEMA_signal_5258), .Z1_t (new_AGEMA_signal_5259), .Z1_f (new_AGEMA_signal_5260) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_26_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_26_U1_Y), .A0_f (new_AGEMA_signal_5258), .A1_t (new_AGEMA_signal_5259), .A1_f (new_AGEMA_signal_5260), .B0_t (Midori_rounds_SR_Result[26]), .B0_f (new_AGEMA_signal_4757), .B1_t (new_AGEMA_signal_4758), .B1_f (new_AGEMA_signal_4759), .Z0_t (Midori_rounds_mul_input[26]), .Z0_f (new_AGEMA_signal_5380), .Z1_t (new_AGEMA_signal_5381), .Z1_f (new_AGEMA_signal_5382) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_27_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[27]), .A0_f (new_AGEMA_signal_4430), .A1_t (new_AGEMA_signal_4431), .A1_f (new_AGEMA_signal_4432), .B0_t (Midori_rounds_sub_ResultXORkey[27]), .B0_f (new_AGEMA_signal_4648), .B1_t (new_AGEMA_signal_4649), .B1_f (new_AGEMA_signal_4650), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_27_U1_X), .Z0_f (new_AGEMA_signal_4975), .Z1_t (new_AGEMA_signal_4976), .Z1_f (new_AGEMA_signal_4977) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_27_U1_X), .B0_f (new_AGEMA_signal_4975), .B1_t (new_AGEMA_signal_4976), .B1_f (new_AGEMA_signal_4977), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_27_U1_Y), .Z0_f (new_AGEMA_signal_5104), .Z1_t (new_AGEMA_signal_5105), .Z1_f (new_AGEMA_signal_5106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_27_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_27_U1_Y), .A0_f (new_AGEMA_signal_5104), .A1_t (new_AGEMA_signal_5105), .A1_f (new_AGEMA_signal_5106), .B0_t (Midori_rounds_SR_Result[27]), .B0_f (new_AGEMA_signal_4430), .B1_t (new_AGEMA_signal_4431), .B1_f (new_AGEMA_signal_4432), .Z0_t (Midori_rounds_mul_input[27]), .Z0_f (new_AGEMA_signal_5261), .Z1_t (new_AGEMA_signal_5262), .Z1_f (new_AGEMA_signal_5263) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_28_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[28]), .A0_f (new_AGEMA_signal_4718), .A1_t (new_AGEMA_signal_4719), .A1_f (new_AGEMA_signal_4720), .B0_t (Midori_rounds_sub_ResultXORkey[28]), .B0_f (new_AGEMA_signal_5803), .B1_t (new_AGEMA_signal_5804), .B1_f (new_AGEMA_signal_5805), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_28_U1_X), .Z0_f (new_AGEMA_signal_6005), .Z1_t (new_AGEMA_signal_6006), .Z1_f (new_AGEMA_signal_6007) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_28_U1_X), .B0_f (new_AGEMA_signal_6005), .B1_t (new_AGEMA_signal_6006), .B1_f (new_AGEMA_signal_6007), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_28_U1_Y), .Z0_f (new_AGEMA_signal_6185), .Z1_t (new_AGEMA_signal_6186), .Z1_f (new_AGEMA_signal_6187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_28_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_28_U1_Y), .A0_f (new_AGEMA_signal_6185), .A1_t (new_AGEMA_signal_6186), .A1_f (new_AGEMA_signal_6187), .B0_t (Midori_rounds_SR_Result[28]), .B0_f (new_AGEMA_signal_4718), .B1_t (new_AGEMA_signal_4719), .B1_f (new_AGEMA_signal_4720), .Z0_t (Midori_rounds_mul_input[28]), .Z0_f (new_AGEMA_signal_6464), .Z1_t (new_AGEMA_signal_6465), .Z1_f (new_AGEMA_signal_6466) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_29_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[29]), .A0_f (new_AGEMA_signal_4361), .A1_t (new_AGEMA_signal_4362), .A1_f (new_AGEMA_signal_4363), .B0_t (Midori_rounds_sub_ResultXORkey[29]), .B0_f (new_AGEMA_signal_4627), .B1_t (new_AGEMA_signal_4628), .B1_f (new_AGEMA_signal_4629), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_29_U1_X), .Z0_f (new_AGEMA_signal_4978), .Z1_t (new_AGEMA_signal_4979), .Z1_f (new_AGEMA_signal_4980) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_29_U1_X), .B0_f (new_AGEMA_signal_4978), .B1_t (new_AGEMA_signal_4979), .B1_f (new_AGEMA_signal_4980), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_29_U1_Y), .Z0_f (new_AGEMA_signal_5107), .Z1_t (new_AGEMA_signal_5108), .Z1_f (new_AGEMA_signal_5109) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_29_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_29_U1_Y), .A0_f (new_AGEMA_signal_5107), .A1_t (new_AGEMA_signal_5108), .A1_f (new_AGEMA_signal_5109), .B0_t (Midori_rounds_SR_Result[29]), .B0_f (new_AGEMA_signal_4361), .B1_t (new_AGEMA_signal_4362), .B1_f (new_AGEMA_signal_4363), .Z0_t (Midori_rounds_mul_input[29]), .Z0_f (new_AGEMA_signal_5264), .Z1_t (new_AGEMA_signal_5265), .Z1_f (new_AGEMA_signal_5266) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_30_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[30]), .A0_f (new_AGEMA_signal_4721), .A1_t (new_AGEMA_signal_4722), .A1_f (new_AGEMA_signal_4723), .B0_t (Midori_rounds_sub_ResultXORkey[30]), .B0_f (new_AGEMA_signal_4914), .B1_t (new_AGEMA_signal_4915), .B1_f (new_AGEMA_signal_4916), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_30_U1_X), .Z0_f (new_AGEMA_signal_5110), .Z1_t (new_AGEMA_signal_5111), .Z1_f (new_AGEMA_signal_5112) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_30_U1_X), .B0_f (new_AGEMA_signal_5110), .B1_t (new_AGEMA_signal_5111), .B1_f (new_AGEMA_signal_5112), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_30_U1_Y), .Z0_f (new_AGEMA_signal_5267), .Z1_t (new_AGEMA_signal_5268), .Z1_f (new_AGEMA_signal_5269) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_30_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_30_U1_Y), .A0_f (new_AGEMA_signal_5267), .A1_t (new_AGEMA_signal_5268), .A1_f (new_AGEMA_signal_5269), .B0_t (Midori_rounds_SR_Result[30]), .B0_f (new_AGEMA_signal_4721), .B1_t (new_AGEMA_signal_4722), .B1_f (new_AGEMA_signal_4723), .Z0_t (Midori_rounds_mul_input[30]), .Z0_f (new_AGEMA_signal_5383), .Z1_t (new_AGEMA_signal_5384), .Z1_f (new_AGEMA_signal_5385) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_31_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[31]), .A0_f (new_AGEMA_signal_4358), .A1_t (new_AGEMA_signal_4359), .A1_f (new_AGEMA_signal_4360), .B0_t (Midori_rounds_sub_ResultXORkey[31]), .B0_f (new_AGEMA_signal_4624), .B1_t (new_AGEMA_signal_4625), .B1_f (new_AGEMA_signal_4626), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_31_U1_X), .Z0_f (new_AGEMA_signal_4981), .Z1_t (new_AGEMA_signal_4982), .Z1_f (new_AGEMA_signal_4983) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_31_U1_X), .B0_f (new_AGEMA_signal_4981), .B1_t (new_AGEMA_signal_4982), .B1_f (new_AGEMA_signal_4983), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_31_U1_Y), .Z0_f (new_AGEMA_signal_5113), .Z1_t (new_AGEMA_signal_5114), .Z1_f (new_AGEMA_signal_5115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_31_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_31_U1_Y), .A0_f (new_AGEMA_signal_5113), .A1_t (new_AGEMA_signal_5114), .A1_f (new_AGEMA_signal_5115), .B0_t (Midori_rounds_SR_Result[31]), .B0_f (new_AGEMA_signal_4358), .B1_t (new_AGEMA_signal_4359), .B1_f (new_AGEMA_signal_4360), .Z0_t (Midori_rounds_mul_input[31]), .Z0_f (new_AGEMA_signal_5270), .Z1_t (new_AGEMA_signal_5271), .Z1_f (new_AGEMA_signal_5272) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_32_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[32]), .A0_f (new_AGEMA_signal_4769), .A1_t (new_AGEMA_signal_4770), .A1_f (new_AGEMA_signal_4771), .B0_t (Midori_rounds_sub_ResultXORkey[32]), .B0_f (new_AGEMA_signal_5984), .B1_t (new_AGEMA_signal_5985), .B1_f (new_AGEMA_signal_5986), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_32_U1_X), .Z0_f (new_AGEMA_signal_6188), .Z1_t (new_AGEMA_signal_6189), .Z1_f (new_AGEMA_signal_6190) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_32_U1_X), .B0_f (new_AGEMA_signal_6188), .B1_t (new_AGEMA_signal_6189), .B1_f (new_AGEMA_signal_6190), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_32_U1_Y), .Z0_f (new_AGEMA_signal_6467), .Z1_t (new_AGEMA_signal_6468), .Z1_f (new_AGEMA_signal_6469) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_32_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_32_U1_Y), .A0_f (new_AGEMA_signal_6467), .A1_t (new_AGEMA_signal_6468), .A1_f (new_AGEMA_signal_6469), .B0_t (Midori_rounds_SR_Result[32]), .B0_f (new_AGEMA_signal_4769), .B1_t (new_AGEMA_signal_4770), .B1_f (new_AGEMA_signal_4771), .Z0_t (Midori_rounds_mul_input[32]), .Z0_f (new_AGEMA_signal_6683), .Z1_t (new_AGEMA_signal_6684), .Z1_f (new_AGEMA_signal_6685) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_33_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[33]), .A0_f (new_AGEMA_signal_4451), .A1_t (new_AGEMA_signal_4452), .A1_f (new_AGEMA_signal_4453), .B0_t (Midori_rounds_sub_ResultXORkey[33]), .B0_f (new_AGEMA_signal_4597), .B1_t (new_AGEMA_signal_4598), .B1_f (new_AGEMA_signal_4599), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_33_U1_X), .Z0_f (new_AGEMA_signal_4984), .Z1_t (new_AGEMA_signal_4985), .Z1_f (new_AGEMA_signal_4986) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_33_U1_X), .B0_f (new_AGEMA_signal_4984), .B1_t (new_AGEMA_signal_4985), .B1_f (new_AGEMA_signal_4986), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_33_U1_Y), .Z0_f (new_AGEMA_signal_5116), .Z1_t (new_AGEMA_signal_5117), .Z1_f (new_AGEMA_signal_5118) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_33_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_33_U1_Y), .A0_f (new_AGEMA_signal_5116), .A1_t (new_AGEMA_signal_5117), .A1_f (new_AGEMA_signal_5118), .B0_t (Midori_rounds_SR_Result[33]), .B0_f (new_AGEMA_signal_4451), .B1_t (new_AGEMA_signal_4452), .B1_f (new_AGEMA_signal_4453), .Z0_t (Midori_rounds_mul_input[33]), .Z0_f (new_AGEMA_signal_5273), .Z1_t (new_AGEMA_signal_5274), .Z1_f (new_AGEMA_signal_5275) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_34_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[34]), .A0_f (new_AGEMA_signal_4766), .A1_t (new_AGEMA_signal_4767), .A1_f (new_AGEMA_signal_4768), .B0_t (Midori_rounds_sub_ResultXORkey[34]), .B0_f (new_AGEMA_signal_4878), .B1_t (new_AGEMA_signal_4879), .B1_f (new_AGEMA_signal_4880), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_34_U1_X), .Z0_f (new_AGEMA_signal_5119), .Z1_t (new_AGEMA_signal_5120), .Z1_f (new_AGEMA_signal_5121) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_34_U1_X), .B0_f (new_AGEMA_signal_5119), .B1_t (new_AGEMA_signal_5120), .B1_f (new_AGEMA_signal_5121), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_34_U1_Y), .Z0_f (new_AGEMA_signal_5276), .Z1_t (new_AGEMA_signal_5277), .Z1_f (new_AGEMA_signal_5278) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_34_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_34_U1_Y), .A0_f (new_AGEMA_signal_5276), .A1_t (new_AGEMA_signal_5277), .A1_f (new_AGEMA_signal_5278), .B0_t (Midori_rounds_SR_Result[34]), .B0_f (new_AGEMA_signal_4766), .B1_t (new_AGEMA_signal_4767), .B1_f (new_AGEMA_signal_4768), .Z0_t (Midori_rounds_mul_input[34]), .Z0_f (new_AGEMA_signal_5386), .Z1_t (new_AGEMA_signal_5387), .Z1_f (new_AGEMA_signal_5388) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_35_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[35]), .A0_f (new_AGEMA_signal_4448), .A1_t (new_AGEMA_signal_4449), .A1_f (new_AGEMA_signal_4450), .B0_t (Midori_rounds_sub_ResultXORkey[35]), .B0_f (new_AGEMA_signal_4594), .B1_t (new_AGEMA_signal_4595), .B1_f (new_AGEMA_signal_4596), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_35_U1_X), .Z0_f (new_AGEMA_signal_4987), .Z1_t (new_AGEMA_signal_4988), .Z1_f (new_AGEMA_signal_4989) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_35_U1_X), .B0_f (new_AGEMA_signal_4987), .B1_t (new_AGEMA_signal_4988), .B1_f (new_AGEMA_signal_4989), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_35_U1_Y), .Z0_f (new_AGEMA_signal_5122), .Z1_t (new_AGEMA_signal_5123), .Z1_f (new_AGEMA_signal_5124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_35_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_35_U1_Y), .A0_f (new_AGEMA_signal_5122), .A1_t (new_AGEMA_signal_5123), .A1_f (new_AGEMA_signal_5124), .B0_t (Midori_rounds_SR_Result[35]), .B0_f (new_AGEMA_signal_4448), .B1_t (new_AGEMA_signal_4449), .B1_f (new_AGEMA_signal_4450), .Z0_t (Midori_rounds_mul_input[35]), .Z0_f (new_AGEMA_signal_5279), .Z1_t (new_AGEMA_signal_5280), .Z1_f (new_AGEMA_signal_5281) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_36_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[36]), .A0_f (new_AGEMA_signal_4706), .A1_t (new_AGEMA_signal_4707), .A1_f (new_AGEMA_signal_4708), .B0_t (Midori_rounds_sub_ResultXORkey[36]), .B0_f (new_AGEMA_signal_5794), .B1_t (new_AGEMA_signal_5795), .B1_f (new_AGEMA_signal_5796), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_36_U1_X), .Z0_f (new_AGEMA_signal_6008), .Z1_t (new_AGEMA_signal_6009), .Z1_f (new_AGEMA_signal_6010) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_36_U1_X), .B0_f (new_AGEMA_signal_6008), .B1_t (new_AGEMA_signal_6009), .B1_f (new_AGEMA_signal_6010), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_36_U1_Y), .Z0_f (new_AGEMA_signal_6191), .Z1_t (new_AGEMA_signal_6192), .Z1_f (new_AGEMA_signal_6193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_36_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_36_U1_Y), .A0_f (new_AGEMA_signal_6191), .A1_t (new_AGEMA_signal_6192), .A1_f (new_AGEMA_signal_6193), .B0_t (Midori_rounds_SR_Result[36]), .B0_f (new_AGEMA_signal_4706), .B1_t (new_AGEMA_signal_4707), .B1_f (new_AGEMA_signal_4708), .Z0_t (Midori_rounds_mul_input[36]), .Z0_f (new_AGEMA_signal_6470), .Z1_t (new_AGEMA_signal_6471), .Z1_f (new_AGEMA_signal_6472) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_37_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[37]), .A0_f (new_AGEMA_signal_4337), .A1_t (new_AGEMA_signal_4338), .A1_f (new_AGEMA_signal_4339), .B0_t (Midori_rounds_sub_ResultXORkey[37]), .B0_f (new_AGEMA_signal_4579), .B1_t (new_AGEMA_signal_4580), .B1_f (new_AGEMA_signal_4581), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_37_U1_X), .Z0_f (new_AGEMA_signal_4990), .Z1_t (new_AGEMA_signal_4991), .Z1_f (new_AGEMA_signal_4992) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_37_U1_X), .B0_f (new_AGEMA_signal_4990), .B1_t (new_AGEMA_signal_4991), .B1_f (new_AGEMA_signal_4992), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_37_U1_Y), .Z0_f (new_AGEMA_signal_5125), .Z1_t (new_AGEMA_signal_5126), .Z1_f (new_AGEMA_signal_5127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_37_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_37_U1_Y), .A0_f (new_AGEMA_signal_5125), .A1_t (new_AGEMA_signal_5126), .A1_f (new_AGEMA_signal_5127), .B0_t (Midori_rounds_SR_Result[37]), .B0_f (new_AGEMA_signal_4337), .B1_t (new_AGEMA_signal_4338), .B1_f (new_AGEMA_signal_4339), .Z0_t (Midori_rounds_mul_input[37]), .Z0_f (new_AGEMA_signal_5282), .Z1_t (new_AGEMA_signal_5283), .Z1_f (new_AGEMA_signal_5284) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_38_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[38]), .A0_f (new_AGEMA_signal_4709), .A1_t (new_AGEMA_signal_4710), .A1_f (new_AGEMA_signal_4711), .B0_t (Midori_rounds_sub_ResultXORkey[38]), .B0_f (new_AGEMA_signal_4887), .B1_t (new_AGEMA_signal_4888), .B1_f (new_AGEMA_signal_4889), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_38_U1_X), .Z0_f (new_AGEMA_signal_5128), .Z1_t (new_AGEMA_signal_5129), .Z1_f (new_AGEMA_signal_5130) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_38_U1_X), .B0_f (new_AGEMA_signal_5128), .B1_t (new_AGEMA_signal_5129), .B1_f (new_AGEMA_signal_5130), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_38_U1_Y), .Z0_f (new_AGEMA_signal_5285), .Z1_t (new_AGEMA_signal_5286), .Z1_f (new_AGEMA_signal_5287) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_38_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_38_U1_Y), .A0_f (new_AGEMA_signal_5285), .A1_t (new_AGEMA_signal_5286), .A1_f (new_AGEMA_signal_5287), .B0_t (Midori_rounds_SR_Result[38]), .B0_f (new_AGEMA_signal_4709), .B1_t (new_AGEMA_signal_4710), .B1_f (new_AGEMA_signal_4711), .Z0_t (Midori_rounds_mul_input[38]), .Z0_f (new_AGEMA_signal_5389), .Z1_t (new_AGEMA_signal_5390), .Z1_f (new_AGEMA_signal_5391) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_39_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[39]), .A0_f (new_AGEMA_signal_4334), .A1_t (new_AGEMA_signal_4335), .A1_f (new_AGEMA_signal_4336), .B0_t (Midori_rounds_sub_ResultXORkey[39]), .B0_f (new_AGEMA_signal_4576), .B1_t (new_AGEMA_signal_4577), .B1_f (new_AGEMA_signal_4578), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_39_U1_X), .Z0_f (new_AGEMA_signal_4993), .Z1_t (new_AGEMA_signal_4994), .Z1_f (new_AGEMA_signal_4995) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_39_U1_X), .B0_f (new_AGEMA_signal_4993), .B1_t (new_AGEMA_signal_4994), .B1_f (new_AGEMA_signal_4995), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_39_U1_Y), .Z0_f (new_AGEMA_signal_5131), .Z1_t (new_AGEMA_signal_5132), .Z1_f (new_AGEMA_signal_5133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_39_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_39_U1_Y), .A0_f (new_AGEMA_signal_5131), .A1_t (new_AGEMA_signal_5132), .A1_f (new_AGEMA_signal_5133), .B0_t (Midori_rounds_SR_Result[39]), .B0_f (new_AGEMA_signal_4334), .B1_t (new_AGEMA_signal_4335), .B1_f (new_AGEMA_signal_4336), .Z0_t (Midori_rounds_mul_input[39]), .Z0_f (new_AGEMA_signal_5288), .Z1_t (new_AGEMA_signal_5289), .Z1_f (new_AGEMA_signal_5290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_40_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[40]), .A0_f (new_AGEMA_signal_4748), .A1_t (new_AGEMA_signal_4749), .A1_f (new_AGEMA_signal_4750), .B0_t (Midori_rounds_sub_ResultXORkey[40]), .B0_f (new_AGEMA_signal_5628), .B1_t (new_AGEMA_signal_5629), .B1_f (new_AGEMA_signal_5630), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_40_U1_X), .Z0_f (new_AGEMA_signal_5870), .Z1_t (new_AGEMA_signal_5871), .Z1_f (new_AGEMA_signal_5872) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_40_U1_X), .B0_f (new_AGEMA_signal_5870), .B1_t (new_AGEMA_signal_5871), .B1_f (new_AGEMA_signal_5872), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_40_U1_Y), .Z0_f (new_AGEMA_signal_6011), .Z1_t (new_AGEMA_signal_6012), .Z1_f (new_AGEMA_signal_6013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_40_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_40_U1_Y), .A0_f (new_AGEMA_signal_6011), .A1_t (new_AGEMA_signal_6012), .A1_f (new_AGEMA_signal_6013), .B0_t (Midori_rounds_SR_Result[40]), .B0_f (new_AGEMA_signal_4748), .B1_t (new_AGEMA_signal_4749), .B1_f (new_AGEMA_signal_4750), .Z0_t (Midori_rounds_mul_input[40]), .Z0_f (new_AGEMA_signal_6194), .Z1_t (new_AGEMA_signal_6195), .Z1_f (new_AGEMA_signal_6196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_41_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[41]), .A0_f (new_AGEMA_signal_4421), .A1_t (new_AGEMA_signal_4422), .A1_f (new_AGEMA_signal_4423), .B0_t (Midori_rounds_sub_ResultXORkey[41]), .B0_f (new_AGEMA_signal_4621), .B1_t (new_AGEMA_signal_4622), .B1_f (new_AGEMA_signal_4623), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_41_U1_X), .Z0_f (new_AGEMA_signal_4996), .Z1_t (new_AGEMA_signal_4997), .Z1_f (new_AGEMA_signal_4998) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_41_U1_X), .B0_f (new_AGEMA_signal_4996), .B1_t (new_AGEMA_signal_4997), .B1_f (new_AGEMA_signal_4998), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_41_U1_Y), .Z0_f (new_AGEMA_signal_5134), .Z1_t (new_AGEMA_signal_5135), .Z1_f (new_AGEMA_signal_5136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_41_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_41_U1_Y), .A0_f (new_AGEMA_signal_5134), .A1_t (new_AGEMA_signal_5135), .A1_f (new_AGEMA_signal_5136), .B0_t (Midori_rounds_SR_Result[41]), .B0_f (new_AGEMA_signal_4421), .B1_t (new_AGEMA_signal_4422), .B1_f (new_AGEMA_signal_4423), .Z0_t (Midori_rounds_mul_input[41]), .Z0_f (new_AGEMA_signal_5291), .Z1_t (new_AGEMA_signal_5292), .Z1_f (new_AGEMA_signal_5293) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_42_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[42]), .A0_f (new_AGEMA_signal_4751), .A1_t (new_AGEMA_signal_4752), .A1_f (new_AGEMA_signal_4753), .B0_t (Midori_rounds_sub_ResultXORkey[42]), .B0_f (new_AGEMA_signal_4905), .B1_t (new_AGEMA_signal_4906), .B1_f (new_AGEMA_signal_4907), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_42_U1_X), .Z0_f (new_AGEMA_signal_5137), .Z1_t (new_AGEMA_signal_5138), .Z1_f (new_AGEMA_signal_5139) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_42_U1_X), .B0_f (new_AGEMA_signal_5137), .B1_t (new_AGEMA_signal_5138), .B1_f (new_AGEMA_signal_5139), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_42_U1_Y), .Z0_f (new_AGEMA_signal_5294), .Z1_t (new_AGEMA_signal_5295), .Z1_f (new_AGEMA_signal_5296) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_42_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_42_U1_Y), .A0_f (new_AGEMA_signal_5294), .A1_t (new_AGEMA_signal_5295), .A1_f (new_AGEMA_signal_5296), .B0_t (Midori_rounds_SR_Result[42]), .B0_f (new_AGEMA_signal_4751), .B1_t (new_AGEMA_signal_4752), .B1_f (new_AGEMA_signal_4753), .Z0_t (Midori_rounds_mul_input[42]), .Z0_f (new_AGEMA_signal_5392), .Z1_t (new_AGEMA_signal_5393), .Z1_f (new_AGEMA_signal_5394) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_43_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[43]), .A0_f (new_AGEMA_signal_4418), .A1_t (new_AGEMA_signal_4419), .A1_f (new_AGEMA_signal_4420), .B0_t (Midori_rounds_sub_ResultXORkey[43]), .B0_f (new_AGEMA_signal_4618), .B1_t (new_AGEMA_signal_4619), .B1_f (new_AGEMA_signal_4620), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_43_U1_X), .Z0_f (new_AGEMA_signal_4999), .Z1_t (new_AGEMA_signal_5000), .Z1_f (new_AGEMA_signal_5001) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_43_U1_X), .B0_f (new_AGEMA_signal_4999), .B1_t (new_AGEMA_signal_5000), .B1_f (new_AGEMA_signal_5001), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_43_U1_Y), .Z0_f (new_AGEMA_signal_5140), .Z1_t (new_AGEMA_signal_5141), .Z1_f (new_AGEMA_signal_5142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_43_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_43_U1_Y), .A0_f (new_AGEMA_signal_5140), .A1_t (new_AGEMA_signal_5141), .A1_f (new_AGEMA_signal_5142), .B0_t (Midori_rounds_SR_Result[43]), .B0_f (new_AGEMA_signal_4418), .B1_t (new_AGEMA_signal_4419), .B1_f (new_AGEMA_signal_4420), .Z0_t (Midori_rounds_mul_input[43]), .Z0_f (new_AGEMA_signal_5297), .Z1_t (new_AGEMA_signal_5298), .Z1_f (new_AGEMA_signal_5299) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_44_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[44]), .A0_f (new_AGEMA_signal_4688), .A1_t (new_AGEMA_signal_4689), .A1_f (new_AGEMA_signal_4690), .B0_t (Midori_rounds_sub_ResultXORkey[44]), .B0_f (new_AGEMA_signal_5345), .B1_t (new_AGEMA_signal_5346), .B1_f (new_AGEMA_signal_5347), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_44_U1_X), .Z0_f (new_AGEMA_signal_5481), .Z1_t (new_AGEMA_signal_5482), .Z1_f (new_AGEMA_signal_5483) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_44_U1_X), .B0_f (new_AGEMA_signal_5481), .B1_t (new_AGEMA_signal_5482), .B1_f (new_AGEMA_signal_5483), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_44_U1_Y), .Z0_f (new_AGEMA_signal_5737), .Z1_t (new_AGEMA_signal_5738), .Z1_f (new_AGEMA_signal_5739) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_44_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_44_U1_Y), .A0_f (new_AGEMA_signal_5737), .A1_t (new_AGEMA_signal_5738), .A1_f (new_AGEMA_signal_5739), .B0_t (Midori_rounds_SR_Result[44]), .B0_f (new_AGEMA_signal_4688), .B1_t (new_AGEMA_signal_4689), .B1_f (new_AGEMA_signal_4690), .Z0_t (Midori_rounds_mul_input[44]), .Z0_f (new_AGEMA_signal_5873), .Z1_t (new_AGEMA_signal_5874), .Z1_f (new_AGEMA_signal_5875) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_45_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[45]), .A0_f (new_AGEMA_signal_4301), .A1_t (new_AGEMA_signal_4302), .A1_f (new_AGEMA_signal_4303), .B0_t (Midori_rounds_sub_ResultXORkey[45]), .B0_f (new_AGEMA_signal_4645), .B1_t (new_AGEMA_signal_4646), .B1_f (new_AGEMA_signal_4647), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_45_U1_X), .Z0_f (new_AGEMA_signal_5002), .Z1_t (new_AGEMA_signal_5003), .Z1_f (new_AGEMA_signal_5004) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_45_U1_X), .B0_f (new_AGEMA_signal_5002), .B1_t (new_AGEMA_signal_5003), .B1_f (new_AGEMA_signal_5004), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_45_U1_Y), .Z0_f (new_AGEMA_signal_5143), .Z1_t (new_AGEMA_signal_5144), .Z1_f (new_AGEMA_signal_5145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_45_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_45_U1_Y), .A0_f (new_AGEMA_signal_5143), .A1_t (new_AGEMA_signal_5144), .A1_f (new_AGEMA_signal_5145), .B0_t (Midori_rounds_SR_Result[45]), .B0_f (new_AGEMA_signal_4301), .B1_t (new_AGEMA_signal_4302), .B1_f (new_AGEMA_signal_4303), .Z0_t (Midori_rounds_mul_input[45]), .Z0_f (new_AGEMA_signal_5300), .Z1_t (new_AGEMA_signal_5301), .Z1_f (new_AGEMA_signal_5302) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_46_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[46]), .A0_f (new_AGEMA_signal_4691), .A1_t (new_AGEMA_signal_4692), .A1_f (new_AGEMA_signal_4693), .B0_t (Midori_rounds_sub_ResultXORkey[46]), .B0_f (new_AGEMA_signal_4911), .B1_t (new_AGEMA_signal_4912), .B1_f (new_AGEMA_signal_4913), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_46_U1_X), .Z0_f (new_AGEMA_signal_5146), .Z1_t (new_AGEMA_signal_5147), .Z1_f (new_AGEMA_signal_5148) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_46_U1_X), .B0_f (new_AGEMA_signal_5146), .B1_t (new_AGEMA_signal_5147), .B1_f (new_AGEMA_signal_5148), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_46_U1_Y), .Z0_f (new_AGEMA_signal_5303), .Z1_t (new_AGEMA_signal_5304), .Z1_f (new_AGEMA_signal_5305) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_46_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_46_U1_Y), .A0_f (new_AGEMA_signal_5303), .A1_t (new_AGEMA_signal_5304), .A1_f (new_AGEMA_signal_5305), .B0_t (Midori_rounds_SR_Result[46]), .B0_f (new_AGEMA_signal_4691), .B1_t (new_AGEMA_signal_4692), .B1_f (new_AGEMA_signal_4693), .Z0_t (Midori_rounds_mul_input[46]), .Z0_f (new_AGEMA_signal_5395), .Z1_t (new_AGEMA_signal_5396), .Z1_f (new_AGEMA_signal_5397) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_47_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[47]), .A0_f (new_AGEMA_signal_4298), .A1_t (new_AGEMA_signal_4299), .A1_f (new_AGEMA_signal_4300), .B0_t (Midori_rounds_sub_ResultXORkey[47]), .B0_f (new_AGEMA_signal_4642), .B1_t (new_AGEMA_signal_4643), .B1_f (new_AGEMA_signal_4644), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_47_U1_X), .Z0_f (new_AGEMA_signal_5005), .Z1_t (new_AGEMA_signal_5006), .Z1_f (new_AGEMA_signal_5007) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_47_U1_X), .B0_f (new_AGEMA_signal_5005), .B1_t (new_AGEMA_signal_5006), .B1_f (new_AGEMA_signal_5007), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_47_U1_Y), .Z0_f (new_AGEMA_signal_5149), .Z1_t (new_AGEMA_signal_5150), .Z1_f (new_AGEMA_signal_5151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_47_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_47_U1_Y), .A0_f (new_AGEMA_signal_5149), .A1_t (new_AGEMA_signal_5150), .A1_f (new_AGEMA_signal_5151), .B0_t (Midori_rounds_SR_Result[47]), .B0_f (new_AGEMA_signal_4298), .B1_t (new_AGEMA_signal_4299), .B1_f (new_AGEMA_signal_4300), .Z0_t (Midori_rounds_mul_input[47]), .Z0_f (new_AGEMA_signal_5306), .Z1_t (new_AGEMA_signal_5307), .Z1_f (new_AGEMA_signal_5308) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_48_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[48]), .A0_f (new_AGEMA_signal_4685), .A1_t (new_AGEMA_signal_4686), .A1_f (new_AGEMA_signal_4687), .B0_t (Midori_rounds_sub_ResultXORkey[48]), .B0_f (new_AGEMA_signal_5981), .B1_t (new_AGEMA_signal_5982), .B1_f (new_AGEMA_signal_5983), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_48_U1_X), .Z0_f (new_AGEMA_signal_6197), .Z1_t (new_AGEMA_signal_6198), .Z1_f (new_AGEMA_signal_6199) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_48_U1_X), .B0_f (new_AGEMA_signal_6197), .B1_t (new_AGEMA_signal_6198), .B1_f (new_AGEMA_signal_6199), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_48_U1_Y), .Z0_f (new_AGEMA_signal_6473), .Z1_t (new_AGEMA_signal_6474), .Z1_f (new_AGEMA_signal_6475) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_48_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_48_U1_Y), .A0_f (new_AGEMA_signal_6473), .A1_t (new_AGEMA_signal_6474), .A1_f (new_AGEMA_signal_6475), .B0_t (Midori_rounds_SR_Result[48]), .B0_f (new_AGEMA_signal_4685), .B1_t (new_AGEMA_signal_4686), .B1_f (new_AGEMA_signal_4687), .Z0_t (Midori_rounds_mul_input[48]), .Z0_f (new_AGEMA_signal_6686), .Z1_t (new_AGEMA_signal_6687), .Z1_f (new_AGEMA_signal_6688) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_49_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[49]), .A0_f (new_AGEMA_signal_4283), .A1_t (new_AGEMA_signal_4284), .A1_f (new_AGEMA_signal_4285), .B0_t (Midori_rounds_sub_ResultXORkey[49]), .B0_f (new_AGEMA_signal_4573), .B1_t (new_AGEMA_signal_4574), .B1_f (new_AGEMA_signal_4575), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_49_U1_X), .Z0_f (new_AGEMA_signal_5008), .Z1_t (new_AGEMA_signal_5009), .Z1_f (new_AGEMA_signal_5010) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_49_U1_X), .B0_f (new_AGEMA_signal_5008), .B1_t (new_AGEMA_signal_5009), .B1_f (new_AGEMA_signal_5010), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_49_U1_Y), .Z0_f (new_AGEMA_signal_5152), .Z1_t (new_AGEMA_signal_5153), .Z1_f (new_AGEMA_signal_5154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_49_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_49_U1_Y), .A0_f (new_AGEMA_signal_5152), .A1_t (new_AGEMA_signal_5153), .A1_f (new_AGEMA_signal_5154), .B0_t (Midori_rounds_SR_Result[49]), .B0_f (new_AGEMA_signal_4283), .B1_t (new_AGEMA_signal_4284), .B1_f (new_AGEMA_signal_4285), .Z0_t (Midori_rounds_mul_input[49]), .Z0_f (new_AGEMA_signal_5309), .Z1_t (new_AGEMA_signal_5310), .Z1_f (new_AGEMA_signal_5311) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_50_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[50]), .A0_f (new_AGEMA_signal_4682), .A1_t (new_AGEMA_signal_4683), .A1_f (new_AGEMA_signal_4684), .B0_t (Midori_rounds_sub_ResultXORkey[50]), .B0_f (new_AGEMA_signal_4884), .B1_t (new_AGEMA_signal_4885), .B1_f (new_AGEMA_signal_4886), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_50_U1_X), .Z0_f (new_AGEMA_signal_5155), .Z1_t (new_AGEMA_signal_5156), .Z1_f (new_AGEMA_signal_5157) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_50_U1_X), .B0_f (new_AGEMA_signal_5155), .B1_t (new_AGEMA_signal_5156), .B1_f (new_AGEMA_signal_5157), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_50_U1_Y), .Z0_f (new_AGEMA_signal_5312), .Z1_t (new_AGEMA_signal_5313), .Z1_f (new_AGEMA_signal_5314) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_50_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_50_U1_Y), .A0_f (new_AGEMA_signal_5312), .A1_t (new_AGEMA_signal_5313), .A1_f (new_AGEMA_signal_5314), .B0_t (Midori_rounds_SR_Result[50]), .B0_f (new_AGEMA_signal_4682), .B1_t (new_AGEMA_signal_4683), .B1_f (new_AGEMA_signal_4684), .Z0_t (Midori_rounds_mul_input[50]), .Z0_f (new_AGEMA_signal_5398), .Z1_t (new_AGEMA_signal_5399), .Z1_f (new_AGEMA_signal_5400) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_51_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[51]), .A0_f (new_AGEMA_signal_4280), .A1_t (new_AGEMA_signal_4281), .A1_f (new_AGEMA_signal_4282), .B0_t (Midori_rounds_sub_ResultXORkey[51]), .B0_f (new_AGEMA_signal_4570), .B1_t (new_AGEMA_signal_4571), .B1_f (new_AGEMA_signal_4572), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_51_U1_X), .Z0_f (new_AGEMA_signal_5011), .Z1_t (new_AGEMA_signal_5012), .Z1_f (new_AGEMA_signal_5013) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_51_U1_X), .B0_f (new_AGEMA_signal_5011), .B1_t (new_AGEMA_signal_5012), .B1_f (new_AGEMA_signal_5013), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_51_U1_Y), .Z0_f (new_AGEMA_signal_5158), .Z1_t (new_AGEMA_signal_5159), .Z1_f (new_AGEMA_signal_5160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_51_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_51_U1_Y), .A0_f (new_AGEMA_signal_5158), .A1_t (new_AGEMA_signal_5159), .A1_f (new_AGEMA_signal_5160), .B0_t (Midori_rounds_SR_Result[51]), .B0_f (new_AGEMA_signal_4280), .B1_t (new_AGEMA_signal_4281), .B1_f (new_AGEMA_signal_4282), .Z0_t (Midori_rounds_mul_input[51]), .Z0_f (new_AGEMA_signal_5315), .Z1_t (new_AGEMA_signal_5316), .Z1_f (new_AGEMA_signal_5317) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_52_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[52]), .A0_f (new_AGEMA_signal_4742), .A1_t (new_AGEMA_signal_4743), .A1_f (new_AGEMA_signal_4744), .B0_t (Midori_rounds_sub_ResultXORkey[52]), .B0_f (new_AGEMA_signal_5788), .B1_t (new_AGEMA_signal_5789), .B1_f (new_AGEMA_signal_5790), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_52_U1_X), .Z0_f (new_AGEMA_signal_6014), .Z1_t (new_AGEMA_signal_6015), .Z1_f (new_AGEMA_signal_6016) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_52_U1_X), .B0_f (new_AGEMA_signal_6014), .B1_t (new_AGEMA_signal_6015), .B1_f (new_AGEMA_signal_6016), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_52_U1_Y), .Z0_f (new_AGEMA_signal_6200), .Z1_t (new_AGEMA_signal_6201), .Z1_f (new_AGEMA_signal_6202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_52_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_52_U1_Y), .A0_f (new_AGEMA_signal_6200), .A1_t (new_AGEMA_signal_6201), .A1_f (new_AGEMA_signal_6202), .B0_t (Midori_rounds_SR_Result[52]), .B0_f (new_AGEMA_signal_4742), .B1_t (new_AGEMA_signal_4743), .B1_f (new_AGEMA_signal_4744), .Z0_t (Midori_rounds_mul_input[52]), .Z0_f (new_AGEMA_signal_6476), .Z1_t (new_AGEMA_signal_6477), .Z1_f (new_AGEMA_signal_6478) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_53_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[53]), .A0_f (new_AGEMA_signal_4409), .A1_t (new_AGEMA_signal_4410), .A1_f (new_AGEMA_signal_4411), .B0_t (Midori_rounds_sub_ResultXORkey[53]), .B0_f (new_AGEMA_signal_4591), .B1_t (new_AGEMA_signal_4592), .B1_f (new_AGEMA_signal_4593), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_53_U1_X), .Z0_f (new_AGEMA_signal_5014), .Z1_t (new_AGEMA_signal_5015), .Z1_f (new_AGEMA_signal_5016) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_53_U1_X), .B0_f (new_AGEMA_signal_5014), .B1_t (new_AGEMA_signal_5015), .B1_f (new_AGEMA_signal_5016), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_53_U1_Y), .Z0_f (new_AGEMA_signal_5161), .Z1_t (new_AGEMA_signal_5162), .Z1_f (new_AGEMA_signal_5163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_53_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_53_U1_Y), .A0_f (new_AGEMA_signal_5161), .A1_t (new_AGEMA_signal_5162), .A1_f (new_AGEMA_signal_5163), .B0_t (Midori_rounds_SR_Result[53]), .B0_f (new_AGEMA_signal_4409), .B1_t (new_AGEMA_signal_4410), .B1_f (new_AGEMA_signal_4411), .Z0_t (Midori_rounds_mul_input[53]), .Z0_f (new_AGEMA_signal_5318), .Z1_t (new_AGEMA_signal_5319), .Z1_f (new_AGEMA_signal_5320) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_54_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[54]), .A0_f (new_AGEMA_signal_4745), .A1_t (new_AGEMA_signal_4746), .A1_f (new_AGEMA_signal_4747), .B0_t (Midori_rounds_sub_ResultXORkey[54]), .B0_f (new_AGEMA_signal_4875), .B1_t (new_AGEMA_signal_4876), .B1_f (new_AGEMA_signal_4877), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_54_U1_X), .Z0_f (new_AGEMA_signal_5164), .Z1_t (new_AGEMA_signal_5165), .Z1_f (new_AGEMA_signal_5166) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_54_U1_X), .B0_f (new_AGEMA_signal_5164), .B1_t (new_AGEMA_signal_5165), .B1_f (new_AGEMA_signal_5166), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_54_U1_Y), .Z0_f (new_AGEMA_signal_5321), .Z1_t (new_AGEMA_signal_5322), .Z1_f (new_AGEMA_signal_5323) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_54_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_54_U1_Y), .A0_f (new_AGEMA_signal_5321), .A1_t (new_AGEMA_signal_5322), .A1_f (new_AGEMA_signal_5323), .B0_t (Midori_rounds_SR_Result[54]), .B0_f (new_AGEMA_signal_4745), .B1_t (new_AGEMA_signal_4746), .B1_f (new_AGEMA_signal_4747), .Z0_t (Midori_rounds_mul_input[54]), .Z0_f (new_AGEMA_signal_5401), .Z1_t (new_AGEMA_signal_5402), .Z1_f (new_AGEMA_signal_5403) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_55_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[55]), .A0_f (new_AGEMA_signal_4406), .A1_t (new_AGEMA_signal_4407), .A1_f (new_AGEMA_signal_4408), .B0_t (Midori_rounds_sub_ResultXORkey[55]), .B0_f (new_AGEMA_signal_4588), .B1_t (new_AGEMA_signal_4589), .B1_f (new_AGEMA_signal_4590), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_55_U1_X), .Z0_f (new_AGEMA_signal_5017), .Z1_t (new_AGEMA_signal_5018), .Z1_f (new_AGEMA_signal_5019) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_55_U1_X), .B0_f (new_AGEMA_signal_5017), .B1_t (new_AGEMA_signal_5018), .B1_f (new_AGEMA_signal_5019), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_55_U1_Y), .Z0_f (new_AGEMA_signal_5167), .Z1_t (new_AGEMA_signal_5168), .Z1_f (new_AGEMA_signal_5169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_55_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_55_U1_Y), .A0_f (new_AGEMA_signal_5167), .A1_t (new_AGEMA_signal_5168), .A1_f (new_AGEMA_signal_5169), .B0_t (Midori_rounds_SR_Result[55]), .B0_f (new_AGEMA_signal_4406), .B1_t (new_AGEMA_signal_4407), .B1_f (new_AGEMA_signal_4408), .Z0_t (Midori_rounds_mul_input[55]), .Z0_f (new_AGEMA_signal_5324), .Z1_t (new_AGEMA_signal_5325), .Z1_f (new_AGEMA_signal_5326) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_56_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[56]), .A0_f (new_AGEMA_signal_4712), .A1_t (new_AGEMA_signal_4713), .A1_f (new_AGEMA_signal_4714), .B0_t (Midori_rounds_sub_ResultXORkey[56]), .B0_f (new_AGEMA_signal_5607), .B1_t (new_AGEMA_signal_5608), .B1_f (new_AGEMA_signal_5609), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_56_U1_X), .Z0_f (new_AGEMA_signal_5876), .Z1_t (new_AGEMA_signal_5877), .Z1_f (new_AGEMA_signal_5878) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_56_U1_X), .B0_f (new_AGEMA_signal_5876), .B1_t (new_AGEMA_signal_5877), .B1_f (new_AGEMA_signal_5878), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_56_U1_Y), .Z0_f (new_AGEMA_signal_6017), .Z1_t (new_AGEMA_signal_6018), .Z1_f (new_AGEMA_signal_6019) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_56_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_56_U1_Y), .A0_f (new_AGEMA_signal_6017), .A1_t (new_AGEMA_signal_6018), .A1_f (new_AGEMA_signal_6019), .B0_t (Midori_rounds_SR_Result[56]), .B0_f (new_AGEMA_signal_4712), .B1_t (new_AGEMA_signal_4713), .B1_f (new_AGEMA_signal_4714), .Z0_t (Midori_rounds_mul_input[56]), .Z0_f (new_AGEMA_signal_6203), .Z1_t (new_AGEMA_signal_6204), .Z1_f (new_AGEMA_signal_6205) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_57_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[57]), .A0_f (new_AGEMA_signal_4349), .A1_t (new_AGEMA_signal_4350), .A1_f (new_AGEMA_signal_4351), .B0_t (Midori_rounds_sub_ResultXORkey[57]), .B0_f (new_AGEMA_signal_4639), .B1_t (new_AGEMA_signal_4640), .B1_f (new_AGEMA_signal_4641), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_57_U1_X), .Z0_f (new_AGEMA_signal_5020), .Z1_t (new_AGEMA_signal_5021), .Z1_f (new_AGEMA_signal_5022) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_57_U1_X), .B0_f (new_AGEMA_signal_5020), .B1_t (new_AGEMA_signal_5021), .B1_f (new_AGEMA_signal_5022), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_57_U1_Y), .Z0_f (new_AGEMA_signal_5170), .Z1_t (new_AGEMA_signal_5171), .Z1_f (new_AGEMA_signal_5172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_57_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_57_U1_Y), .A0_f (new_AGEMA_signal_5170), .A1_t (new_AGEMA_signal_5171), .A1_f (new_AGEMA_signal_5172), .B0_t (Midori_rounds_SR_Result[57]), .B0_f (new_AGEMA_signal_4349), .B1_t (new_AGEMA_signal_4350), .B1_f (new_AGEMA_signal_4351), .Z0_t (Midori_rounds_mul_input[57]), .Z0_f (new_AGEMA_signal_5327), .Z1_t (new_AGEMA_signal_5328), .Z1_f (new_AGEMA_signal_5329) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_58_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[58]), .A0_f (new_AGEMA_signal_4715), .A1_t (new_AGEMA_signal_4716), .A1_f (new_AGEMA_signal_4717), .B0_t (Midori_rounds_sub_ResultXORkey[58]), .B0_f (new_AGEMA_signal_4908), .B1_t (new_AGEMA_signal_4909), .B1_f (new_AGEMA_signal_4910), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_58_U1_X), .Z0_f (new_AGEMA_signal_5173), .Z1_t (new_AGEMA_signal_5174), .Z1_f (new_AGEMA_signal_5175) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_58_U1_X), .B0_f (new_AGEMA_signal_5173), .B1_t (new_AGEMA_signal_5174), .B1_f (new_AGEMA_signal_5175), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_58_U1_Y), .Z0_f (new_AGEMA_signal_5330), .Z1_t (new_AGEMA_signal_5331), .Z1_f (new_AGEMA_signal_5332) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_58_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_58_U1_Y), .A0_f (new_AGEMA_signal_5330), .A1_t (new_AGEMA_signal_5331), .A1_f (new_AGEMA_signal_5332), .B0_t (Midori_rounds_SR_Result[58]), .B0_f (new_AGEMA_signal_4715), .B1_t (new_AGEMA_signal_4716), .B1_f (new_AGEMA_signal_4717), .Z0_t (Midori_rounds_mul_input[58]), .Z0_f (new_AGEMA_signal_5404), .Z1_t (new_AGEMA_signal_5405), .Z1_f (new_AGEMA_signal_5406) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_59_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[59]), .A0_f (new_AGEMA_signal_4346), .A1_t (new_AGEMA_signal_4347), .A1_f (new_AGEMA_signal_4348), .B0_t (Midori_rounds_sub_ResultXORkey[59]), .B0_f (new_AGEMA_signal_4636), .B1_t (new_AGEMA_signal_4637), .B1_f (new_AGEMA_signal_4638), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_59_U1_X), .Z0_f (new_AGEMA_signal_5023), .Z1_t (new_AGEMA_signal_5024), .Z1_f (new_AGEMA_signal_5025) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_59_U1_X), .B0_f (new_AGEMA_signal_5023), .B1_t (new_AGEMA_signal_5024), .B1_f (new_AGEMA_signal_5025), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_59_U1_Y), .Z0_f (new_AGEMA_signal_5176), .Z1_t (new_AGEMA_signal_5177), .Z1_f (new_AGEMA_signal_5178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_59_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_59_U1_Y), .A0_f (new_AGEMA_signal_5176), .A1_t (new_AGEMA_signal_5177), .A1_f (new_AGEMA_signal_5178), .B0_t (Midori_rounds_SR_Result[59]), .B0_f (new_AGEMA_signal_4346), .B1_t (new_AGEMA_signal_4347), .B1_f (new_AGEMA_signal_4348), .Z0_t (Midori_rounds_mul_input[59]), .Z0_f (new_AGEMA_signal_5333), .Z1_t (new_AGEMA_signal_5334), .Z1_f (new_AGEMA_signal_5335) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_60_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[60]), .A0_f (new_AGEMA_signal_4772), .A1_t (new_AGEMA_signal_4773), .A1_f (new_AGEMA_signal_4774), .B0_t (Midori_rounds_sub_ResultXORkey[60]), .B0_f (new_AGEMA_signal_5604), .B1_t (new_AGEMA_signal_5605), .B1_f (new_AGEMA_signal_5606), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_60_U1_X), .Z0_f (new_AGEMA_signal_5879), .Z1_t (new_AGEMA_signal_5880), .Z1_f (new_AGEMA_signal_5881) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_60_U1_X), .B0_f (new_AGEMA_signal_5879), .B1_t (new_AGEMA_signal_5880), .B1_f (new_AGEMA_signal_5881), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_60_U1_Y), .Z0_f (new_AGEMA_signal_6020), .Z1_t (new_AGEMA_signal_6021), .Z1_f (new_AGEMA_signal_6022) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_60_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_60_U1_Y), .A0_f (new_AGEMA_signal_6020), .A1_t (new_AGEMA_signal_6021), .A1_f (new_AGEMA_signal_6022), .B0_t (Midori_rounds_SR_Result[60]), .B0_f (new_AGEMA_signal_4772), .B1_t (new_AGEMA_signal_4773), .B1_f (new_AGEMA_signal_4774), .Z0_t (Midori_rounds_mul_input[60]), .Z0_f (new_AGEMA_signal_6206), .Z1_t (new_AGEMA_signal_6207), .Z1_f (new_AGEMA_signal_6208) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_61_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[61]), .A0_f (new_AGEMA_signal_4469), .A1_t (new_AGEMA_signal_4470), .A1_f (new_AGEMA_signal_4471), .B0_t (Midori_rounds_sub_ResultXORkey[61]), .B0_f (new_AGEMA_signal_4633), .B1_t (new_AGEMA_signal_4634), .B1_f (new_AGEMA_signal_4635), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_61_U1_X), .Z0_f (new_AGEMA_signal_5026), .Z1_t (new_AGEMA_signal_5027), .Z1_f (new_AGEMA_signal_5028) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_61_U1_X), .B0_f (new_AGEMA_signal_5026), .B1_t (new_AGEMA_signal_5027), .B1_f (new_AGEMA_signal_5028), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_61_U1_Y), .Z0_f (new_AGEMA_signal_5179), .Z1_t (new_AGEMA_signal_5180), .Z1_f (new_AGEMA_signal_5181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_61_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_61_U1_Y), .A0_f (new_AGEMA_signal_5179), .A1_t (new_AGEMA_signal_5180), .A1_f (new_AGEMA_signal_5181), .B0_t (Midori_rounds_SR_Result[61]), .B0_f (new_AGEMA_signal_4469), .B1_t (new_AGEMA_signal_4470), .B1_f (new_AGEMA_signal_4471), .Z0_t (Midori_rounds_mul_input[61]), .Z0_f (new_AGEMA_signal_5336), .Z1_t (new_AGEMA_signal_5337), .Z1_f (new_AGEMA_signal_5338) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_62_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[62]), .A0_f (new_AGEMA_signal_4775), .A1_t (new_AGEMA_signal_4776), .A1_f (new_AGEMA_signal_4777), .B0_t (Midori_rounds_sub_ResultXORkey[62]), .B0_f (new_AGEMA_signal_4902), .B1_t (new_AGEMA_signal_4903), .B1_f (new_AGEMA_signal_4904), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_62_U1_X), .Z0_f (new_AGEMA_signal_5182), .Z1_t (new_AGEMA_signal_5183), .Z1_f (new_AGEMA_signal_5184) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_62_U1_X), .B0_f (new_AGEMA_signal_5182), .B1_t (new_AGEMA_signal_5183), .B1_f (new_AGEMA_signal_5184), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_62_U1_Y), .Z0_f (new_AGEMA_signal_5339), .Z1_t (new_AGEMA_signal_5340), .Z1_f (new_AGEMA_signal_5341) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_62_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_62_U1_Y), .A0_f (new_AGEMA_signal_5339), .A1_t (new_AGEMA_signal_5340), .A1_f (new_AGEMA_signal_5341), .B0_t (Midori_rounds_SR_Result[62]), .B0_f (new_AGEMA_signal_4775), .B1_t (new_AGEMA_signal_4776), .B1_f (new_AGEMA_signal_4777), .Z0_t (Midori_rounds_mul_input[62]), .Z0_f (new_AGEMA_signal_5407), .Z1_t (new_AGEMA_signal_5408), .Z1_f (new_AGEMA_signal_5409) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_63_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[63]), .A0_f (new_AGEMA_signal_4466), .A1_t (new_AGEMA_signal_4467), .A1_f (new_AGEMA_signal_4468), .B0_t (Midori_rounds_sub_ResultXORkey[63]), .B0_f (new_AGEMA_signal_4630), .B1_t (new_AGEMA_signal_4631), .B1_f (new_AGEMA_signal_4632), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_63_U1_X), .Z0_f (new_AGEMA_signal_5029), .Z1_t (new_AGEMA_signal_5030), .Z1_f (new_AGEMA_signal_5031) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_63_U1_X), .B0_f (new_AGEMA_signal_5029), .B1_t (new_AGEMA_signal_5030), .B1_f (new_AGEMA_signal_5031), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_63_U1_Y), .Z0_f (new_AGEMA_signal_5185), .Z1_t (new_AGEMA_signal_5186), .Z1_f (new_AGEMA_signal_5187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_63_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_63_U1_Y), .A0_f (new_AGEMA_signal_5185), .A1_t (new_AGEMA_signal_5186), .A1_f (new_AGEMA_signal_5187), .B0_t (Midori_rounds_SR_Result[63]), .B0_f (new_AGEMA_signal_4466), .B1_t (new_AGEMA_signal_4467), .B1_f (new_AGEMA_signal_4468), .Z0_t (Midori_rounds_mul_input[63]), .Z0_f (new_AGEMA_signal_5342), .Z1_t (new_AGEMA_signal_5343), .Z1_f (new_AGEMA_signal_5344) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U24 ( .A0_t (Midori_rounds_mul_input[59]), .A0_f (new_AGEMA_signal_5333), .A1_t (new_AGEMA_signal_5334), .A1_f (new_AGEMA_signal_5335), .B0_t (Midori_rounds_mul_MC1_n8), .B0_f (new_AGEMA_signal_5410), .B1_t (new_AGEMA_signal_5411), .B1_f (new_AGEMA_signal_5412), .Z0_t (Midori_rounds_SR_Inv_Result[63]), .Z0_f (new_AGEMA_signal_5484), .Z1_t (new_AGEMA_signal_5485), .Z1_f (new_AGEMA_signal_5486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U23 ( .A0_t (Midori_rounds_mul_input[63]), .A0_f (new_AGEMA_signal_5342), .A1_t (new_AGEMA_signal_5343), .A1_f (new_AGEMA_signal_5344), .B0_t (Midori_rounds_mul_MC1_n8), .B0_f (new_AGEMA_signal_5410), .B1_t (new_AGEMA_signal_5411), .B1_f (new_AGEMA_signal_5412), .Z0_t (Midori_rounds_SR_Inv_Result[23]), .Z0_f (new_AGEMA_signal_5487), .Z1_t (new_AGEMA_signal_5488), .Z1_f (new_AGEMA_signal_5489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U22 ( .A0_t (Midori_rounds_mul_input[55]), .A0_f (new_AGEMA_signal_5324), .A1_t (new_AGEMA_signal_5325), .A1_f (new_AGEMA_signal_5326), .B0_t (Midori_rounds_mul_input[51]), .B0_f (new_AGEMA_signal_5315), .B1_t (new_AGEMA_signal_5316), .B1_f (new_AGEMA_signal_5317), .Z0_t (Midori_rounds_mul_MC1_n8), .Z0_f (new_AGEMA_signal_5410), .Z1_t (new_AGEMA_signal_5411), .Z1_f (new_AGEMA_signal_5412) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U21 ( .A0_t (Midori_rounds_mul_input[58]), .A0_f (new_AGEMA_signal_5404), .A1_t (new_AGEMA_signal_5405), .A1_f (new_AGEMA_signal_5406), .B0_t (Midori_rounds_mul_MC1_n7), .B0_f (new_AGEMA_signal_5490), .B1_t (new_AGEMA_signal_5491), .B1_f (new_AGEMA_signal_5492), .Z0_t (Midori_rounds_SR_Inv_Result[62]), .Z0_f (new_AGEMA_signal_5740), .Z1_t (new_AGEMA_signal_5741), .Z1_f (new_AGEMA_signal_5742) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U20 ( .A0_t (Midori_rounds_mul_input[62]), .A0_f (new_AGEMA_signal_5407), .A1_t (new_AGEMA_signal_5408), .A1_f (new_AGEMA_signal_5409), .B0_t (Midori_rounds_mul_MC1_n7), .B0_f (new_AGEMA_signal_5490), .B1_t (new_AGEMA_signal_5491), .B1_f (new_AGEMA_signal_5492), .Z0_t (Midori_rounds_SR_Inv_Result[22]), .Z0_f (new_AGEMA_signal_5743), .Z1_t (new_AGEMA_signal_5744), .Z1_f (new_AGEMA_signal_5745) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U19 ( .A0_t (Midori_rounds_mul_input[54]), .A0_f (new_AGEMA_signal_5401), .A1_t (new_AGEMA_signal_5402), .A1_f (new_AGEMA_signal_5403), .B0_t (Midori_rounds_mul_input[50]), .B0_f (new_AGEMA_signal_5398), .B1_t (new_AGEMA_signal_5399), .B1_f (new_AGEMA_signal_5400), .Z0_t (Midori_rounds_mul_MC1_n7), .Z0_f (new_AGEMA_signal_5490), .Z1_t (new_AGEMA_signal_5491), .Z1_f (new_AGEMA_signal_5492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U18 ( .A0_t (Midori_rounds_mul_input[56]), .A0_f (new_AGEMA_signal_6203), .A1_t (new_AGEMA_signal_6204), .A1_f (new_AGEMA_signal_6205), .B0_t (Midori_rounds_mul_MC1_n6), .B0_f (new_AGEMA_signal_6758), .B1_t (new_AGEMA_signal_6759), .B1_f (new_AGEMA_signal_6760), .Z0_t (Midori_rounds_SR_Inv_Result[60]), .Z0_f (new_AGEMA_signal_6797), .Z1_t (new_AGEMA_signal_6798), .Z1_f (new_AGEMA_signal_6799) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U17 ( .A0_t (Midori_rounds_mul_input[60]), .A0_f (new_AGEMA_signal_6206), .A1_t (new_AGEMA_signal_6207), .A1_f (new_AGEMA_signal_6208), .B0_t (Midori_rounds_mul_MC1_n6), .B0_f (new_AGEMA_signal_6758), .B1_t (new_AGEMA_signal_6759), .B1_f (new_AGEMA_signal_6760), .Z0_t (Midori_rounds_SR_Inv_Result[20]), .Z0_f (new_AGEMA_signal_6800), .Z1_t (new_AGEMA_signal_6801), .Z1_f (new_AGEMA_signal_6802) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U16 ( .A0_t (Midori_rounds_mul_input[52]), .A0_f (new_AGEMA_signal_6476), .A1_t (new_AGEMA_signal_6477), .A1_f (new_AGEMA_signal_6478), .B0_t (Midori_rounds_mul_input[48]), .B0_f (new_AGEMA_signal_6686), .B1_t (new_AGEMA_signal_6687), .B1_f (new_AGEMA_signal_6688), .Z0_t (Midori_rounds_mul_MC1_n6), .Z0_f (new_AGEMA_signal_6758), .Z1_t (new_AGEMA_signal_6759), .Z1_f (new_AGEMA_signal_6760) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U15 ( .A0_t (Midori_rounds_mul_input[51]), .A0_f (new_AGEMA_signal_5315), .A1_t (new_AGEMA_signal_5316), .A1_f (new_AGEMA_signal_5317), .B0_t (Midori_rounds_mul_MC1_n5), .B0_f (new_AGEMA_signal_5413), .B1_t (new_AGEMA_signal_5414), .B1_f (new_AGEMA_signal_5415), .Z0_t (Midori_rounds_SR_Inv_Result[43]), .Z0_f (new_AGEMA_signal_5493), .Z1_t (new_AGEMA_signal_5494), .Z1_f (new_AGEMA_signal_5495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U14 ( .A0_t (Midori_rounds_mul_input[55]), .A0_f (new_AGEMA_signal_5324), .A1_t (new_AGEMA_signal_5325), .A1_f (new_AGEMA_signal_5326), .B0_t (Midori_rounds_mul_MC1_n5), .B0_f (new_AGEMA_signal_5413), .B1_t (new_AGEMA_signal_5414), .B1_f (new_AGEMA_signal_5415), .Z0_t (Midori_rounds_SR_Inv_Result[3]), .Z0_f (new_AGEMA_signal_5496), .Z1_t (new_AGEMA_signal_5497), .Z1_f (new_AGEMA_signal_5498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U13 ( .A0_t (Midori_rounds_mul_input[59]), .A0_f (new_AGEMA_signal_5333), .A1_t (new_AGEMA_signal_5334), .A1_f (new_AGEMA_signal_5335), .B0_t (Midori_rounds_mul_input[63]), .B0_f (new_AGEMA_signal_5342), .B1_t (new_AGEMA_signal_5343), .B1_f (new_AGEMA_signal_5344), .Z0_t (Midori_rounds_mul_MC1_n5), .Z0_f (new_AGEMA_signal_5413), .Z1_t (new_AGEMA_signal_5414), .Z1_f (new_AGEMA_signal_5415) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U12 ( .A0_t (Midori_rounds_mul_input[57]), .A0_f (new_AGEMA_signal_5327), .A1_t (new_AGEMA_signal_5328), .A1_f (new_AGEMA_signal_5329), .B0_t (Midori_rounds_mul_MC1_n4), .B0_f (new_AGEMA_signal_5416), .B1_t (new_AGEMA_signal_5417), .B1_f (new_AGEMA_signal_5418), .Z0_t (Midori_rounds_SR_Inv_Result[61]), .Z0_f (new_AGEMA_signal_5499), .Z1_t (new_AGEMA_signal_5500), .Z1_f (new_AGEMA_signal_5501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U11 ( .A0_t (Midori_rounds_mul_input[61]), .A0_f (new_AGEMA_signal_5336), .A1_t (new_AGEMA_signal_5337), .A1_f (new_AGEMA_signal_5338), .B0_t (Midori_rounds_mul_MC1_n4), .B0_f (new_AGEMA_signal_5416), .B1_t (new_AGEMA_signal_5417), .B1_f (new_AGEMA_signal_5418), .Z0_t (Midori_rounds_SR_Inv_Result[21]), .Z0_f (new_AGEMA_signal_5502), .Z1_t (new_AGEMA_signal_5503), .Z1_f (new_AGEMA_signal_5504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U10 ( .A0_t (Midori_rounds_mul_input[53]), .A0_f (new_AGEMA_signal_5318), .A1_t (new_AGEMA_signal_5319), .A1_f (new_AGEMA_signal_5320), .B0_t (Midori_rounds_mul_input[49]), .B0_f (new_AGEMA_signal_5309), .B1_t (new_AGEMA_signal_5310), .B1_f (new_AGEMA_signal_5311), .Z0_t (Midori_rounds_mul_MC1_n4), .Z0_f (new_AGEMA_signal_5416), .Z1_t (new_AGEMA_signal_5417), .Z1_f (new_AGEMA_signal_5418) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U9 ( .A0_t (Midori_rounds_mul_input[50]), .A0_f (new_AGEMA_signal_5398), .A1_t (new_AGEMA_signal_5399), .A1_f (new_AGEMA_signal_5400), .B0_t (Midori_rounds_mul_MC1_n3), .B0_f (new_AGEMA_signal_5505), .B1_t (new_AGEMA_signal_5506), .B1_f (new_AGEMA_signal_5507), .Z0_t (Midori_rounds_SR_Inv_Result[42]), .Z0_f (new_AGEMA_signal_5746), .Z1_t (new_AGEMA_signal_5747), .Z1_f (new_AGEMA_signal_5748) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U8 ( .A0_t (Midori_rounds_mul_input[54]), .A0_f (new_AGEMA_signal_5401), .A1_t (new_AGEMA_signal_5402), .A1_f (new_AGEMA_signal_5403), .B0_t (Midori_rounds_mul_MC1_n3), .B0_f (new_AGEMA_signal_5505), .B1_t (new_AGEMA_signal_5506), .B1_f (new_AGEMA_signal_5507), .Z0_t (Midori_rounds_SR_Inv_Result[2]), .Z0_f (new_AGEMA_signal_5749), .Z1_t (new_AGEMA_signal_5750), .Z1_f (new_AGEMA_signal_5751) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U7 ( .A0_t (Midori_rounds_mul_input[58]), .A0_f (new_AGEMA_signal_5404), .A1_t (new_AGEMA_signal_5405), .A1_f (new_AGEMA_signal_5406), .B0_t (Midori_rounds_mul_input[62]), .B0_f (new_AGEMA_signal_5407), .B1_t (new_AGEMA_signal_5408), .B1_f (new_AGEMA_signal_5409), .Z0_t (Midori_rounds_mul_MC1_n3), .Z0_f (new_AGEMA_signal_5505), .Z1_t (new_AGEMA_signal_5506), .Z1_f (new_AGEMA_signal_5507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U6 ( .A0_t (Midori_rounds_mul_input[49]), .A0_f (new_AGEMA_signal_5309), .A1_t (new_AGEMA_signal_5310), .A1_f (new_AGEMA_signal_5311), .B0_t (Midori_rounds_mul_MC1_n2), .B0_f (new_AGEMA_signal_5419), .B1_t (new_AGEMA_signal_5420), .B1_f (new_AGEMA_signal_5421), .Z0_t (Midori_rounds_SR_Inv_Result[41]), .Z0_f (new_AGEMA_signal_5508), .Z1_t (new_AGEMA_signal_5509), .Z1_f (new_AGEMA_signal_5510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U5 ( .A0_t (Midori_rounds_mul_input[53]), .A0_f (new_AGEMA_signal_5318), .A1_t (new_AGEMA_signal_5319), .A1_f (new_AGEMA_signal_5320), .B0_t (Midori_rounds_mul_MC1_n2), .B0_f (new_AGEMA_signal_5419), .B1_t (new_AGEMA_signal_5420), .B1_f (new_AGEMA_signal_5421), .Z0_t (Midori_rounds_SR_Inv_Result[1]), .Z0_f (new_AGEMA_signal_5511), .Z1_t (new_AGEMA_signal_5512), .Z1_f (new_AGEMA_signal_5513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U4 ( .A0_t (Midori_rounds_mul_input[57]), .A0_f (new_AGEMA_signal_5327), .A1_t (new_AGEMA_signal_5328), .A1_f (new_AGEMA_signal_5329), .B0_t (Midori_rounds_mul_input[61]), .B0_f (new_AGEMA_signal_5336), .B1_t (new_AGEMA_signal_5337), .B1_f (new_AGEMA_signal_5338), .Z0_t (Midori_rounds_mul_MC1_n2), .Z0_f (new_AGEMA_signal_5419), .Z1_t (new_AGEMA_signal_5420), .Z1_f (new_AGEMA_signal_5421) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U3 ( .A0_t (Midori_rounds_mul_input[48]), .A0_f (new_AGEMA_signal_6686), .A1_t (new_AGEMA_signal_6687), .A1_f (new_AGEMA_signal_6688), .B0_t (Midori_rounds_mul_MC1_n1), .B0_f (new_AGEMA_signal_6479), .B1_t (new_AGEMA_signal_6480), .B1_f (new_AGEMA_signal_6481), .Z0_t (Midori_rounds_SR_Inv_Result[40]), .Z0_f (new_AGEMA_signal_6761), .Z1_t (new_AGEMA_signal_6762), .Z1_f (new_AGEMA_signal_6763) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U2 ( .A0_t (Midori_rounds_mul_input[52]), .A0_f (new_AGEMA_signal_6476), .A1_t (new_AGEMA_signal_6477), .A1_f (new_AGEMA_signal_6478), .B0_t (Midori_rounds_mul_MC1_n1), .B0_f (new_AGEMA_signal_6479), .B1_t (new_AGEMA_signal_6480), .B1_f (new_AGEMA_signal_6481), .Z0_t (Midori_rounds_SR_Inv_Result[0]), .Z0_f (new_AGEMA_signal_6689), .Z1_t (new_AGEMA_signal_6690), .Z1_f (new_AGEMA_signal_6691) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U1 ( .A0_t (Midori_rounds_mul_input[56]), .A0_f (new_AGEMA_signal_6203), .A1_t (new_AGEMA_signal_6204), .A1_f (new_AGEMA_signal_6205), .B0_t (Midori_rounds_mul_input[60]), .B0_f (new_AGEMA_signal_6206), .B1_t (new_AGEMA_signal_6207), .B1_f (new_AGEMA_signal_6208), .Z0_t (Midori_rounds_mul_MC1_n1), .Z0_f (new_AGEMA_signal_6479), .Z1_t (new_AGEMA_signal_6480), .Z1_f (new_AGEMA_signal_6481) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U24 ( .A0_t (Midori_rounds_mul_input[43]), .A0_f (new_AGEMA_signal_5297), .A1_t (new_AGEMA_signal_5298), .A1_f (new_AGEMA_signal_5299), .B0_t (Midori_rounds_mul_MC2_n8), .B0_f (new_AGEMA_signal_5422), .B1_t (new_AGEMA_signal_5423), .B1_f (new_AGEMA_signal_5424), .Z0_t (Midori_rounds_SR_Inv_Result[7]), .Z0_f (new_AGEMA_signal_5514), .Z1_t (new_AGEMA_signal_5515), .Z1_f (new_AGEMA_signal_5516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U23 ( .A0_t (Midori_rounds_mul_input[47]), .A0_f (new_AGEMA_signal_5306), .A1_t (new_AGEMA_signal_5307), .A1_f (new_AGEMA_signal_5308), .B0_t (Midori_rounds_mul_MC2_n8), .B0_f (new_AGEMA_signal_5422), .B1_t (new_AGEMA_signal_5423), .B1_f (new_AGEMA_signal_5424), .Z0_t (Midori_rounds_SR_Inv_Result[47]), .Z0_f (new_AGEMA_signal_5517), .Z1_t (new_AGEMA_signal_5518), .Z1_f (new_AGEMA_signal_5519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U22 ( .A0_t (Midori_rounds_mul_input[39]), .A0_f (new_AGEMA_signal_5288), .A1_t (new_AGEMA_signal_5289), .A1_f (new_AGEMA_signal_5290), .B0_t (Midori_rounds_mul_input[35]), .B0_f (new_AGEMA_signal_5279), .B1_t (new_AGEMA_signal_5280), .B1_f (new_AGEMA_signal_5281), .Z0_t (Midori_rounds_mul_MC2_n8), .Z0_f (new_AGEMA_signal_5422), .Z1_t (new_AGEMA_signal_5423), .Z1_f (new_AGEMA_signal_5424) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U21 ( .A0_t (Midori_rounds_mul_input[42]), .A0_f (new_AGEMA_signal_5392), .A1_t (new_AGEMA_signal_5393), .A1_f (new_AGEMA_signal_5394), .B0_t (Midori_rounds_mul_MC2_n7), .B0_f (new_AGEMA_signal_5520), .B1_t (new_AGEMA_signal_5521), .B1_f (new_AGEMA_signal_5522), .Z0_t (Midori_rounds_SR_Inv_Result[6]), .Z0_f (new_AGEMA_signal_5752), .Z1_t (new_AGEMA_signal_5753), .Z1_f (new_AGEMA_signal_5754) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U20 ( .A0_t (Midori_rounds_mul_input[46]), .A0_f (new_AGEMA_signal_5395), .A1_t (new_AGEMA_signal_5396), .A1_f (new_AGEMA_signal_5397), .B0_t (Midori_rounds_mul_MC2_n7), .B0_f (new_AGEMA_signal_5520), .B1_t (new_AGEMA_signal_5521), .B1_f (new_AGEMA_signal_5522), .Z0_t (Midori_rounds_SR_Inv_Result[46]), .Z0_f (new_AGEMA_signal_5755), .Z1_t (new_AGEMA_signal_5756), .Z1_f (new_AGEMA_signal_5757) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U19 ( .A0_t (Midori_rounds_mul_input[38]), .A0_f (new_AGEMA_signal_5389), .A1_t (new_AGEMA_signal_5390), .A1_f (new_AGEMA_signal_5391), .B0_t (Midori_rounds_mul_input[34]), .B0_f (new_AGEMA_signal_5386), .B1_t (new_AGEMA_signal_5387), .B1_f (new_AGEMA_signal_5388), .Z0_t (Midori_rounds_mul_MC2_n7), .Z0_f (new_AGEMA_signal_5520), .Z1_t (new_AGEMA_signal_5521), .Z1_f (new_AGEMA_signal_5522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U18 ( .A0_t (Midori_rounds_mul_input[40]), .A0_f (new_AGEMA_signal_6194), .A1_t (new_AGEMA_signal_6195), .A1_f (new_AGEMA_signal_6196), .B0_t (Midori_rounds_mul_MC2_n6), .B0_f (new_AGEMA_signal_6764), .B1_t (new_AGEMA_signal_6765), .B1_f (new_AGEMA_signal_6766), .Z0_t (Midori_rounds_SR_Inv_Result[4]), .Z0_f (new_AGEMA_signal_6803), .Z1_t (new_AGEMA_signal_6804), .Z1_f (new_AGEMA_signal_6805) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U17 ( .A0_t (Midori_rounds_mul_input[44]), .A0_f (new_AGEMA_signal_5873), .A1_t (new_AGEMA_signal_5874), .A1_f (new_AGEMA_signal_5875), .B0_t (Midori_rounds_mul_MC2_n6), .B0_f (new_AGEMA_signal_6764), .B1_t (new_AGEMA_signal_6765), .B1_f (new_AGEMA_signal_6766), .Z0_t (Midori_rounds_SR_Inv_Result[44]), .Z0_f (new_AGEMA_signal_6806), .Z1_t (new_AGEMA_signal_6807), .Z1_f (new_AGEMA_signal_6808) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U16 ( .A0_t (Midori_rounds_mul_input[36]), .A0_f (new_AGEMA_signal_6470), .A1_t (new_AGEMA_signal_6471), .A1_f (new_AGEMA_signal_6472), .B0_t (Midori_rounds_mul_input[32]), .B0_f (new_AGEMA_signal_6683), .B1_t (new_AGEMA_signal_6684), .B1_f (new_AGEMA_signal_6685), .Z0_t (Midori_rounds_mul_MC2_n6), .Z0_f (new_AGEMA_signal_6764), .Z1_t (new_AGEMA_signal_6765), .Z1_f (new_AGEMA_signal_6766) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U15 ( .A0_t (Midori_rounds_mul_input[35]), .A0_f (new_AGEMA_signal_5279), .A1_t (new_AGEMA_signal_5280), .A1_f (new_AGEMA_signal_5281), .B0_t (Midori_rounds_mul_MC2_n5), .B0_f (new_AGEMA_signal_5425), .B1_t (new_AGEMA_signal_5426), .B1_f (new_AGEMA_signal_5427), .Z0_t (Midori_rounds_SR_Inv_Result[19]), .Z0_f (new_AGEMA_signal_5523), .Z1_t (new_AGEMA_signal_5524), .Z1_f (new_AGEMA_signal_5525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U14 ( .A0_t (Midori_rounds_mul_input[39]), .A0_f (new_AGEMA_signal_5288), .A1_t (new_AGEMA_signal_5289), .A1_f (new_AGEMA_signal_5290), .B0_t (Midori_rounds_mul_MC2_n5), .B0_f (new_AGEMA_signal_5425), .B1_t (new_AGEMA_signal_5426), .B1_f (new_AGEMA_signal_5427), .Z0_t (Midori_rounds_SR_Inv_Result[59]), .Z0_f (new_AGEMA_signal_5526), .Z1_t (new_AGEMA_signal_5527), .Z1_f (new_AGEMA_signal_5528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U13 ( .A0_t (Midori_rounds_mul_input[43]), .A0_f (new_AGEMA_signal_5297), .A1_t (new_AGEMA_signal_5298), .A1_f (new_AGEMA_signal_5299), .B0_t (Midori_rounds_mul_input[47]), .B0_f (new_AGEMA_signal_5306), .B1_t (new_AGEMA_signal_5307), .B1_f (new_AGEMA_signal_5308), .Z0_t (Midori_rounds_mul_MC2_n5), .Z0_f (new_AGEMA_signal_5425), .Z1_t (new_AGEMA_signal_5426), .Z1_f (new_AGEMA_signal_5427) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U12 ( .A0_t (Midori_rounds_mul_input[41]), .A0_f (new_AGEMA_signal_5291), .A1_t (new_AGEMA_signal_5292), .A1_f (new_AGEMA_signal_5293), .B0_t (Midori_rounds_mul_MC2_n4), .B0_f (new_AGEMA_signal_5428), .B1_t (new_AGEMA_signal_5429), .B1_f (new_AGEMA_signal_5430), .Z0_t (Midori_rounds_SR_Inv_Result[5]), .Z0_f (new_AGEMA_signal_5529), .Z1_t (new_AGEMA_signal_5530), .Z1_f (new_AGEMA_signal_5531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U11 ( .A0_t (Midori_rounds_mul_input[45]), .A0_f (new_AGEMA_signal_5300), .A1_t (new_AGEMA_signal_5301), .A1_f (new_AGEMA_signal_5302), .B0_t (Midori_rounds_mul_MC2_n4), .B0_f (new_AGEMA_signal_5428), .B1_t (new_AGEMA_signal_5429), .B1_f (new_AGEMA_signal_5430), .Z0_t (Midori_rounds_SR_Inv_Result[45]), .Z0_f (new_AGEMA_signal_5532), .Z1_t (new_AGEMA_signal_5533), .Z1_f (new_AGEMA_signal_5534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U10 ( .A0_t (Midori_rounds_mul_input[37]), .A0_f (new_AGEMA_signal_5282), .A1_t (new_AGEMA_signal_5283), .A1_f (new_AGEMA_signal_5284), .B0_t (Midori_rounds_mul_input[33]), .B0_f (new_AGEMA_signal_5273), .B1_t (new_AGEMA_signal_5274), .B1_f (new_AGEMA_signal_5275), .Z0_t (Midori_rounds_mul_MC2_n4), .Z0_f (new_AGEMA_signal_5428), .Z1_t (new_AGEMA_signal_5429), .Z1_f (new_AGEMA_signal_5430) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U9 ( .A0_t (Midori_rounds_mul_input[34]), .A0_f (new_AGEMA_signal_5386), .A1_t (new_AGEMA_signal_5387), .A1_f (new_AGEMA_signal_5388), .B0_t (Midori_rounds_mul_MC2_n3), .B0_f (new_AGEMA_signal_5535), .B1_t (new_AGEMA_signal_5536), .B1_f (new_AGEMA_signal_5537), .Z0_t (Midori_rounds_SR_Inv_Result[18]), .Z0_f (new_AGEMA_signal_5758), .Z1_t (new_AGEMA_signal_5759), .Z1_f (new_AGEMA_signal_5760) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U8 ( .A0_t (Midori_rounds_mul_input[38]), .A0_f (new_AGEMA_signal_5389), .A1_t (new_AGEMA_signal_5390), .A1_f (new_AGEMA_signal_5391), .B0_t (Midori_rounds_mul_MC2_n3), .B0_f (new_AGEMA_signal_5535), .B1_t (new_AGEMA_signal_5536), .B1_f (new_AGEMA_signal_5537), .Z0_t (Midori_rounds_SR_Inv_Result[58]), .Z0_f (new_AGEMA_signal_5761), .Z1_t (new_AGEMA_signal_5762), .Z1_f (new_AGEMA_signal_5763) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U7 ( .A0_t (Midori_rounds_mul_input[42]), .A0_f (new_AGEMA_signal_5392), .A1_t (new_AGEMA_signal_5393), .A1_f (new_AGEMA_signal_5394), .B0_t (Midori_rounds_mul_input[46]), .B0_f (new_AGEMA_signal_5395), .B1_t (new_AGEMA_signal_5396), .B1_f (new_AGEMA_signal_5397), .Z0_t (Midori_rounds_mul_MC2_n3), .Z0_f (new_AGEMA_signal_5535), .Z1_t (new_AGEMA_signal_5536), .Z1_f (new_AGEMA_signal_5537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U6 ( .A0_t (Midori_rounds_mul_input[33]), .A0_f (new_AGEMA_signal_5273), .A1_t (new_AGEMA_signal_5274), .A1_f (new_AGEMA_signal_5275), .B0_t (Midori_rounds_mul_MC2_n2), .B0_f (new_AGEMA_signal_5431), .B1_t (new_AGEMA_signal_5432), .B1_f (new_AGEMA_signal_5433), .Z0_t (Midori_rounds_SR_Inv_Result[17]), .Z0_f (new_AGEMA_signal_5538), .Z1_t (new_AGEMA_signal_5539), .Z1_f (new_AGEMA_signal_5540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U5 ( .A0_t (Midori_rounds_mul_input[37]), .A0_f (new_AGEMA_signal_5282), .A1_t (new_AGEMA_signal_5283), .A1_f (new_AGEMA_signal_5284), .B0_t (Midori_rounds_mul_MC2_n2), .B0_f (new_AGEMA_signal_5431), .B1_t (new_AGEMA_signal_5432), .B1_f (new_AGEMA_signal_5433), .Z0_t (Midori_rounds_SR_Inv_Result[57]), .Z0_f (new_AGEMA_signal_5541), .Z1_t (new_AGEMA_signal_5542), .Z1_f (new_AGEMA_signal_5543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U4 ( .A0_t (Midori_rounds_mul_input[41]), .A0_f (new_AGEMA_signal_5291), .A1_t (new_AGEMA_signal_5292), .A1_f (new_AGEMA_signal_5293), .B0_t (Midori_rounds_mul_input[45]), .B0_f (new_AGEMA_signal_5300), .B1_t (new_AGEMA_signal_5301), .B1_f (new_AGEMA_signal_5302), .Z0_t (Midori_rounds_mul_MC2_n2), .Z0_f (new_AGEMA_signal_5431), .Z1_t (new_AGEMA_signal_5432), .Z1_f (new_AGEMA_signal_5433) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U3 ( .A0_t (Midori_rounds_mul_input[32]), .A0_f (new_AGEMA_signal_6683), .A1_t (new_AGEMA_signal_6684), .A1_f (new_AGEMA_signal_6685), .B0_t (Midori_rounds_mul_MC2_n1), .B0_f (new_AGEMA_signal_6482), .B1_t (new_AGEMA_signal_6483), .B1_f (new_AGEMA_signal_6484), .Z0_t (Midori_rounds_SR_Inv_Result[16]), .Z0_f (new_AGEMA_signal_6767), .Z1_t (new_AGEMA_signal_6768), .Z1_f (new_AGEMA_signal_6769) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U2 ( .A0_t (Midori_rounds_mul_input[36]), .A0_f (new_AGEMA_signal_6470), .A1_t (new_AGEMA_signal_6471), .A1_f (new_AGEMA_signal_6472), .B0_t (Midori_rounds_mul_MC2_n1), .B0_f (new_AGEMA_signal_6482), .B1_t (new_AGEMA_signal_6483), .B1_f (new_AGEMA_signal_6484), .Z0_t (Midori_rounds_SR_Inv_Result[56]), .Z0_f (new_AGEMA_signal_6692), .Z1_t (new_AGEMA_signal_6693), .Z1_f (new_AGEMA_signal_6694) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U1 ( .A0_t (Midori_rounds_mul_input[40]), .A0_f (new_AGEMA_signal_6194), .A1_t (new_AGEMA_signal_6195), .A1_f (new_AGEMA_signal_6196), .B0_t (Midori_rounds_mul_input[44]), .B0_f (new_AGEMA_signal_5873), .B1_t (new_AGEMA_signal_5874), .B1_f (new_AGEMA_signal_5875), .Z0_t (Midori_rounds_mul_MC2_n1), .Z0_f (new_AGEMA_signal_6482), .Z1_t (new_AGEMA_signal_6483), .Z1_f (new_AGEMA_signal_6484) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U24 ( .A0_t (Midori_rounds_mul_input[27]), .A0_f (new_AGEMA_signal_5261), .A1_t (new_AGEMA_signal_5262), .A1_f (new_AGEMA_signal_5263), .B0_t (Midori_rounds_mul_MC3_n8), .B0_f (new_AGEMA_signal_5434), .B1_t (new_AGEMA_signal_5435), .B1_f (new_AGEMA_signal_5436), .Z0_t (Midori_rounds_SR_Inv_Result[27]), .Z0_f (new_AGEMA_signal_5544), .Z1_t (new_AGEMA_signal_5545), .Z1_f (new_AGEMA_signal_5546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U23 ( .A0_t (Midori_rounds_mul_input[31]), .A0_f (new_AGEMA_signal_5270), .A1_t (new_AGEMA_signal_5271), .A1_f (new_AGEMA_signal_5272), .B0_t (Midori_rounds_mul_MC3_n8), .B0_f (new_AGEMA_signal_5434), .B1_t (new_AGEMA_signal_5435), .B1_f (new_AGEMA_signal_5436), .Z0_t (Midori_rounds_SR_Inv_Result[51]), .Z0_f (new_AGEMA_signal_5547), .Z1_t (new_AGEMA_signal_5548), .Z1_f (new_AGEMA_signal_5549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U22 ( .A0_t (Midori_rounds_mul_input[23]), .A0_f (new_AGEMA_signal_5252), .A1_t (new_AGEMA_signal_5253), .A1_f (new_AGEMA_signal_5254), .B0_t (Midori_rounds_mul_input[19]), .B0_f (new_AGEMA_signal_5243), .B1_t (new_AGEMA_signal_5244), .B1_f (new_AGEMA_signal_5245), .Z0_t (Midori_rounds_mul_MC3_n8), .Z0_f (new_AGEMA_signal_5434), .Z1_t (new_AGEMA_signal_5435), .Z1_f (new_AGEMA_signal_5436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U21 ( .A0_t (Midori_rounds_mul_input[26]), .A0_f (new_AGEMA_signal_5380), .A1_t (new_AGEMA_signal_5381), .A1_f (new_AGEMA_signal_5382), .B0_t (Midori_rounds_mul_MC3_n7), .B0_f (new_AGEMA_signal_5550), .B1_t (new_AGEMA_signal_5551), .B1_f (new_AGEMA_signal_5552), .Z0_t (Midori_rounds_SR_Inv_Result[26]), .Z0_f (new_AGEMA_signal_5764), .Z1_t (new_AGEMA_signal_5765), .Z1_f (new_AGEMA_signal_5766) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U20 ( .A0_t (Midori_rounds_mul_input[30]), .A0_f (new_AGEMA_signal_5383), .A1_t (new_AGEMA_signal_5384), .A1_f (new_AGEMA_signal_5385), .B0_t (Midori_rounds_mul_MC3_n7), .B0_f (new_AGEMA_signal_5550), .B1_t (new_AGEMA_signal_5551), .B1_f (new_AGEMA_signal_5552), .Z0_t (Midori_rounds_SR_Inv_Result[50]), .Z0_f (new_AGEMA_signal_5767), .Z1_t (new_AGEMA_signal_5768), .Z1_f (new_AGEMA_signal_5769) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U19 ( .A0_t (Midori_rounds_mul_input[22]), .A0_f (new_AGEMA_signal_5377), .A1_t (new_AGEMA_signal_5378), .A1_f (new_AGEMA_signal_5379), .B0_t (Midori_rounds_mul_input[18]), .B0_f (new_AGEMA_signal_5374), .B1_t (new_AGEMA_signal_5375), .B1_f (new_AGEMA_signal_5376), .Z0_t (Midori_rounds_mul_MC3_n7), .Z0_f (new_AGEMA_signal_5550), .Z1_t (new_AGEMA_signal_5551), .Z1_f (new_AGEMA_signal_5552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U18 ( .A0_t (Midori_rounds_mul_input[24]), .A0_f (new_AGEMA_signal_6002), .A1_t (new_AGEMA_signal_6003), .A1_f (new_AGEMA_signal_6004), .B0_t (Midori_rounds_mul_MC3_n6), .B0_f (new_AGEMA_signal_6770), .B1_t (new_AGEMA_signal_6771), .B1_f (new_AGEMA_signal_6772), .Z0_t (Midori_rounds_SR_Inv_Result[24]), .Z0_f (new_AGEMA_signal_6809), .Z1_t (new_AGEMA_signal_6810), .Z1_f (new_AGEMA_signal_6811) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U17 ( .A0_t (Midori_rounds_mul_input[28]), .A0_f (new_AGEMA_signal_6464), .A1_t (new_AGEMA_signal_6465), .A1_f (new_AGEMA_signal_6466), .B0_t (Midori_rounds_mul_MC3_n6), .B0_f (new_AGEMA_signal_6770), .B1_t (new_AGEMA_signal_6771), .B1_f (new_AGEMA_signal_6772), .Z0_t (Midori_rounds_SR_Inv_Result[48]), .Z0_f (new_AGEMA_signal_6812), .Z1_t (new_AGEMA_signal_6813), .Z1_f (new_AGEMA_signal_6814) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U16 ( .A0_t (Midori_rounds_mul_input[20]), .A0_f (new_AGEMA_signal_6182), .A1_t (new_AGEMA_signal_6183), .A1_f (new_AGEMA_signal_6184), .B0_t (Midori_rounds_mul_input[16]), .B0_f (new_AGEMA_signal_6680), .B1_t (new_AGEMA_signal_6681), .B1_f (new_AGEMA_signal_6682), .Z0_t (Midori_rounds_mul_MC3_n6), .Z0_f (new_AGEMA_signal_6770), .Z1_t (new_AGEMA_signal_6771), .Z1_f (new_AGEMA_signal_6772) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U15 ( .A0_t (Midori_rounds_mul_input[19]), .A0_f (new_AGEMA_signal_5243), .A1_t (new_AGEMA_signal_5244), .A1_f (new_AGEMA_signal_5245), .B0_t (Midori_rounds_mul_MC3_n5), .B0_f (new_AGEMA_signal_5437), .B1_t (new_AGEMA_signal_5438), .B1_f (new_AGEMA_signal_5439), .Z0_t (Midori_rounds_SR_Inv_Result[15]), .Z0_f (new_AGEMA_signal_5553), .Z1_t (new_AGEMA_signal_5554), .Z1_f (new_AGEMA_signal_5555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U14 ( .A0_t (Midori_rounds_mul_input[23]), .A0_f (new_AGEMA_signal_5252), .A1_t (new_AGEMA_signal_5253), .A1_f (new_AGEMA_signal_5254), .B0_t (Midori_rounds_mul_MC3_n5), .B0_f (new_AGEMA_signal_5437), .B1_t (new_AGEMA_signal_5438), .B1_f (new_AGEMA_signal_5439), .Z0_t (Midori_rounds_SR_Inv_Result[39]), .Z0_f (new_AGEMA_signal_5556), .Z1_t (new_AGEMA_signal_5557), .Z1_f (new_AGEMA_signal_5558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U13 ( .A0_t (Midori_rounds_mul_input[27]), .A0_f (new_AGEMA_signal_5261), .A1_t (new_AGEMA_signal_5262), .A1_f (new_AGEMA_signal_5263), .B0_t (Midori_rounds_mul_input[31]), .B0_f (new_AGEMA_signal_5270), .B1_t (new_AGEMA_signal_5271), .B1_f (new_AGEMA_signal_5272), .Z0_t (Midori_rounds_mul_MC3_n5), .Z0_f (new_AGEMA_signal_5437), .Z1_t (new_AGEMA_signal_5438), .Z1_f (new_AGEMA_signal_5439) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U12 ( .A0_t (Midori_rounds_mul_input[25]), .A0_f (new_AGEMA_signal_5255), .A1_t (new_AGEMA_signal_5256), .A1_f (new_AGEMA_signal_5257), .B0_t (Midori_rounds_mul_MC3_n4), .B0_f (new_AGEMA_signal_5440), .B1_t (new_AGEMA_signal_5441), .B1_f (new_AGEMA_signal_5442), .Z0_t (Midori_rounds_SR_Inv_Result[25]), .Z0_f (new_AGEMA_signal_5559), .Z1_t (new_AGEMA_signal_5560), .Z1_f (new_AGEMA_signal_5561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U11 ( .A0_t (Midori_rounds_mul_input[29]), .A0_f (new_AGEMA_signal_5264), .A1_t (new_AGEMA_signal_5265), .A1_f (new_AGEMA_signal_5266), .B0_t (Midori_rounds_mul_MC3_n4), .B0_f (new_AGEMA_signal_5440), .B1_t (new_AGEMA_signal_5441), .B1_f (new_AGEMA_signal_5442), .Z0_t (Midori_rounds_SR_Inv_Result[49]), .Z0_f (new_AGEMA_signal_5562), .Z1_t (new_AGEMA_signal_5563), .Z1_f (new_AGEMA_signal_5564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U10 ( .A0_t (Midori_rounds_mul_input[21]), .A0_f (new_AGEMA_signal_5246), .A1_t (new_AGEMA_signal_5247), .A1_f (new_AGEMA_signal_5248), .B0_t (Midori_rounds_mul_input[17]), .B0_f (new_AGEMA_signal_5237), .B1_t (new_AGEMA_signal_5238), .B1_f (new_AGEMA_signal_5239), .Z0_t (Midori_rounds_mul_MC3_n4), .Z0_f (new_AGEMA_signal_5440), .Z1_t (new_AGEMA_signal_5441), .Z1_f (new_AGEMA_signal_5442) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U9 ( .A0_t (Midori_rounds_mul_input[18]), .A0_f (new_AGEMA_signal_5374), .A1_t (new_AGEMA_signal_5375), .A1_f (new_AGEMA_signal_5376), .B0_t (Midori_rounds_mul_MC3_n3), .B0_f (new_AGEMA_signal_5565), .B1_t (new_AGEMA_signal_5566), .B1_f (new_AGEMA_signal_5567), .Z0_t (Midori_rounds_SR_Inv_Result[14]), .Z0_f (new_AGEMA_signal_5770), .Z1_t (new_AGEMA_signal_5771), .Z1_f (new_AGEMA_signal_5772) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U8 ( .A0_t (Midori_rounds_mul_input[22]), .A0_f (new_AGEMA_signal_5377), .A1_t (new_AGEMA_signal_5378), .A1_f (new_AGEMA_signal_5379), .B0_t (Midori_rounds_mul_MC3_n3), .B0_f (new_AGEMA_signal_5565), .B1_t (new_AGEMA_signal_5566), .B1_f (new_AGEMA_signal_5567), .Z0_t (Midori_rounds_SR_Inv_Result[38]), .Z0_f (new_AGEMA_signal_5773), .Z1_t (new_AGEMA_signal_5774), .Z1_f (new_AGEMA_signal_5775) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U7 ( .A0_t (Midori_rounds_mul_input[26]), .A0_f (new_AGEMA_signal_5380), .A1_t (new_AGEMA_signal_5381), .A1_f (new_AGEMA_signal_5382), .B0_t (Midori_rounds_mul_input[30]), .B0_f (new_AGEMA_signal_5383), .B1_t (new_AGEMA_signal_5384), .B1_f (new_AGEMA_signal_5385), .Z0_t (Midori_rounds_mul_MC3_n3), .Z0_f (new_AGEMA_signal_5565), .Z1_t (new_AGEMA_signal_5566), .Z1_f (new_AGEMA_signal_5567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U6 ( .A0_t (Midori_rounds_mul_input[17]), .A0_f (new_AGEMA_signal_5237), .A1_t (new_AGEMA_signal_5238), .A1_f (new_AGEMA_signal_5239), .B0_t (Midori_rounds_mul_MC3_n2), .B0_f (new_AGEMA_signal_5443), .B1_t (new_AGEMA_signal_5444), .B1_f (new_AGEMA_signal_5445), .Z0_t (Midori_rounds_SR_Inv_Result[13]), .Z0_f (new_AGEMA_signal_5568), .Z1_t (new_AGEMA_signal_5569), .Z1_f (new_AGEMA_signal_5570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U5 ( .A0_t (Midori_rounds_mul_input[21]), .A0_f (new_AGEMA_signal_5246), .A1_t (new_AGEMA_signal_5247), .A1_f (new_AGEMA_signal_5248), .B0_t (Midori_rounds_mul_MC3_n2), .B0_f (new_AGEMA_signal_5443), .B1_t (new_AGEMA_signal_5444), .B1_f (new_AGEMA_signal_5445), .Z0_t (Midori_rounds_SR_Inv_Result[37]), .Z0_f (new_AGEMA_signal_5571), .Z1_t (new_AGEMA_signal_5572), .Z1_f (new_AGEMA_signal_5573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U4 ( .A0_t (Midori_rounds_mul_input[25]), .A0_f (new_AGEMA_signal_5255), .A1_t (new_AGEMA_signal_5256), .A1_f (new_AGEMA_signal_5257), .B0_t (Midori_rounds_mul_input[29]), .B0_f (new_AGEMA_signal_5264), .B1_t (new_AGEMA_signal_5265), .B1_f (new_AGEMA_signal_5266), .Z0_t (Midori_rounds_mul_MC3_n2), .Z0_f (new_AGEMA_signal_5443), .Z1_t (new_AGEMA_signal_5444), .Z1_f (new_AGEMA_signal_5445) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U3 ( .A0_t (Midori_rounds_mul_input[16]), .A0_f (new_AGEMA_signal_6680), .A1_t (new_AGEMA_signal_6681), .A1_f (new_AGEMA_signal_6682), .B0_t (Midori_rounds_mul_MC3_n1), .B0_f (new_AGEMA_signal_6695), .B1_t (new_AGEMA_signal_6696), .B1_f (new_AGEMA_signal_6697), .Z0_t (Midori_rounds_SR_Inv_Result[12]), .Z0_f (new_AGEMA_signal_6773), .Z1_t (new_AGEMA_signal_6774), .Z1_f (new_AGEMA_signal_6775) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U2 ( .A0_t (Midori_rounds_mul_input[20]), .A0_f (new_AGEMA_signal_6182), .A1_t (new_AGEMA_signal_6183), .A1_f (new_AGEMA_signal_6184), .B0_t (Midori_rounds_mul_MC3_n1), .B0_f (new_AGEMA_signal_6695), .B1_t (new_AGEMA_signal_6696), .B1_f (new_AGEMA_signal_6697), .Z0_t (Midori_rounds_SR_Inv_Result[36]), .Z0_f (new_AGEMA_signal_6776), .Z1_t (new_AGEMA_signal_6777), .Z1_f (new_AGEMA_signal_6778) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U1 ( .A0_t (Midori_rounds_mul_input[24]), .A0_f (new_AGEMA_signal_6002), .A1_t (new_AGEMA_signal_6003), .A1_f (new_AGEMA_signal_6004), .B0_t (Midori_rounds_mul_input[28]), .B0_f (new_AGEMA_signal_6464), .B1_t (new_AGEMA_signal_6465), .B1_f (new_AGEMA_signal_6466), .Z0_t (Midori_rounds_mul_MC3_n1), .Z0_f (new_AGEMA_signal_6695), .Z1_t (new_AGEMA_signal_6696), .Z1_f (new_AGEMA_signal_6697) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U24 ( .A0_t (Midori_rounds_mul_input[11]), .A0_f (new_AGEMA_signal_5225), .A1_t (new_AGEMA_signal_5226), .A1_f (new_AGEMA_signal_5227), .B0_t (Midori_rounds_mul_MC4_n8), .B0_f (new_AGEMA_signal_5446), .B1_t (new_AGEMA_signal_5447), .B1_f (new_AGEMA_signal_5448), .Z0_t (Midori_rounds_SR_Inv_Result[35]), .Z0_f (new_AGEMA_signal_5574), .Z1_t (new_AGEMA_signal_5575), .Z1_f (new_AGEMA_signal_5576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U23 ( .A0_t (Midori_rounds_mul_input[15]), .A0_f (new_AGEMA_signal_5234), .A1_t (new_AGEMA_signal_5235), .A1_f (new_AGEMA_signal_5236), .B0_t (Midori_rounds_mul_MC4_n8), .B0_f (new_AGEMA_signal_5446), .B1_t (new_AGEMA_signal_5447), .B1_f (new_AGEMA_signal_5448), .Z0_t (Midori_rounds_SR_Inv_Result[11]), .Z0_f (new_AGEMA_signal_5577), .Z1_t (new_AGEMA_signal_5578), .Z1_f (new_AGEMA_signal_5579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U22 ( .A0_t (Midori_rounds_mul_input[7]), .A0_f (new_AGEMA_signal_5216), .A1_t (new_AGEMA_signal_5217), .A1_f (new_AGEMA_signal_5218), .B0_t (Midori_rounds_mul_input[3]), .B0_f (new_AGEMA_signal_5207), .B1_t (new_AGEMA_signal_5208), .B1_f (new_AGEMA_signal_5209), .Z0_t (Midori_rounds_mul_MC4_n8), .Z0_f (new_AGEMA_signal_5446), .Z1_t (new_AGEMA_signal_5447), .Z1_f (new_AGEMA_signal_5448) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U21 ( .A0_t (Midori_rounds_mul_input[10]), .A0_f (new_AGEMA_signal_5368), .A1_t (new_AGEMA_signal_5369), .A1_f (new_AGEMA_signal_5370), .B0_t (Midori_rounds_mul_MC4_n7), .B0_f (new_AGEMA_signal_5580), .B1_t (new_AGEMA_signal_5581), .B1_f (new_AGEMA_signal_5582), .Z0_t (Midori_rounds_SR_Inv_Result[34]), .Z0_f (new_AGEMA_signal_5776), .Z1_t (new_AGEMA_signal_5777), .Z1_f (new_AGEMA_signal_5778) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U20 ( .A0_t (Midori_rounds_mul_input[14]), .A0_f (new_AGEMA_signal_5371), .A1_t (new_AGEMA_signal_5372), .A1_f (new_AGEMA_signal_5373), .B0_t (Midori_rounds_mul_MC4_n7), .B0_f (new_AGEMA_signal_5580), .B1_t (new_AGEMA_signal_5581), .B1_f (new_AGEMA_signal_5582), .Z0_t (Midori_rounds_SR_Inv_Result[10]), .Z0_f (new_AGEMA_signal_5779), .Z1_t (new_AGEMA_signal_5780), .Z1_f (new_AGEMA_signal_5781) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U19 ( .A0_t (Midori_rounds_mul_input[6]), .A0_f (new_AGEMA_signal_5365), .A1_t (new_AGEMA_signal_5366), .A1_f (new_AGEMA_signal_5367), .B0_t (Midori_rounds_mul_input[2]), .B0_f (new_AGEMA_signal_5362), .B1_t (new_AGEMA_signal_5363), .B1_f (new_AGEMA_signal_5364), .Z0_t (Midori_rounds_mul_MC4_n7), .Z0_f (new_AGEMA_signal_5580), .Z1_t (new_AGEMA_signal_5581), .Z1_f (new_AGEMA_signal_5582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U18 ( .A0_t (Midori_rounds_mul_input[8]), .A0_f (new_AGEMA_signal_6455), .A1_t (new_AGEMA_signal_6456), .A1_f (new_AGEMA_signal_6457), .B0_t (Midori_rounds_mul_MC4_n6), .B0_f (new_AGEMA_signal_6815), .B1_t (new_AGEMA_signal_6816), .B1_f (new_AGEMA_signal_6817), .Z0_t (Midori_rounds_SR_Inv_Result[32]), .Z0_f (new_AGEMA_signal_6842), .Z1_t (new_AGEMA_signal_6843), .Z1_f (new_AGEMA_signal_6844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U17 ( .A0_t (Midori_rounds_mul_input[12]), .A0_f (new_AGEMA_signal_6458), .A1_t (new_AGEMA_signal_6459), .A1_f (new_AGEMA_signal_6460), .B0_t (Midori_rounds_mul_MC4_n6), .B0_f (new_AGEMA_signal_6815), .B1_t (new_AGEMA_signal_6816), .B1_f (new_AGEMA_signal_6817), .Z0_t (Midori_rounds_SR_Inv_Result[8]), .Z0_f (new_AGEMA_signal_6845), .Z1_t (new_AGEMA_signal_6846), .Z1_f (new_AGEMA_signal_6847) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U16 ( .A0_t (Midori_rounds_mul_input[4]), .A0_f (new_AGEMA_signal_6755), .A1_t (new_AGEMA_signal_6756), .A1_f (new_AGEMA_signal_6757), .B0_t (Midori_rounds_mul_input[0]), .B0_f (new_AGEMA_signal_6449), .B1_t (new_AGEMA_signal_6450), .B1_f (new_AGEMA_signal_6451), .Z0_t (Midori_rounds_mul_MC4_n6), .Z0_f (new_AGEMA_signal_6815), .Z1_t (new_AGEMA_signal_6816), .Z1_f (new_AGEMA_signal_6817) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U15 ( .A0_t (Midori_rounds_mul_input[3]), .A0_f (new_AGEMA_signal_5207), .A1_t (new_AGEMA_signal_5208), .A1_f (new_AGEMA_signal_5209), .B0_t (Midori_rounds_mul_MC4_n5), .B0_f (new_AGEMA_signal_5449), .B1_t (new_AGEMA_signal_5450), .B1_f (new_AGEMA_signal_5451), .Z0_t (Midori_rounds_SR_Inv_Result[55]), .Z0_f (new_AGEMA_signal_5583), .Z1_t (new_AGEMA_signal_5584), .Z1_f (new_AGEMA_signal_5585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U14 ( .A0_t (Midori_rounds_mul_input[7]), .A0_f (new_AGEMA_signal_5216), .A1_t (new_AGEMA_signal_5217), .A1_f (new_AGEMA_signal_5218), .B0_t (Midori_rounds_mul_MC4_n5), .B0_f (new_AGEMA_signal_5449), .B1_t (new_AGEMA_signal_5450), .B1_f (new_AGEMA_signal_5451), .Z0_t (Midori_rounds_SR_Inv_Result[31]), .Z0_f (new_AGEMA_signal_5586), .Z1_t (new_AGEMA_signal_5587), .Z1_f (new_AGEMA_signal_5588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U13 ( .A0_t (Midori_rounds_mul_input[11]), .A0_f (new_AGEMA_signal_5225), .A1_t (new_AGEMA_signal_5226), .A1_f (new_AGEMA_signal_5227), .B0_t (Midori_rounds_mul_input[15]), .B0_f (new_AGEMA_signal_5234), .B1_t (new_AGEMA_signal_5235), .B1_f (new_AGEMA_signal_5236), .Z0_t (Midori_rounds_mul_MC4_n5), .Z0_f (new_AGEMA_signal_5449), .Z1_t (new_AGEMA_signal_5450), .Z1_f (new_AGEMA_signal_5451) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U12 ( .A0_t (Midori_rounds_mul_input[9]), .A0_f (new_AGEMA_signal_5219), .A1_t (new_AGEMA_signal_5220), .A1_f (new_AGEMA_signal_5221), .B0_t (Midori_rounds_mul_MC4_n4), .B0_f (new_AGEMA_signal_5452), .B1_t (new_AGEMA_signal_5453), .B1_f (new_AGEMA_signal_5454), .Z0_t (Midori_rounds_SR_Inv_Result[33]), .Z0_f (new_AGEMA_signal_5589), .Z1_t (new_AGEMA_signal_5590), .Z1_f (new_AGEMA_signal_5591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U11 ( .A0_t (Midori_rounds_mul_input[13]), .A0_f (new_AGEMA_signal_5228), .A1_t (new_AGEMA_signal_5229), .A1_f (new_AGEMA_signal_5230), .B0_t (Midori_rounds_mul_MC4_n4), .B0_f (new_AGEMA_signal_5452), .B1_t (new_AGEMA_signal_5453), .B1_f (new_AGEMA_signal_5454), .Z0_t (Midori_rounds_SR_Inv_Result[9]), .Z0_f (new_AGEMA_signal_5592), .Z1_t (new_AGEMA_signal_5593), .Z1_f (new_AGEMA_signal_5594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U10 ( .A0_t (Midori_rounds_mul_input[5]), .A0_f (new_AGEMA_signal_5210), .A1_t (new_AGEMA_signal_5211), .A1_f (new_AGEMA_signal_5212), .B0_t (Midori_rounds_mul_input[1]), .B0_f (new_AGEMA_signal_5201), .B1_t (new_AGEMA_signal_5202), .B1_f (new_AGEMA_signal_5203), .Z0_t (Midori_rounds_mul_MC4_n4), .Z0_f (new_AGEMA_signal_5452), .Z1_t (new_AGEMA_signal_5453), .Z1_f (new_AGEMA_signal_5454) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U9 ( .A0_t (Midori_rounds_mul_input[2]), .A0_f (new_AGEMA_signal_5362), .A1_t (new_AGEMA_signal_5363), .A1_f (new_AGEMA_signal_5364), .B0_t (Midori_rounds_mul_MC4_n3), .B0_f (new_AGEMA_signal_5595), .B1_t (new_AGEMA_signal_5596), .B1_f (new_AGEMA_signal_5597), .Z0_t (Midori_rounds_SR_Inv_Result[54]), .Z0_f (new_AGEMA_signal_5782), .Z1_t (new_AGEMA_signal_5783), .Z1_f (new_AGEMA_signal_5784) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U8 ( .A0_t (Midori_rounds_mul_input[6]), .A0_f (new_AGEMA_signal_5365), .A1_t (new_AGEMA_signal_5366), .A1_f (new_AGEMA_signal_5367), .B0_t (Midori_rounds_mul_MC4_n3), .B0_f (new_AGEMA_signal_5595), .B1_t (new_AGEMA_signal_5596), .B1_f (new_AGEMA_signal_5597), .Z0_t (Midori_rounds_SR_Inv_Result[30]), .Z0_f (new_AGEMA_signal_5785), .Z1_t (new_AGEMA_signal_5786), .Z1_f (new_AGEMA_signal_5787) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U7 ( .A0_t (Midori_rounds_mul_input[10]), .A0_f (new_AGEMA_signal_5368), .A1_t (new_AGEMA_signal_5369), .A1_f (new_AGEMA_signal_5370), .B0_t (Midori_rounds_mul_input[14]), .B0_f (new_AGEMA_signal_5371), .B1_t (new_AGEMA_signal_5372), .B1_f (new_AGEMA_signal_5373), .Z0_t (Midori_rounds_mul_MC4_n3), .Z0_f (new_AGEMA_signal_5595), .Z1_t (new_AGEMA_signal_5596), .Z1_f (new_AGEMA_signal_5597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U6 ( .A0_t (Midori_rounds_mul_input[1]), .A0_f (new_AGEMA_signal_5201), .A1_t (new_AGEMA_signal_5202), .A1_f (new_AGEMA_signal_5203), .B0_t (Midori_rounds_mul_MC4_n2), .B0_f (new_AGEMA_signal_5455), .B1_t (new_AGEMA_signal_5456), .B1_f (new_AGEMA_signal_5457), .Z0_t (Midori_rounds_SR_Inv_Result[53]), .Z0_f (new_AGEMA_signal_5598), .Z1_t (new_AGEMA_signal_5599), .Z1_f (new_AGEMA_signal_5600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U5 ( .A0_t (Midori_rounds_mul_input[5]), .A0_f (new_AGEMA_signal_5210), .A1_t (new_AGEMA_signal_5211), .A1_f (new_AGEMA_signal_5212), .B0_t (Midori_rounds_mul_MC4_n2), .B0_f (new_AGEMA_signal_5455), .B1_t (new_AGEMA_signal_5456), .B1_f (new_AGEMA_signal_5457), .Z0_t (Midori_rounds_SR_Inv_Result[29]), .Z0_f (new_AGEMA_signal_5601), .Z1_t (new_AGEMA_signal_5602), .Z1_f (new_AGEMA_signal_5603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U4 ( .A0_t (Midori_rounds_mul_input[9]), .A0_f (new_AGEMA_signal_5219), .A1_t (new_AGEMA_signal_5220), .A1_f (new_AGEMA_signal_5221), .B0_t (Midori_rounds_mul_input[13]), .B0_f (new_AGEMA_signal_5228), .B1_t (new_AGEMA_signal_5229), .B1_f (new_AGEMA_signal_5230), .Z0_t (Midori_rounds_mul_MC4_n2), .Z0_f (new_AGEMA_signal_5455), .Z1_t (new_AGEMA_signal_5456), .Z1_f (new_AGEMA_signal_5457) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U3 ( .A0_t (Midori_rounds_mul_input[0]), .A0_f (new_AGEMA_signal_6449), .A1_t (new_AGEMA_signal_6450), .A1_f (new_AGEMA_signal_6451), .B0_t (Midori_rounds_mul_MC4_n1), .B0_f (new_AGEMA_signal_6698), .B1_t (new_AGEMA_signal_6699), .B1_f (new_AGEMA_signal_6700), .Z0_t (Midori_rounds_SR_Inv_Result[52]), .Z0_f (new_AGEMA_signal_6779), .Z1_t (new_AGEMA_signal_6780), .Z1_f (new_AGEMA_signal_6781) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U2 ( .A0_t (Midori_rounds_mul_input[4]), .A0_f (new_AGEMA_signal_6755), .A1_t (new_AGEMA_signal_6756), .A1_f (new_AGEMA_signal_6757), .B0_t (Midori_rounds_mul_MC4_n1), .B0_f (new_AGEMA_signal_6698), .B1_t (new_AGEMA_signal_6699), .B1_f (new_AGEMA_signal_6700), .Z0_t (Midori_rounds_SR_Inv_Result[28]), .Z0_f (new_AGEMA_signal_6818), .Z1_t (new_AGEMA_signal_6819), .Z1_f (new_AGEMA_signal_6820) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U1 ( .A0_t (Midori_rounds_mul_input[8]), .A0_f (new_AGEMA_signal_6455), .A1_t (new_AGEMA_signal_6456), .A1_f (new_AGEMA_signal_6457), .B0_t (Midori_rounds_mul_input[12]), .B0_f (new_AGEMA_signal_6458), .B1_t (new_AGEMA_signal_6459), .B1_f (new_AGEMA_signal_6460), .Z0_t (Midori_rounds_mul_MC4_n1), .Z0_f (new_AGEMA_signal_6698), .Z1_t (new_AGEMA_signal_6699), .Z1_f (new_AGEMA_signal_6700) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_0_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[0]), .A0_f (new_AGEMA_signal_6836), .A1_t (new_AGEMA_signal_6837), .A1_f (new_AGEMA_signal_6838), .B0_t (Midori_rounds_SR_Inv_Result[0]), .B0_f (new_AGEMA_signal_6689), .B1_t (new_AGEMA_signal_6690), .B1_f (new_AGEMA_signal_6691), .Z0_t (Midori_rounds_Res_Inst_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_6872), .Z1_t (new_AGEMA_signal_6873), .Z1_f (new_AGEMA_signal_6874) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_6872), .B1_t (new_AGEMA_signal_6873), .B1_f (new_AGEMA_signal_6874), .Z0_t (Midori_rounds_Res_Inst_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_6914), .Z1_t (new_AGEMA_signal_6915), .Z1_f (new_AGEMA_signal_6916) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_0_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_6914), .A1_t (new_AGEMA_signal_6915), .A1_f (new_AGEMA_signal_6916), .B0_t (Midori_rounds_mul_ResultXORkey[0]), .B0_f (new_AGEMA_signal_6836), .B1_t (new_AGEMA_signal_6837), .B1_f (new_AGEMA_signal_6838), .Z0_t (Midori_rounds_round_Result[0]), .Z0_f (new_AGEMA_signal_6980), .Z1_t (new_AGEMA_signal_6981), .Z1_f (new_AGEMA_signal_6982) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_1_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[1]), .A0_f (new_AGEMA_signal_5727), .A1_t (new_AGEMA_signal_5728), .A1_f (new_AGEMA_signal_5729), .B0_t (Midori_rounds_SR_Inv_Result[1]), .B0_f (new_AGEMA_signal_5511), .B1_t (new_AGEMA_signal_5512), .B1_f (new_AGEMA_signal_5513), .Z0_t (Midori_rounds_Res_Inst_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_5882), .Z1_t (new_AGEMA_signal_5883), .Z1_f (new_AGEMA_signal_5884) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_5882), .B1_t (new_AGEMA_signal_5883), .B1_f (new_AGEMA_signal_5884), .Z0_t (Midori_rounds_Res_Inst_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_6023), .Z1_t (new_AGEMA_signal_6024), .Z1_f (new_AGEMA_signal_6025) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_1_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_6023), .A1_t (new_AGEMA_signal_6024), .A1_f (new_AGEMA_signal_6025), .B0_t (Midori_rounds_mul_ResultXORkey[1]), .B0_f (new_AGEMA_signal_5727), .B1_t (new_AGEMA_signal_5728), .B1_f (new_AGEMA_signal_5729), .Z0_t (Midori_rounds_round_Result[1]), .Z0_f (new_AGEMA_signal_6209), .Z1_t (new_AGEMA_signal_6210), .Z1_f (new_AGEMA_signal_6211) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_2_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[2]), .A0_f (new_AGEMA_signal_5860), .A1_t (new_AGEMA_signal_5861), .A1_f (new_AGEMA_signal_5862), .B0_t (Midori_rounds_SR_Inv_Result[2]), .B0_f (new_AGEMA_signal_5749), .B1_t (new_AGEMA_signal_5750), .B1_f (new_AGEMA_signal_5751), .Z0_t (Midori_rounds_Res_Inst_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_6026), .Z1_t (new_AGEMA_signal_6027), .Z1_f (new_AGEMA_signal_6028) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_6026), .B1_t (new_AGEMA_signal_6027), .B1_f (new_AGEMA_signal_6028), .Z0_t (Midori_rounds_Res_Inst_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_6212), .Z1_t (new_AGEMA_signal_6213), .Z1_f (new_AGEMA_signal_6214) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_2_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_6212), .A1_t (new_AGEMA_signal_6213), .A1_f (new_AGEMA_signal_6214), .B0_t (Midori_rounds_mul_ResultXORkey[2]), .B0_f (new_AGEMA_signal_5860), .B1_t (new_AGEMA_signal_5861), .B1_f (new_AGEMA_signal_5862), .Z0_t (Midori_rounds_round_Result[2]), .Z0_f (new_AGEMA_signal_6485), .Z1_t (new_AGEMA_signal_6486), .Z1_f (new_AGEMA_signal_6487) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_3_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[3]), .A0_f (new_AGEMA_signal_5724), .A1_t (new_AGEMA_signal_5725), .A1_f (new_AGEMA_signal_5726), .B0_t (Midori_rounds_SR_Inv_Result[3]), .B0_f (new_AGEMA_signal_5496), .B1_t (new_AGEMA_signal_5497), .B1_f (new_AGEMA_signal_5498), .Z0_t (Midori_rounds_Res_Inst_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_5885), .Z1_t (new_AGEMA_signal_5886), .Z1_f (new_AGEMA_signal_5887) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_5885), .B1_t (new_AGEMA_signal_5886), .B1_f (new_AGEMA_signal_5887), .Z0_t (Midori_rounds_Res_Inst_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_6029), .Z1_t (new_AGEMA_signal_6030), .Z1_f (new_AGEMA_signal_6031) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_3_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_6029), .A1_t (new_AGEMA_signal_6030), .A1_f (new_AGEMA_signal_6031), .B0_t (Midori_rounds_mul_ResultXORkey[3]), .B0_f (new_AGEMA_signal_5724), .B1_t (new_AGEMA_signal_5725), .B1_f (new_AGEMA_signal_5726), .Z0_t (Midori_rounds_round_Result[3]), .Z0_f (new_AGEMA_signal_6215), .Z1_t (new_AGEMA_signal_6216), .Z1_f (new_AGEMA_signal_6217) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_4_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[4]), .A0_f (new_AGEMA_signal_6782), .A1_t (new_AGEMA_signal_6783), .A1_f (new_AGEMA_signal_6784), .B0_t (Midori_rounds_SR_Inv_Result[4]), .B0_f (new_AGEMA_signal_6803), .B1_t (new_AGEMA_signal_6804), .B1_f (new_AGEMA_signal_6805), .Z0_t (Midori_rounds_Res_Inst_mux_inst_4_U1_X), .Z0_f (new_AGEMA_signal_6848), .Z1_t (new_AGEMA_signal_6849), .Z1_f (new_AGEMA_signal_6850) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_4_U1_X), .B0_f (new_AGEMA_signal_6848), .B1_t (new_AGEMA_signal_6849), .B1_f (new_AGEMA_signal_6850), .Z0_t (Midori_rounds_Res_Inst_mux_inst_4_U1_Y), .Z0_f (new_AGEMA_signal_6875), .Z1_t (new_AGEMA_signal_6876), .Z1_f (new_AGEMA_signal_6877) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_4_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_4_U1_Y), .A0_f (new_AGEMA_signal_6875), .A1_t (new_AGEMA_signal_6876), .A1_f (new_AGEMA_signal_6877), .B0_t (Midori_rounds_mul_ResultXORkey[4]), .B0_f (new_AGEMA_signal_6782), .B1_t (new_AGEMA_signal_6783), .B1_f (new_AGEMA_signal_6784), .Z0_t (Midori_rounds_round_Result[4]), .Z0_f (new_AGEMA_signal_6917), .Z1_t (new_AGEMA_signal_6918), .Z1_f (new_AGEMA_signal_6919) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_5_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[5]), .A0_f (new_AGEMA_signal_5721), .A1_t (new_AGEMA_signal_5722), .A1_f (new_AGEMA_signal_5723), .B0_t (Midori_rounds_SR_Inv_Result[5]), .B0_f (new_AGEMA_signal_5529), .B1_t (new_AGEMA_signal_5530), .B1_f (new_AGEMA_signal_5531), .Z0_t (Midori_rounds_Res_Inst_mux_inst_5_U1_X), .Z0_f (new_AGEMA_signal_5888), .Z1_t (new_AGEMA_signal_5889), .Z1_f (new_AGEMA_signal_5890) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_5_U1_X), .B0_f (new_AGEMA_signal_5888), .B1_t (new_AGEMA_signal_5889), .B1_f (new_AGEMA_signal_5890), .Z0_t (Midori_rounds_Res_Inst_mux_inst_5_U1_Y), .Z0_f (new_AGEMA_signal_6032), .Z1_t (new_AGEMA_signal_6033), .Z1_f (new_AGEMA_signal_6034) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_5_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_5_U1_Y), .A0_f (new_AGEMA_signal_6032), .A1_t (new_AGEMA_signal_6033), .A1_f (new_AGEMA_signal_6034), .B0_t (Midori_rounds_mul_ResultXORkey[5]), .B0_f (new_AGEMA_signal_5721), .B1_t (new_AGEMA_signal_5722), .B1_f (new_AGEMA_signal_5723), .Z0_t (Midori_rounds_round_Result[5]), .Z0_f (new_AGEMA_signal_6218), .Z1_t (new_AGEMA_signal_6219), .Z1_f (new_AGEMA_signal_6220) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_6_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[6]), .A0_f (new_AGEMA_signal_5857), .A1_t (new_AGEMA_signal_5858), .A1_f (new_AGEMA_signal_5859), .B0_t (Midori_rounds_SR_Inv_Result[6]), .B0_f (new_AGEMA_signal_5752), .B1_t (new_AGEMA_signal_5753), .B1_f (new_AGEMA_signal_5754), .Z0_t (Midori_rounds_Res_Inst_mux_inst_6_U1_X), .Z0_f (new_AGEMA_signal_6035), .Z1_t (new_AGEMA_signal_6036), .Z1_f (new_AGEMA_signal_6037) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_6_U1_X), .B0_f (new_AGEMA_signal_6035), .B1_t (new_AGEMA_signal_6036), .B1_f (new_AGEMA_signal_6037), .Z0_t (Midori_rounds_Res_Inst_mux_inst_6_U1_Y), .Z0_f (new_AGEMA_signal_6221), .Z1_t (new_AGEMA_signal_6222), .Z1_f (new_AGEMA_signal_6223) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_6_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_6_U1_Y), .A0_f (new_AGEMA_signal_6221), .A1_t (new_AGEMA_signal_6222), .A1_f (new_AGEMA_signal_6223), .B0_t (Midori_rounds_mul_ResultXORkey[6]), .B0_f (new_AGEMA_signal_5857), .B1_t (new_AGEMA_signal_5858), .B1_f (new_AGEMA_signal_5859), .Z0_t (Midori_rounds_round_Result[6]), .Z0_f (new_AGEMA_signal_6488), .Z1_t (new_AGEMA_signal_6489), .Z1_f (new_AGEMA_signal_6490) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_7_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[7]), .A0_f (new_AGEMA_signal_5718), .A1_t (new_AGEMA_signal_5719), .A1_f (new_AGEMA_signal_5720), .B0_t (Midori_rounds_SR_Inv_Result[7]), .B0_f (new_AGEMA_signal_5514), .B1_t (new_AGEMA_signal_5515), .B1_f (new_AGEMA_signal_5516), .Z0_t (Midori_rounds_Res_Inst_mux_inst_7_U1_X), .Z0_f (new_AGEMA_signal_5891), .Z1_t (new_AGEMA_signal_5892), .Z1_f (new_AGEMA_signal_5893) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_7_U1_X), .B0_f (new_AGEMA_signal_5891), .B1_t (new_AGEMA_signal_5892), .B1_f (new_AGEMA_signal_5893), .Z0_t (Midori_rounds_Res_Inst_mux_inst_7_U1_Y), .Z0_f (new_AGEMA_signal_6038), .Z1_t (new_AGEMA_signal_6039), .Z1_f (new_AGEMA_signal_6040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_7_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_7_U1_Y), .A0_f (new_AGEMA_signal_6038), .A1_t (new_AGEMA_signal_6039), .A1_f (new_AGEMA_signal_6040), .B0_t (Midori_rounds_mul_ResultXORkey[7]), .B0_f (new_AGEMA_signal_5718), .B1_t (new_AGEMA_signal_5719), .B1_f (new_AGEMA_signal_5720), .Z0_t (Midori_rounds_round_Result[7]), .Z0_f (new_AGEMA_signal_6224), .Z1_t (new_AGEMA_signal_6225), .Z1_f (new_AGEMA_signal_6226) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_8_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[8]), .A0_f (new_AGEMA_signal_6869), .A1_t (new_AGEMA_signal_6870), .A1_f (new_AGEMA_signal_6871), .B0_t (Midori_rounds_SR_Inv_Result[8]), .B0_f (new_AGEMA_signal_6845), .B1_t (new_AGEMA_signal_6846), .B1_f (new_AGEMA_signal_6847), .Z0_t (Midori_rounds_Res_Inst_mux_inst_8_U1_X), .Z0_f (new_AGEMA_signal_6920), .Z1_t (new_AGEMA_signal_6921), .Z1_f (new_AGEMA_signal_6922) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_8_U1_X), .B0_f (new_AGEMA_signal_6920), .B1_t (new_AGEMA_signal_6921), .B1_f (new_AGEMA_signal_6922), .Z0_t (Midori_rounds_Res_Inst_mux_inst_8_U1_Y), .Z0_f (new_AGEMA_signal_6983), .Z1_t (new_AGEMA_signal_6984), .Z1_f (new_AGEMA_signal_6985) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_8_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_8_U1_Y), .A0_f (new_AGEMA_signal_6983), .A1_t (new_AGEMA_signal_6984), .A1_f (new_AGEMA_signal_6985), .B0_t (Midori_rounds_mul_ResultXORkey[8]), .B0_f (new_AGEMA_signal_6869), .B1_t (new_AGEMA_signal_6870), .B1_f (new_AGEMA_signal_6871), .Z0_t (Midori_rounds_round_Result[8]), .Z0_f (new_AGEMA_signal_7052), .Z1_t (new_AGEMA_signal_7053), .Z1_f (new_AGEMA_signal_7054) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_9_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[9]), .A0_f (new_AGEMA_signal_5715), .A1_t (new_AGEMA_signal_5716), .A1_f (new_AGEMA_signal_5717), .B0_t (Midori_rounds_SR_Inv_Result[9]), .B0_f (new_AGEMA_signal_5592), .B1_t (new_AGEMA_signal_5593), .B1_f (new_AGEMA_signal_5594), .Z0_t (Midori_rounds_Res_Inst_mux_inst_9_U1_X), .Z0_f (new_AGEMA_signal_5894), .Z1_t (new_AGEMA_signal_5895), .Z1_f (new_AGEMA_signal_5896) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_9_U1_X), .B0_f (new_AGEMA_signal_5894), .B1_t (new_AGEMA_signal_5895), .B1_f (new_AGEMA_signal_5896), .Z0_t (Midori_rounds_Res_Inst_mux_inst_9_U1_Y), .Z0_f (new_AGEMA_signal_6041), .Z1_t (new_AGEMA_signal_6042), .Z1_f (new_AGEMA_signal_6043) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_9_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_9_U1_Y), .A0_f (new_AGEMA_signal_6041), .A1_t (new_AGEMA_signal_6042), .A1_f (new_AGEMA_signal_6043), .B0_t (Midori_rounds_mul_ResultXORkey[9]), .B0_f (new_AGEMA_signal_5715), .B1_t (new_AGEMA_signal_5716), .B1_f (new_AGEMA_signal_5717), .Z0_t (Midori_rounds_round_Result[9]), .Z0_f (new_AGEMA_signal_6227), .Z1_t (new_AGEMA_signal_6228), .Z1_f (new_AGEMA_signal_6229) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_10_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[10]), .A0_f (new_AGEMA_signal_5854), .A1_t (new_AGEMA_signal_5855), .A1_f (new_AGEMA_signal_5856), .B0_t (Midori_rounds_SR_Inv_Result[10]), .B0_f (new_AGEMA_signal_5779), .B1_t (new_AGEMA_signal_5780), .B1_f (new_AGEMA_signal_5781), .Z0_t (Midori_rounds_Res_Inst_mux_inst_10_U1_X), .Z0_f (new_AGEMA_signal_6044), .Z1_t (new_AGEMA_signal_6045), .Z1_f (new_AGEMA_signal_6046) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_10_U1_X), .B0_f (new_AGEMA_signal_6044), .B1_t (new_AGEMA_signal_6045), .B1_f (new_AGEMA_signal_6046), .Z0_t (Midori_rounds_Res_Inst_mux_inst_10_U1_Y), .Z0_f (new_AGEMA_signal_6230), .Z1_t (new_AGEMA_signal_6231), .Z1_f (new_AGEMA_signal_6232) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_10_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_10_U1_Y), .A0_f (new_AGEMA_signal_6230), .A1_t (new_AGEMA_signal_6231), .A1_f (new_AGEMA_signal_6232), .B0_t (Midori_rounds_mul_ResultXORkey[10]), .B0_f (new_AGEMA_signal_5854), .B1_t (new_AGEMA_signal_5855), .B1_f (new_AGEMA_signal_5856), .Z0_t (Midori_rounds_round_Result[10]), .Z0_f (new_AGEMA_signal_6491), .Z1_t (new_AGEMA_signal_6492), .Z1_f (new_AGEMA_signal_6493) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_11_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[11]), .A0_f (new_AGEMA_signal_5712), .A1_t (new_AGEMA_signal_5713), .A1_f (new_AGEMA_signal_5714), .B0_t (Midori_rounds_SR_Inv_Result[11]), .B0_f (new_AGEMA_signal_5577), .B1_t (new_AGEMA_signal_5578), .B1_f (new_AGEMA_signal_5579), .Z0_t (Midori_rounds_Res_Inst_mux_inst_11_U1_X), .Z0_f (new_AGEMA_signal_5897), .Z1_t (new_AGEMA_signal_5898), .Z1_f (new_AGEMA_signal_5899) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_11_U1_X), .B0_f (new_AGEMA_signal_5897), .B1_t (new_AGEMA_signal_5898), .B1_f (new_AGEMA_signal_5899), .Z0_t (Midori_rounds_Res_Inst_mux_inst_11_U1_Y), .Z0_f (new_AGEMA_signal_6047), .Z1_t (new_AGEMA_signal_6048), .Z1_f (new_AGEMA_signal_6049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_11_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_11_U1_Y), .A0_f (new_AGEMA_signal_6047), .A1_t (new_AGEMA_signal_6048), .A1_f (new_AGEMA_signal_6049), .B0_t (Midori_rounds_mul_ResultXORkey[11]), .B0_f (new_AGEMA_signal_5712), .B1_t (new_AGEMA_signal_5713), .B1_f (new_AGEMA_signal_5714), .Z0_t (Midori_rounds_round_Result[11]), .Z0_f (new_AGEMA_signal_6233), .Z1_t (new_AGEMA_signal_6234), .Z1_f (new_AGEMA_signal_6235) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_12_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[12]), .A0_f (new_AGEMA_signal_6866), .A1_t (new_AGEMA_signal_6867), .A1_f (new_AGEMA_signal_6868), .B0_t (Midori_rounds_SR_Inv_Result[12]), .B0_f (new_AGEMA_signal_6773), .B1_t (new_AGEMA_signal_6774), .B1_f (new_AGEMA_signal_6775), .Z0_t (Midori_rounds_Res_Inst_mux_inst_12_U1_X), .Z0_f (new_AGEMA_signal_6923), .Z1_t (new_AGEMA_signal_6924), .Z1_f (new_AGEMA_signal_6925) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_12_U1_X), .B0_f (new_AGEMA_signal_6923), .B1_t (new_AGEMA_signal_6924), .B1_f (new_AGEMA_signal_6925), .Z0_t (Midori_rounds_Res_Inst_mux_inst_12_U1_Y), .Z0_f (new_AGEMA_signal_6986), .Z1_t (new_AGEMA_signal_6987), .Z1_f (new_AGEMA_signal_6988) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_12_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_12_U1_Y), .A0_f (new_AGEMA_signal_6986), .A1_t (new_AGEMA_signal_6987), .A1_f (new_AGEMA_signal_6988), .B0_t (Midori_rounds_mul_ResultXORkey[12]), .B0_f (new_AGEMA_signal_6866), .B1_t (new_AGEMA_signal_6867), .B1_f (new_AGEMA_signal_6868), .Z0_t (Midori_rounds_round_Result[12]), .Z0_f (new_AGEMA_signal_7055), .Z1_t (new_AGEMA_signal_7056), .Z1_f (new_AGEMA_signal_7057) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_13_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[13]), .A0_f (new_AGEMA_signal_5709), .A1_t (new_AGEMA_signal_5710), .A1_f (new_AGEMA_signal_5711), .B0_t (Midori_rounds_SR_Inv_Result[13]), .B0_f (new_AGEMA_signal_5568), .B1_t (new_AGEMA_signal_5569), .B1_f (new_AGEMA_signal_5570), .Z0_t (Midori_rounds_Res_Inst_mux_inst_13_U1_X), .Z0_f (new_AGEMA_signal_5900), .Z1_t (new_AGEMA_signal_5901), .Z1_f (new_AGEMA_signal_5902) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_13_U1_X), .B0_f (new_AGEMA_signal_5900), .B1_t (new_AGEMA_signal_5901), .B1_f (new_AGEMA_signal_5902), .Z0_t (Midori_rounds_Res_Inst_mux_inst_13_U1_Y), .Z0_f (new_AGEMA_signal_6050), .Z1_t (new_AGEMA_signal_6051), .Z1_f (new_AGEMA_signal_6052) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_13_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_13_U1_Y), .A0_f (new_AGEMA_signal_6050), .A1_t (new_AGEMA_signal_6051), .A1_f (new_AGEMA_signal_6052), .B0_t (Midori_rounds_mul_ResultXORkey[13]), .B0_f (new_AGEMA_signal_5709), .B1_t (new_AGEMA_signal_5710), .B1_f (new_AGEMA_signal_5711), .Z0_t (Midori_rounds_round_Result[13]), .Z0_f (new_AGEMA_signal_6236), .Z1_t (new_AGEMA_signal_6237), .Z1_f (new_AGEMA_signal_6238) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_14_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[14]), .A0_f (new_AGEMA_signal_5851), .A1_t (new_AGEMA_signal_5852), .A1_f (new_AGEMA_signal_5853), .B0_t (Midori_rounds_SR_Inv_Result[14]), .B0_f (new_AGEMA_signal_5770), .B1_t (new_AGEMA_signal_5771), .B1_f (new_AGEMA_signal_5772), .Z0_t (Midori_rounds_Res_Inst_mux_inst_14_U1_X), .Z0_f (new_AGEMA_signal_6053), .Z1_t (new_AGEMA_signal_6054), .Z1_f (new_AGEMA_signal_6055) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_14_U1_X), .B0_f (new_AGEMA_signal_6053), .B1_t (new_AGEMA_signal_6054), .B1_f (new_AGEMA_signal_6055), .Z0_t (Midori_rounds_Res_Inst_mux_inst_14_U1_Y), .Z0_f (new_AGEMA_signal_6239), .Z1_t (new_AGEMA_signal_6240), .Z1_f (new_AGEMA_signal_6241) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_14_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_14_U1_Y), .A0_f (new_AGEMA_signal_6239), .A1_t (new_AGEMA_signal_6240), .A1_f (new_AGEMA_signal_6241), .B0_t (Midori_rounds_mul_ResultXORkey[14]), .B0_f (new_AGEMA_signal_5851), .B1_t (new_AGEMA_signal_5852), .B1_f (new_AGEMA_signal_5853), .Z0_t (Midori_rounds_round_Result[14]), .Z0_f (new_AGEMA_signal_6494), .Z1_t (new_AGEMA_signal_6495), .Z1_f (new_AGEMA_signal_6496) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_15_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[15]), .A0_f (new_AGEMA_signal_5706), .A1_t (new_AGEMA_signal_5707), .A1_f (new_AGEMA_signal_5708), .B0_t (Midori_rounds_SR_Inv_Result[15]), .B0_f (new_AGEMA_signal_5553), .B1_t (new_AGEMA_signal_5554), .B1_f (new_AGEMA_signal_5555), .Z0_t (Midori_rounds_Res_Inst_mux_inst_15_U1_X), .Z0_f (new_AGEMA_signal_5903), .Z1_t (new_AGEMA_signal_5904), .Z1_f (new_AGEMA_signal_5905) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_15_U1_X), .B0_f (new_AGEMA_signal_5903), .B1_t (new_AGEMA_signal_5904), .B1_f (new_AGEMA_signal_5905), .Z0_t (Midori_rounds_Res_Inst_mux_inst_15_U1_Y), .Z0_f (new_AGEMA_signal_6056), .Z1_t (new_AGEMA_signal_6057), .Z1_f (new_AGEMA_signal_6058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_15_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_15_U1_Y), .A0_f (new_AGEMA_signal_6056), .A1_t (new_AGEMA_signal_6057), .A1_f (new_AGEMA_signal_6058), .B0_t (Midori_rounds_mul_ResultXORkey[15]), .B0_f (new_AGEMA_signal_5706), .B1_t (new_AGEMA_signal_5707), .B1_f (new_AGEMA_signal_5708), .Z0_t (Midori_rounds_round_Result[15]), .Z0_f (new_AGEMA_signal_6242), .Z1_t (new_AGEMA_signal_6243), .Z1_f (new_AGEMA_signal_6244) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_16_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[16]), .A0_f (new_AGEMA_signal_6794), .A1_t (new_AGEMA_signal_6795), .A1_f (new_AGEMA_signal_6796), .B0_t (Midori_rounds_SR_Inv_Result[16]), .B0_f (new_AGEMA_signal_6767), .B1_t (new_AGEMA_signal_6768), .B1_f (new_AGEMA_signal_6769), .Z0_t (Midori_rounds_Res_Inst_mux_inst_16_U1_X), .Z0_f (new_AGEMA_signal_6851), .Z1_t (new_AGEMA_signal_6852), .Z1_f (new_AGEMA_signal_6853) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_16_U1_X), .B0_f (new_AGEMA_signal_6851), .B1_t (new_AGEMA_signal_6852), .B1_f (new_AGEMA_signal_6853), .Z0_t (Midori_rounds_Res_Inst_mux_inst_16_U1_Y), .Z0_f (new_AGEMA_signal_6878), .Z1_t (new_AGEMA_signal_6879), .Z1_f (new_AGEMA_signal_6880) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_16_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_16_U1_Y), .A0_f (new_AGEMA_signal_6878), .A1_t (new_AGEMA_signal_6879), .A1_f (new_AGEMA_signal_6880), .B0_t (Midori_rounds_mul_ResultXORkey[16]), .B0_f (new_AGEMA_signal_6794), .B1_t (new_AGEMA_signal_6795), .B1_f (new_AGEMA_signal_6796), .Z0_t (Midori_rounds_round_Result[16]), .Z0_f (new_AGEMA_signal_6926), .Z1_t (new_AGEMA_signal_6927), .Z1_f (new_AGEMA_signal_6928) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_17_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[17]), .A0_f (new_AGEMA_signal_5703), .A1_t (new_AGEMA_signal_5704), .A1_f (new_AGEMA_signal_5705), .B0_t (Midori_rounds_SR_Inv_Result[17]), .B0_f (new_AGEMA_signal_5538), .B1_t (new_AGEMA_signal_5539), .B1_f (new_AGEMA_signal_5540), .Z0_t (Midori_rounds_Res_Inst_mux_inst_17_U1_X), .Z0_f (new_AGEMA_signal_5906), .Z1_t (new_AGEMA_signal_5907), .Z1_f (new_AGEMA_signal_5908) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_17_U1_X), .B0_f (new_AGEMA_signal_5906), .B1_t (new_AGEMA_signal_5907), .B1_f (new_AGEMA_signal_5908), .Z0_t (Midori_rounds_Res_Inst_mux_inst_17_U1_Y), .Z0_f (new_AGEMA_signal_6059), .Z1_t (new_AGEMA_signal_6060), .Z1_f (new_AGEMA_signal_6061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_17_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_17_U1_Y), .A0_f (new_AGEMA_signal_6059), .A1_t (new_AGEMA_signal_6060), .A1_f (new_AGEMA_signal_6061), .B0_t (Midori_rounds_mul_ResultXORkey[17]), .B0_f (new_AGEMA_signal_5703), .B1_t (new_AGEMA_signal_5704), .B1_f (new_AGEMA_signal_5705), .Z0_t (Midori_rounds_round_Result[17]), .Z0_f (new_AGEMA_signal_6245), .Z1_t (new_AGEMA_signal_6246), .Z1_f (new_AGEMA_signal_6247) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_18_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[18]), .A0_f (new_AGEMA_signal_5848), .A1_t (new_AGEMA_signal_5849), .A1_f (new_AGEMA_signal_5850), .B0_t (Midori_rounds_SR_Inv_Result[18]), .B0_f (new_AGEMA_signal_5758), .B1_t (new_AGEMA_signal_5759), .B1_f (new_AGEMA_signal_5760), .Z0_t (Midori_rounds_Res_Inst_mux_inst_18_U1_X), .Z0_f (new_AGEMA_signal_6062), .Z1_t (new_AGEMA_signal_6063), .Z1_f (new_AGEMA_signal_6064) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_18_U1_X), .B0_f (new_AGEMA_signal_6062), .B1_t (new_AGEMA_signal_6063), .B1_f (new_AGEMA_signal_6064), .Z0_t (Midori_rounds_Res_Inst_mux_inst_18_U1_Y), .Z0_f (new_AGEMA_signal_6248), .Z1_t (new_AGEMA_signal_6249), .Z1_f (new_AGEMA_signal_6250) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_18_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_18_U1_Y), .A0_f (new_AGEMA_signal_6248), .A1_t (new_AGEMA_signal_6249), .A1_f (new_AGEMA_signal_6250), .B0_t (Midori_rounds_mul_ResultXORkey[18]), .B0_f (new_AGEMA_signal_5848), .B1_t (new_AGEMA_signal_5849), .B1_f (new_AGEMA_signal_5850), .Z0_t (Midori_rounds_round_Result[18]), .Z0_f (new_AGEMA_signal_6497), .Z1_t (new_AGEMA_signal_6498), .Z1_f (new_AGEMA_signal_6499) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_19_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[19]), .A0_f (new_AGEMA_signal_5700), .A1_t (new_AGEMA_signal_5701), .A1_f (new_AGEMA_signal_5702), .B0_t (Midori_rounds_SR_Inv_Result[19]), .B0_f (new_AGEMA_signal_5523), .B1_t (new_AGEMA_signal_5524), .B1_f (new_AGEMA_signal_5525), .Z0_t (Midori_rounds_Res_Inst_mux_inst_19_U1_X), .Z0_f (new_AGEMA_signal_5909), .Z1_t (new_AGEMA_signal_5910), .Z1_f (new_AGEMA_signal_5911) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_19_U1_X), .B0_f (new_AGEMA_signal_5909), .B1_t (new_AGEMA_signal_5910), .B1_f (new_AGEMA_signal_5911), .Z0_t (Midori_rounds_Res_Inst_mux_inst_19_U1_Y), .Z0_f (new_AGEMA_signal_6065), .Z1_t (new_AGEMA_signal_6066), .Z1_f (new_AGEMA_signal_6067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_19_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_19_U1_Y), .A0_f (new_AGEMA_signal_6065), .A1_t (new_AGEMA_signal_6066), .A1_f (new_AGEMA_signal_6067), .B0_t (Midori_rounds_mul_ResultXORkey[19]), .B0_f (new_AGEMA_signal_5700), .B1_t (new_AGEMA_signal_5701), .B1_f (new_AGEMA_signal_5702), .Z0_t (Midori_rounds_round_Result[19]), .Z0_f (new_AGEMA_signal_6251), .Z1_t (new_AGEMA_signal_6252), .Z1_f (new_AGEMA_signal_6253) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_20_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[20]), .A0_f (new_AGEMA_signal_6791), .A1_t (new_AGEMA_signal_6792), .A1_f (new_AGEMA_signal_6793), .B0_t (Midori_rounds_SR_Inv_Result[20]), .B0_f (new_AGEMA_signal_6800), .B1_t (new_AGEMA_signal_6801), .B1_f (new_AGEMA_signal_6802), .Z0_t (Midori_rounds_Res_Inst_mux_inst_20_U1_X), .Z0_f (new_AGEMA_signal_6854), .Z1_t (new_AGEMA_signal_6855), .Z1_f (new_AGEMA_signal_6856) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_20_U1_X), .B0_f (new_AGEMA_signal_6854), .B1_t (new_AGEMA_signal_6855), .B1_f (new_AGEMA_signal_6856), .Z0_t (Midori_rounds_Res_Inst_mux_inst_20_U1_Y), .Z0_f (new_AGEMA_signal_6881), .Z1_t (new_AGEMA_signal_6882), .Z1_f (new_AGEMA_signal_6883) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_20_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_20_U1_Y), .A0_f (new_AGEMA_signal_6881), .A1_t (new_AGEMA_signal_6882), .A1_f (new_AGEMA_signal_6883), .B0_t (Midori_rounds_mul_ResultXORkey[20]), .B0_f (new_AGEMA_signal_6791), .B1_t (new_AGEMA_signal_6792), .B1_f (new_AGEMA_signal_6793), .Z0_t (Midori_rounds_round_Result[20]), .Z0_f (new_AGEMA_signal_6929), .Z1_t (new_AGEMA_signal_6930), .Z1_f (new_AGEMA_signal_6931) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_21_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[21]), .A0_f (new_AGEMA_signal_5697), .A1_t (new_AGEMA_signal_5698), .A1_f (new_AGEMA_signal_5699), .B0_t (Midori_rounds_SR_Inv_Result[21]), .B0_f (new_AGEMA_signal_5502), .B1_t (new_AGEMA_signal_5503), .B1_f (new_AGEMA_signal_5504), .Z0_t (Midori_rounds_Res_Inst_mux_inst_21_U1_X), .Z0_f (new_AGEMA_signal_5912), .Z1_t (new_AGEMA_signal_5913), .Z1_f (new_AGEMA_signal_5914) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_21_U1_X), .B0_f (new_AGEMA_signal_5912), .B1_t (new_AGEMA_signal_5913), .B1_f (new_AGEMA_signal_5914), .Z0_t (Midori_rounds_Res_Inst_mux_inst_21_U1_Y), .Z0_f (new_AGEMA_signal_6068), .Z1_t (new_AGEMA_signal_6069), .Z1_f (new_AGEMA_signal_6070) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_21_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_21_U1_Y), .A0_f (new_AGEMA_signal_6068), .A1_t (new_AGEMA_signal_6069), .A1_f (new_AGEMA_signal_6070), .B0_t (Midori_rounds_mul_ResultXORkey[21]), .B0_f (new_AGEMA_signal_5697), .B1_t (new_AGEMA_signal_5698), .B1_f (new_AGEMA_signal_5699), .Z0_t (Midori_rounds_round_Result[21]), .Z0_f (new_AGEMA_signal_6254), .Z1_t (new_AGEMA_signal_6255), .Z1_f (new_AGEMA_signal_6256) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_22_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[22]), .A0_f (new_AGEMA_signal_5845), .A1_t (new_AGEMA_signal_5846), .A1_f (new_AGEMA_signal_5847), .B0_t (Midori_rounds_SR_Inv_Result[22]), .B0_f (new_AGEMA_signal_5743), .B1_t (new_AGEMA_signal_5744), .B1_f (new_AGEMA_signal_5745), .Z0_t (Midori_rounds_Res_Inst_mux_inst_22_U1_X), .Z0_f (new_AGEMA_signal_6071), .Z1_t (new_AGEMA_signal_6072), .Z1_f (new_AGEMA_signal_6073) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_22_U1_X), .B0_f (new_AGEMA_signal_6071), .B1_t (new_AGEMA_signal_6072), .B1_f (new_AGEMA_signal_6073), .Z0_t (Midori_rounds_Res_Inst_mux_inst_22_U1_Y), .Z0_f (new_AGEMA_signal_6257), .Z1_t (new_AGEMA_signal_6258), .Z1_f (new_AGEMA_signal_6259) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_22_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_22_U1_Y), .A0_f (new_AGEMA_signal_6257), .A1_t (new_AGEMA_signal_6258), .A1_f (new_AGEMA_signal_6259), .B0_t (Midori_rounds_mul_ResultXORkey[22]), .B0_f (new_AGEMA_signal_5845), .B1_t (new_AGEMA_signal_5846), .B1_f (new_AGEMA_signal_5847), .Z0_t (Midori_rounds_round_Result[22]), .Z0_f (new_AGEMA_signal_6500), .Z1_t (new_AGEMA_signal_6501), .Z1_f (new_AGEMA_signal_6502) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_23_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[23]), .A0_f (new_AGEMA_signal_5694), .A1_t (new_AGEMA_signal_5695), .A1_f (new_AGEMA_signal_5696), .B0_t (Midori_rounds_SR_Inv_Result[23]), .B0_f (new_AGEMA_signal_5487), .B1_t (new_AGEMA_signal_5488), .B1_f (new_AGEMA_signal_5489), .Z0_t (Midori_rounds_Res_Inst_mux_inst_23_U1_X), .Z0_f (new_AGEMA_signal_5915), .Z1_t (new_AGEMA_signal_5916), .Z1_f (new_AGEMA_signal_5917) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_23_U1_X), .B0_f (new_AGEMA_signal_5915), .B1_t (new_AGEMA_signal_5916), .B1_f (new_AGEMA_signal_5917), .Z0_t (Midori_rounds_Res_Inst_mux_inst_23_U1_Y), .Z0_f (new_AGEMA_signal_6074), .Z1_t (new_AGEMA_signal_6075), .Z1_f (new_AGEMA_signal_6076) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_23_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_23_U1_Y), .A0_f (new_AGEMA_signal_6074), .A1_t (new_AGEMA_signal_6075), .A1_f (new_AGEMA_signal_6076), .B0_t (Midori_rounds_mul_ResultXORkey[23]), .B0_f (new_AGEMA_signal_5694), .B1_t (new_AGEMA_signal_5695), .B1_f (new_AGEMA_signal_5696), .Z0_t (Midori_rounds_round_Result[23]), .Z0_f (new_AGEMA_signal_6260), .Z1_t (new_AGEMA_signal_6261), .Z1_f (new_AGEMA_signal_6262) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_24_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[24]), .A0_f (new_AGEMA_signal_6833), .A1_t (new_AGEMA_signal_6834), .A1_f (new_AGEMA_signal_6835), .B0_t (Midori_rounds_SR_Inv_Result[24]), .B0_f (new_AGEMA_signal_6809), .B1_t (new_AGEMA_signal_6810), .B1_f (new_AGEMA_signal_6811), .Z0_t (Midori_rounds_Res_Inst_mux_inst_24_U1_X), .Z0_f (new_AGEMA_signal_6884), .Z1_t (new_AGEMA_signal_6885), .Z1_f (new_AGEMA_signal_6886) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_24_U1_X), .B0_f (new_AGEMA_signal_6884), .B1_t (new_AGEMA_signal_6885), .B1_f (new_AGEMA_signal_6886), .Z0_t (Midori_rounds_Res_Inst_mux_inst_24_U1_Y), .Z0_f (new_AGEMA_signal_6932), .Z1_t (new_AGEMA_signal_6933), .Z1_f (new_AGEMA_signal_6934) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_24_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_24_U1_Y), .A0_f (new_AGEMA_signal_6932), .A1_t (new_AGEMA_signal_6933), .A1_f (new_AGEMA_signal_6934), .B0_t (Midori_rounds_mul_ResultXORkey[24]), .B0_f (new_AGEMA_signal_6833), .B1_t (new_AGEMA_signal_6834), .B1_f (new_AGEMA_signal_6835), .Z0_t (Midori_rounds_round_Result[24]), .Z0_f (new_AGEMA_signal_6989), .Z1_t (new_AGEMA_signal_6990), .Z1_f (new_AGEMA_signal_6991) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_25_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[25]), .A0_f (new_AGEMA_signal_5691), .A1_t (new_AGEMA_signal_5692), .A1_f (new_AGEMA_signal_5693), .B0_t (Midori_rounds_SR_Inv_Result[25]), .B0_f (new_AGEMA_signal_5559), .B1_t (new_AGEMA_signal_5560), .B1_f (new_AGEMA_signal_5561), .Z0_t (Midori_rounds_Res_Inst_mux_inst_25_U1_X), .Z0_f (new_AGEMA_signal_5918), .Z1_t (new_AGEMA_signal_5919), .Z1_f (new_AGEMA_signal_5920) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_25_U1_X), .B0_f (new_AGEMA_signal_5918), .B1_t (new_AGEMA_signal_5919), .B1_f (new_AGEMA_signal_5920), .Z0_t (Midori_rounds_Res_Inst_mux_inst_25_U1_Y), .Z0_f (new_AGEMA_signal_6077), .Z1_t (new_AGEMA_signal_6078), .Z1_f (new_AGEMA_signal_6079) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_25_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_25_U1_Y), .A0_f (new_AGEMA_signal_6077), .A1_t (new_AGEMA_signal_6078), .A1_f (new_AGEMA_signal_6079), .B0_t (Midori_rounds_mul_ResultXORkey[25]), .B0_f (new_AGEMA_signal_5691), .B1_t (new_AGEMA_signal_5692), .B1_f (new_AGEMA_signal_5693), .Z0_t (Midori_rounds_round_Result[25]), .Z0_f (new_AGEMA_signal_6263), .Z1_t (new_AGEMA_signal_6264), .Z1_f (new_AGEMA_signal_6265) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_26_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[26]), .A0_f (new_AGEMA_signal_5842), .A1_t (new_AGEMA_signal_5843), .A1_f (new_AGEMA_signal_5844), .B0_t (Midori_rounds_SR_Inv_Result[26]), .B0_f (new_AGEMA_signal_5764), .B1_t (new_AGEMA_signal_5765), .B1_f (new_AGEMA_signal_5766), .Z0_t (Midori_rounds_Res_Inst_mux_inst_26_U1_X), .Z0_f (new_AGEMA_signal_6080), .Z1_t (new_AGEMA_signal_6081), .Z1_f (new_AGEMA_signal_6082) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_26_U1_X), .B0_f (new_AGEMA_signal_6080), .B1_t (new_AGEMA_signal_6081), .B1_f (new_AGEMA_signal_6082), .Z0_t (Midori_rounds_Res_Inst_mux_inst_26_U1_Y), .Z0_f (new_AGEMA_signal_6266), .Z1_t (new_AGEMA_signal_6267), .Z1_f (new_AGEMA_signal_6268) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_26_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_26_U1_Y), .A0_f (new_AGEMA_signal_6266), .A1_t (new_AGEMA_signal_6267), .A1_f (new_AGEMA_signal_6268), .B0_t (Midori_rounds_mul_ResultXORkey[26]), .B0_f (new_AGEMA_signal_5842), .B1_t (new_AGEMA_signal_5843), .B1_f (new_AGEMA_signal_5844), .Z0_t (Midori_rounds_round_Result[26]), .Z0_f (new_AGEMA_signal_6503), .Z1_t (new_AGEMA_signal_6504), .Z1_f (new_AGEMA_signal_6505) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_27_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[27]), .A0_f (new_AGEMA_signal_5688), .A1_t (new_AGEMA_signal_5689), .A1_f (new_AGEMA_signal_5690), .B0_t (Midori_rounds_SR_Inv_Result[27]), .B0_f (new_AGEMA_signal_5544), .B1_t (new_AGEMA_signal_5545), .B1_f (new_AGEMA_signal_5546), .Z0_t (Midori_rounds_Res_Inst_mux_inst_27_U1_X), .Z0_f (new_AGEMA_signal_5921), .Z1_t (new_AGEMA_signal_5922), .Z1_f (new_AGEMA_signal_5923) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_27_U1_X), .B0_f (new_AGEMA_signal_5921), .B1_t (new_AGEMA_signal_5922), .B1_f (new_AGEMA_signal_5923), .Z0_t (Midori_rounds_Res_Inst_mux_inst_27_U1_Y), .Z0_f (new_AGEMA_signal_6083), .Z1_t (new_AGEMA_signal_6084), .Z1_f (new_AGEMA_signal_6085) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_27_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_27_U1_Y), .A0_f (new_AGEMA_signal_6083), .A1_t (new_AGEMA_signal_6084), .A1_f (new_AGEMA_signal_6085), .B0_t (Midori_rounds_mul_ResultXORkey[27]), .B0_f (new_AGEMA_signal_5688), .B1_t (new_AGEMA_signal_5689), .B1_f (new_AGEMA_signal_5690), .Z0_t (Midori_rounds_round_Result[27]), .Z0_f (new_AGEMA_signal_6269), .Z1_t (new_AGEMA_signal_6270), .Z1_f (new_AGEMA_signal_6271) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_28_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[28]), .A0_f (new_AGEMA_signal_6827), .A1_t (new_AGEMA_signal_6828), .A1_f (new_AGEMA_signal_6829), .B0_t (Midori_rounds_SR_Inv_Result[28]), .B0_f (new_AGEMA_signal_6818), .B1_t (new_AGEMA_signal_6819), .B1_f (new_AGEMA_signal_6820), .Z0_t (Midori_rounds_Res_Inst_mux_inst_28_U1_X), .Z0_f (new_AGEMA_signal_6887), .Z1_t (new_AGEMA_signal_6888), .Z1_f (new_AGEMA_signal_6889) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_28_U1_X), .B0_f (new_AGEMA_signal_6887), .B1_t (new_AGEMA_signal_6888), .B1_f (new_AGEMA_signal_6889), .Z0_t (Midori_rounds_Res_Inst_mux_inst_28_U1_Y), .Z0_f (new_AGEMA_signal_6935), .Z1_t (new_AGEMA_signal_6936), .Z1_f (new_AGEMA_signal_6937) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_28_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_28_U1_Y), .A0_f (new_AGEMA_signal_6935), .A1_t (new_AGEMA_signal_6936), .A1_f (new_AGEMA_signal_6937), .B0_t (Midori_rounds_mul_ResultXORkey[28]), .B0_f (new_AGEMA_signal_6827), .B1_t (new_AGEMA_signal_6828), .B1_f (new_AGEMA_signal_6829), .Z0_t (Midori_rounds_round_Result[28]), .Z0_f (new_AGEMA_signal_6992), .Z1_t (new_AGEMA_signal_6993), .Z1_f (new_AGEMA_signal_6994) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_29_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[29]), .A0_f (new_AGEMA_signal_5685), .A1_t (new_AGEMA_signal_5686), .A1_f (new_AGEMA_signal_5687), .B0_t (Midori_rounds_SR_Inv_Result[29]), .B0_f (new_AGEMA_signal_5601), .B1_t (new_AGEMA_signal_5602), .B1_f (new_AGEMA_signal_5603), .Z0_t (Midori_rounds_Res_Inst_mux_inst_29_U1_X), .Z0_f (new_AGEMA_signal_5924), .Z1_t (new_AGEMA_signal_5925), .Z1_f (new_AGEMA_signal_5926) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_29_U1_X), .B0_f (new_AGEMA_signal_5924), .B1_t (new_AGEMA_signal_5925), .B1_f (new_AGEMA_signal_5926), .Z0_t (Midori_rounds_Res_Inst_mux_inst_29_U1_Y), .Z0_f (new_AGEMA_signal_6086), .Z1_t (new_AGEMA_signal_6087), .Z1_f (new_AGEMA_signal_6088) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_29_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_29_U1_Y), .A0_f (new_AGEMA_signal_6086), .A1_t (new_AGEMA_signal_6087), .A1_f (new_AGEMA_signal_6088), .B0_t (Midori_rounds_mul_ResultXORkey[29]), .B0_f (new_AGEMA_signal_5685), .B1_t (new_AGEMA_signal_5686), .B1_f (new_AGEMA_signal_5687), .Z0_t (Midori_rounds_round_Result[29]), .Z0_f (new_AGEMA_signal_6272), .Z1_t (new_AGEMA_signal_6273), .Z1_f (new_AGEMA_signal_6274) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_30_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[30]), .A0_f (new_AGEMA_signal_5839), .A1_t (new_AGEMA_signal_5840), .A1_f (new_AGEMA_signal_5841), .B0_t (Midori_rounds_SR_Inv_Result[30]), .B0_f (new_AGEMA_signal_5785), .B1_t (new_AGEMA_signal_5786), .B1_f (new_AGEMA_signal_5787), .Z0_t (Midori_rounds_Res_Inst_mux_inst_30_U1_X), .Z0_f (new_AGEMA_signal_6089), .Z1_t (new_AGEMA_signal_6090), .Z1_f (new_AGEMA_signal_6091) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_30_U1_X), .B0_f (new_AGEMA_signal_6089), .B1_t (new_AGEMA_signal_6090), .B1_f (new_AGEMA_signal_6091), .Z0_t (Midori_rounds_Res_Inst_mux_inst_30_U1_Y), .Z0_f (new_AGEMA_signal_6275), .Z1_t (new_AGEMA_signal_6276), .Z1_f (new_AGEMA_signal_6277) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_30_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_30_U1_Y), .A0_f (new_AGEMA_signal_6275), .A1_t (new_AGEMA_signal_6276), .A1_f (new_AGEMA_signal_6277), .B0_t (Midori_rounds_mul_ResultXORkey[30]), .B0_f (new_AGEMA_signal_5839), .B1_t (new_AGEMA_signal_5840), .B1_f (new_AGEMA_signal_5841), .Z0_t (Midori_rounds_round_Result[30]), .Z0_f (new_AGEMA_signal_6506), .Z1_t (new_AGEMA_signal_6507), .Z1_f (new_AGEMA_signal_6508) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_31_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[31]), .A0_f (new_AGEMA_signal_5682), .A1_t (new_AGEMA_signal_5683), .A1_f (new_AGEMA_signal_5684), .B0_t (Midori_rounds_SR_Inv_Result[31]), .B0_f (new_AGEMA_signal_5586), .B1_t (new_AGEMA_signal_5587), .B1_f (new_AGEMA_signal_5588), .Z0_t (Midori_rounds_Res_Inst_mux_inst_31_U1_X), .Z0_f (new_AGEMA_signal_5927), .Z1_t (new_AGEMA_signal_5928), .Z1_f (new_AGEMA_signal_5929) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_31_U1_X), .B0_f (new_AGEMA_signal_5927), .B1_t (new_AGEMA_signal_5928), .B1_f (new_AGEMA_signal_5929), .Z0_t (Midori_rounds_Res_Inst_mux_inst_31_U1_Y), .Z0_f (new_AGEMA_signal_6092), .Z1_t (new_AGEMA_signal_6093), .Z1_f (new_AGEMA_signal_6094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_31_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_31_U1_Y), .A0_f (new_AGEMA_signal_6092), .A1_t (new_AGEMA_signal_6093), .A1_f (new_AGEMA_signal_6094), .B0_t (Midori_rounds_mul_ResultXORkey[31]), .B0_f (new_AGEMA_signal_5682), .B1_t (new_AGEMA_signal_5683), .B1_f (new_AGEMA_signal_5684), .Z0_t (Midori_rounds_round_Result[31]), .Z0_f (new_AGEMA_signal_6278), .Z1_t (new_AGEMA_signal_6279), .Z1_f (new_AGEMA_signal_6280) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_32_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[32]), .A0_f (new_AGEMA_signal_6704), .A1_t (new_AGEMA_signal_6705), .A1_f (new_AGEMA_signal_6706), .B0_t (Midori_rounds_SR_Inv_Result[32]), .B0_f (new_AGEMA_signal_6842), .B1_t (new_AGEMA_signal_6843), .B1_f (new_AGEMA_signal_6844), .Z0_t (Midori_rounds_Res_Inst_mux_inst_32_U1_X), .Z0_f (new_AGEMA_signal_6890), .Z1_t (new_AGEMA_signal_6891), .Z1_f (new_AGEMA_signal_6892) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_32_U1_X), .B0_f (new_AGEMA_signal_6890), .B1_t (new_AGEMA_signal_6891), .B1_f (new_AGEMA_signal_6892), .Z0_t (Midori_rounds_Res_Inst_mux_inst_32_U1_Y), .Z0_f (new_AGEMA_signal_6938), .Z1_t (new_AGEMA_signal_6939), .Z1_f (new_AGEMA_signal_6940) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_32_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_32_U1_Y), .A0_f (new_AGEMA_signal_6938), .A1_t (new_AGEMA_signal_6939), .A1_f (new_AGEMA_signal_6940), .B0_t (Midori_rounds_mul_ResultXORkey[32]), .B0_f (new_AGEMA_signal_6704), .B1_t (new_AGEMA_signal_6705), .B1_f (new_AGEMA_signal_6706), .Z0_t (Midori_rounds_round_Result[32]), .Z0_f (new_AGEMA_signal_6995), .Z1_t (new_AGEMA_signal_6996), .Z1_f (new_AGEMA_signal_6997) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_33_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[33]), .A0_f (new_AGEMA_signal_5679), .A1_t (new_AGEMA_signal_5680), .A1_f (new_AGEMA_signal_5681), .B0_t (Midori_rounds_SR_Inv_Result[33]), .B0_f (new_AGEMA_signal_5589), .B1_t (new_AGEMA_signal_5590), .B1_f (new_AGEMA_signal_5591), .Z0_t (Midori_rounds_Res_Inst_mux_inst_33_U1_X), .Z0_f (new_AGEMA_signal_5930), .Z1_t (new_AGEMA_signal_5931), .Z1_f (new_AGEMA_signal_5932) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_33_U1_X), .B0_f (new_AGEMA_signal_5930), .B1_t (new_AGEMA_signal_5931), .B1_f (new_AGEMA_signal_5932), .Z0_t (Midori_rounds_Res_Inst_mux_inst_33_U1_Y), .Z0_f (new_AGEMA_signal_6095), .Z1_t (new_AGEMA_signal_6096), .Z1_f (new_AGEMA_signal_6097) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_33_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_33_U1_Y), .A0_f (new_AGEMA_signal_6095), .A1_t (new_AGEMA_signal_6096), .A1_f (new_AGEMA_signal_6097), .B0_t (Midori_rounds_mul_ResultXORkey[33]), .B0_f (new_AGEMA_signal_5679), .B1_t (new_AGEMA_signal_5680), .B1_f (new_AGEMA_signal_5681), .Z0_t (Midori_rounds_round_Result[33]), .Z0_f (new_AGEMA_signal_6281), .Z1_t (new_AGEMA_signal_6282), .Z1_f (new_AGEMA_signal_6283) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_34_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[34]), .A0_f (new_AGEMA_signal_5836), .A1_t (new_AGEMA_signal_5837), .A1_f (new_AGEMA_signal_5838), .B0_t (Midori_rounds_SR_Inv_Result[34]), .B0_f (new_AGEMA_signal_5776), .B1_t (new_AGEMA_signal_5777), .B1_f (new_AGEMA_signal_5778), .Z0_t (Midori_rounds_Res_Inst_mux_inst_34_U1_X), .Z0_f (new_AGEMA_signal_6098), .Z1_t (new_AGEMA_signal_6099), .Z1_f (new_AGEMA_signal_6100) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_34_U1_X), .B0_f (new_AGEMA_signal_6098), .B1_t (new_AGEMA_signal_6099), .B1_f (new_AGEMA_signal_6100), .Z0_t (Midori_rounds_Res_Inst_mux_inst_34_U1_Y), .Z0_f (new_AGEMA_signal_6284), .Z1_t (new_AGEMA_signal_6285), .Z1_f (new_AGEMA_signal_6286) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_34_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_34_U1_Y), .A0_f (new_AGEMA_signal_6284), .A1_t (new_AGEMA_signal_6285), .A1_f (new_AGEMA_signal_6286), .B0_t (Midori_rounds_mul_ResultXORkey[34]), .B0_f (new_AGEMA_signal_5836), .B1_t (new_AGEMA_signal_5837), .B1_f (new_AGEMA_signal_5838), .Z0_t (Midori_rounds_round_Result[34]), .Z0_f (new_AGEMA_signal_6509), .Z1_t (new_AGEMA_signal_6510), .Z1_f (new_AGEMA_signal_6511) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_35_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[35]), .A0_f (new_AGEMA_signal_5676), .A1_t (new_AGEMA_signal_5677), .A1_f (new_AGEMA_signal_5678), .B0_t (Midori_rounds_SR_Inv_Result[35]), .B0_f (new_AGEMA_signal_5574), .B1_t (new_AGEMA_signal_5575), .B1_f (new_AGEMA_signal_5576), .Z0_t (Midori_rounds_Res_Inst_mux_inst_35_U1_X), .Z0_f (new_AGEMA_signal_5933), .Z1_t (new_AGEMA_signal_5934), .Z1_f (new_AGEMA_signal_5935) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_35_U1_X), .B0_f (new_AGEMA_signal_5933), .B1_t (new_AGEMA_signal_5934), .B1_f (new_AGEMA_signal_5935), .Z0_t (Midori_rounds_Res_Inst_mux_inst_35_U1_Y), .Z0_f (new_AGEMA_signal_6101), .Z1_t (new_AGEMA_signal_6102), .Z1_f (new_AGEMA_signal_6103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_35_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_35_U1_Y), .A0_f (new_AGEMA_signal_6101), .A1_t (new_AGEMA_signal_6102), .A1_f (new_AGEMA_signal_6103), .B0_t (Midori_rounds_mul_ResultXORkey[35]), .B0_f (new_AGEMA_signal_5676), .B1_t (new_AGEMA_signal_5677), .B1_f (new_AGEMA_signal_5678), .Z0_t (Midori_rounds_round_Result[35]), .Z0_f (new_AGEMA_signal_6287), .Z1_t (new_AGEMA_signal_6288), .Z1_f (new_AGEMA_signal_6289) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_36_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[36]), .A0_f (new_AGEMA_signal_6788), .A1_t (new_AGEMA_signal_6789), .A1_f (new_AGEMA_signal_6790), .B0_t (Midori_rounds_SR_Inv_Result[36]), .B0_f (new_AGEMA_signal_6776), .B1_t (new_AGEMA_signal_6777), .B1_f (new_AGEMA_signal_6778), .Z0_t (Midori_rounds_Res_Inst_mux_inst_36_U1_X), .Z0_f (new_AGEMA_signal_6857), .Z1_t (new_AGEMA_signal_6858), .Z1_f (new_AGEMA_signal_6859) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_36_U1_X), .B0_f (new_AGEMA_signal_6857), .B1_t (new_AGEMA_signal_6858), .B1_f (new_AGEMA_signal_6859), .Z0_t (Midori_rounds_Res_Inst_mux_inst_36_U1_Y), .Z0_f (new_AGEMA_signal_6893), .Z1_t (new_AGEMA_signal_6894), .Z1_f (new_AGEMA_signal_6895) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_36_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_36_U1_Y), .A0_f (new_AGEMA_signal_6893), .A1_t (new_AGEMA_signal_6894), .A1_f (new_AGEMA_signal_6895), .B0_t (Midori_rounds_mul_ResultXORkey[36]), .B0_f (new_AGEMA_signal_6788), .B1_t (new_AGEMA_signal_6789), .B1_f (new_AGEMA_signal_6790), .Z0_t (Midori_rounds_round_Result[36]), .Z0_f (new_AGEMA_signal_6941), .Z1_t (new_AGEMA_signal_6942), .Z1_f (new_AGEMA_signal_6943) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_37_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[37]), .A0_f (new_AGEMA_signal_5673), .A1_t (new_AGEMA_signal_5674), .A1_f (new_AGEMA_signal_5675), .B0_t (Midori_rounds_SR_Inv_Result[37]), .B0_f (new_AGEMA_signal_5571), .B1_t (new_AGEMA_signal_5572), .B1_f (new_AGEMA_signal_5573), .Z0_t (Midori_rounds_Res_Inst_mux_inst_37_U1_X), .Z0_f (new_AGEMA_signal_5936), .Z1_t (new_AGEMA_signal_5937), .Z1_f (new_AGEMA_signal_5938) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_37_U1_X), .B0_f (new_AGEMA_signal_5936), .B1_t (new_AGEMA_signal_5937), .B1_f (new_AGEMA_signal_5938), .Z0_t (Midori_rounds_Res_Inst_mux_inst_37_U1_Y), .Z0_f (new_AGEMA_signal_6104), .Z1_t (new_AGEMA_signal_6105), .Z1_f (new_AGEMA_signal_6106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_37_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_37_U1_Y), .A0_f (new_AGEMA_signal_6104), .A1_t (new_AGEMA_signal_6105), .A1_f (new_AGEMA_signal_6106), .B0_t (Midori_rounds_mul_ResultXORkey[37]), .B0_f (new_AGEMA_signal_5673), .B1_t (new_AGEMA_signal_5674), .B1_f (new_AGEMA_signal_5675), .Z0_t (Midori_rounds_round_Result[37]), .Z0_f (new_AGEMA_signal_6290), .Z1_t (new_AGEMA_signal_6291), .Z1_f (new_AGEMA_signal_6292) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_38_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[38]), .A0_f (new_AGEMA_signal_5833), .A1_t (new_AGEMA_signal_5834), .A1_f (new_AGEMA_signal_5835), .B0_t (Midori_rounds_SR_Inv_Result[38]), .B0_f (new_AGEMA_signal_5773), .B1_t (new_AGEMA_signal_5774), .B1_f (new_AGEMA_signal_5775), .Z0_t (Midori_rounds_Res_Inst_mux_inst_38_U1_X), .Z0_f (new_AGEMA_signal_6107), .Z1_t (new_AGEMA_signal_6108), .Z1_f (new_AGEMA_signal_6109) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_38_U1_X), .B0_f (new_AGEMA_signal_6107), .B1_t (new_AGEMA_signal_6108), .B1_f (new_AGEMA_signal_6109), .Z0_t (Midori_rounds_Res_Inst_mux_inst_38_U1_Y), .Z0_f (new_AGEMA_signal_6293), .Z1_t (new_AGEMA_signal_6294), .Z1_f (new_AGEMA_signal_6295) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_38_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_38_U1_Y), .A0_f (new_AGEMA_signal_6293), .A1_t (new_AGEMA_signal_6294), .A1_f (new_AGEMA_signal_6295), .B0_t (Midori_rounds_mul_ResultXORkey[38]), .B0_f (new_AGEMA_signal_5833), .B1_t (new_AGEMA_signal_5834), .B1_f (new_AGEMA_signal_5835), .Z0_t (Midori_rounds_round_Result[38]), .Z0_f (new_AGEMA_signal_6512), .Z1_t (new_AGEMA_signal_6513), .Z1_f (new_AGEMA_signal_6514) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_39_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[39]), .A0_f (new_AGEMA_signal_5670), .A1_t (new_AGEMA_signal_5671), .A1_f (new_AGEMA_signal_5672), .B0_t (Midori_rounds_SR_Inv_Result[39]), .B0_f (new_AGEMA_signal_5556), .B1_t (new_AGEMA_signal_5557), .B1_f (new_AGEMA_signal_5558), .Z0_t (Midori_rounds_Res_Inst_mux_inst_39_U1_X), .Z0_f (new_AGEMA_signal_5939), .Z1_t (new_AGEMA_signal_5940), .Z1_f (new_AGEMA_signal_5941) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_39_U1_X), .B0_f (new_AGEMA_signal_5939), .B1_t (new_AGEMA_signal_5940), .B1_f (new_AGEMA_signal_5941), .Z0_t (Midori_rounds_Res_Inst_mux_inst_39_U1_Y), .Z0_f (new_AGEMA_signal_6110), .Z1_t (new_AGEMA_signal_6111), .Z1_f (new_AGEMA_signal_6112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_39_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_39_U1_Y), .A0_f (new_AGEMA_signal_6110), .A1_t (new_AGEMA_signal_6111), .A1_f (new_AGEMA_signal_6112), .B0_t (Midori_rounds_mul_ResultXORkey[39]), .B0_f (new_AGEMA_signal_5670), .B1_t (new_AGEMA_signal_5671), .B1_f (new_AGEMA_signal_5672), .Z0_t (Midori_rounds_round_Result[39]), .Z0_f (new_AGEMA_signal_6296), .Z1_t (new_AGEMA_signal_6297), .Z1_f (new_AGEMA_signal_6298) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_40_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[40]), .A0_f (new_AGEMA_signal_6839), .A1_t (new_AGEMA_signal_6840), .A1_f (new_AGEMA_signal_6841), .B0_t (Midori_rounds_SR_Inv_Result[40]), .B0_f (new_AGEMA_signal_6761), .B1_t (new_AGEMA_signal_6762), .B1_f (new_AGEMA_signal_6763), .Z0_t (Midori_rounds_Res_Inst_mux_inst_40_U1_X), .Z0_f (new_AGEMA_signal_6896), .Z1_t (new_AGEMA_signal_6897), .Z1_f (new_AGEMA_signal_6898) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_40_U1_X), .B0_f (new_AGEMA_signal_6896), .B1_t (new_AGEMA_signal_6897), .B1_f (new_AGEMA_signal_6898), .Z0_t (Midori_rounds_Res_Inst_mux_inst_40_U1_Y), .Z0_f (new_AGEMA_signal_6944), .Z1_t (new_AGEMA_signal_6945), .Z1_f (new_AGEMA_signal_6946) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_40_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_40_U1_Y), .A0_f (new_AGEMA_signal_6944), .A1_t (new_AGEMA_signal_6945), .A1_f (new_AGEMA_signal_6946), .B0_t (Midori_rounds_mul_ResultXORkey[40]), .B0_f (new_AGEMA_signal_6839), .B1_t (new_AGEMA_signal_6840), .B1_f (new_AGEMA_signal_6841), .Z0_t (Midori_rounds_round_Result[40]), .Z0_f (new_AGEMA_signal_6998), .Z1_t (new_AGEMA_signal_6999), .Z1_f (new_AGEMA_signal_7000) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_41_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[41]), .A0_f (new_AGEMA_signal_5667), .A1_t (new_AGEMA_signal_5668), .A1_f (new_AGEMA_signal_5669), .B0_t (Midori_rounds_SR_Inv_Result[41]), .B0_f (new_AGEMA_signal_5508), .B1_t (new_AGEMA_signal_5509), .B1_f (new_AGEMA_signal_5510), .Z0_t (Midori_rounds_Res_Inst_mux_inst_41_U1_X), .Z0_f (new_AGEMA_signal_5942), .Z1_t (new_AGEMA_signal_5943), .Z1_f (new_AGEMA_signal_5944) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_41_U1_X), .B0_f (new_AGEMA_signal_5942), .B1_t (new_AGEMA_signal_5943), .B1_f (new_AGEMA_signal_5944), .Z0_t (Midori_rounds_Res_Inst_mux_inst_41_U1_Y), .Z0_f (new_AGEMA_signal_6113), .Z1_t (new_AGEMA_signal_6114), .Z1_f (new_AGEMA_signal_6115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_41_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_41_U1_Y), .A0_f (new_AGEMA_signal_6113), .A1_t (new_AGEMA_signal_6114), .A1_f (new_AGEMA_signal_6115), .B0_t (Midori_rounds_mul_ResultXORkey[41]), .B0_f (new_AGEMA_signal_5667), .B1_t (new_AGEMA_signal_5668), .B1_f (new_AGEMA_signal_5669), .Z0_t (Midori_rounds_round_Result[41]), .Z0_f (new_AGEMA_signal_6299), .Z1_t (new_AGEMA_signal_6300), .Z1_f (new_AGEMA_signal_6301) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_42_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[42]), .A0_f (new_AGEMA_signal_5830), .A1_t (new_AGEMA_signal_5831), .A1_f (new_AGEMA_signal_5832), .B0_t (Midori_rounds_SR_Inv_Result[42]), .B0_f (new_AGEMA_signal_5746), .B1_t (new_AGEMA_signal_5747), .B1_f (new_AGEMA_signal_5748), .Z0_t (Midori_rounds_Res_Inst_mux_inst_42_U1_X), .Z0_f (new_AGEMA_signal_6116), .Z1_t (new_AGEMA_signal_6117), .Z1_f (new_AGEMA_signal_6118) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_42_U1_X), .B0_f (new_AGEMA_signal_6116), .B1_t (new_AGEMA_signal_6117), .B1_f (new_AGEMA_signal_6118), .Z0_t (Midori_rounds_Res_Inst_mux_inst_42_U1_Y), .Z0_f (new_AGEMA_signal_6302), .Z1_t (new_AGEMA_signal_6303), .Z1_f (new_AGEMA_signal_6304) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_42_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_42_U1_Y), .A0_f (new_AGEMA_signal_6302), .A1_t (new_AGEMA_signal_6303), .A1_f (new_AGEMA_signal_6304), .B0_t (Midori_rounds_mul_ResultXORkey[42]), .B0_f (new_AGEMA_signal_5830), .B1_t (new_AGEMA_signal_5831), .B1_f (new_AGEMA_signal_5832), .Z0_t (Midori_rounds_round_Result[42]), .Z0_f (new_AGEMA_signal_6515), .Z1_t (new_AGEMA_signal_6516), .Z1_f (new_AGEMA_signal_6517) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_43_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[43]), .A0_f (new_AGEMA_signal_5664), .A1_t (new_AGEMA_signal_5665), .A1_f (new_AGEMA_signal_5666), .B0_t (Midori_rounds_SR_Inv_Result[43]), .B0_f (new_AGEMA_signal_5493), .B1_t (new_AGEMA_signal_5494), .B1_f (new_AGEMA_signal_5495), .Z0_t (Midori_rounds_Res_Inst_mux_inst_43_U1_X), .Z0_f (new_AGEMA_signal_5945), .Z1_t (new_AGEMA_signal_5946), .Z1_f (new_AGEMA_signal_5947) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_43_U1_X), .B0_f (new_AGEMA_signal_5945), .B1_t (new_AGEMA_signal_5946), .B1_f (new_AGEMA_signal_5947), .Z0_t (Midori_rounds_Res_Inst_mux_inst_43_U1_Y), .Z0_f (new_AGEMA_signal_6119), .Z1_t (new_AGEMA_signal_6120), .Z1_f (new_AGEMA_signal_6121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_43_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_43_U1_Y), .A0_f (new_AGEMA_signal_6119), .A1_t (new_AGEMA_signal_6120), .A1_f (new_AGEMA_signal_6121), .B0_t (Midori_rounds_mul_ResultXORkey[43]), .B0_f (new_AGEMA_signal_5664), .B1_t (new_AGEMA_signal_5665), .B1_f (new_AGEMA_signal_5666), .Z0_t (Midori_rounds_round_Result[43]), .Z0_f (new_AGEMA_signal_6305), .Z1_t (new_AGEMA_signal_6306), .Z1_f (new_AGEMA_signal_6307) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_44_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[44]), .A0_f (new_AGEMA_signal_6830), .A1_t (new_AGEMA_signal_6831), .A1_f (new_AGEMA_signal_6832), .B0_t (Midori_rounds_SR_Inv_Result[44]), .B0_f (new_AGEMA_signal_6806), .B1_t (new_AGEMA_signal_6807), .B1_f (new_AGEMA_signal_6808), .Z0_t (Midori_rounds_Res_Inst_mux_inst_44_U1_X), .Z0_f (new_AGEMA_signal_6899), .Z1_t (new_AGEMA_signal_6900), .Z1_f (new_AGEMA_signal_6901) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_44_U1_X), .B0_f (new_AGEMA_signal_6899), .B1_t (new_AGEMA_signal_6900), .B1_f (new_AGEMA_signal_6901), .Z0_t (Midori_rounds_Res_Inst_mux_inst_44_U1_Y), .Z0_f (new_AGEMA_signal_6947), .Z1_t (new_AGEMA_signal_6948), .Z1_f (new_AGEMA_signal_6949) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_44_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_44_U1_Y), .A0_f (new_AGEMA_signal_6947), .A1_t (new_AGEMA_signal_6948), .A1_f (new_AGEMA_signal_6949), .B0_t (Midori_rounds_mul_ResultXORkey[44]), .B0_f (new_AGEMA_signal_6830), .B1_t (new_AGEMA_signal_6831), .B1_f (new_AGEMA_signal_6832), .Z0_t (Midori_rounds_round_Result[44]), .Z0_f (new_AGEMA_signal_7001), .Z1_t (new_AGEMA_signal_7002), .Z1_f (new_AGEMA_signal_7003) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_45_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[45]), .A0_f (new_AGEMA_signal_5661), .A1_t (new_AGEMA_signal_5662), .A1_f (new_AGEMA_signal_5663), .B0_t (Midori_rounds_SR_Inv_Result[45]), .B0_f (new_AGEMA_signal_5532), .B1_t (new_AGEMA_signal_5533), .B1_f (new_AGEMA_signal_5534), .Z0_t (Midori_rounds_Res_Inst_mux_inst_45_U1_X), .Z0_f (new_AGEMA_signal_5948), .Z1_t (new_AGEMA_signal_5949), .Z1_f (new_AGEMA_signal_5950) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_45_U1_X), .B0_f (new_AGEMA_signal_5948), .B1_t (new_AGEMA_signal_5949), .B1_f (new_AGEMA_signal_5950), .Z0_t (Midori_rounds_Res_Inst_mux_inst_45_U1_Y), .Z0_f (new_AGEMA_signal_6122), .Z1_t (new_AGEMA_signal_6123), .Z1_f (new_AGEMA_signal_6124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_45_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_45_U1_Y), .A0_f (new_AGEMA_signal_6122), .A1_t (new_AGEMA_signal_6123), .A1_f (new_AGEMA_signal_6124), .B0_t (Midori_rounds_mul_ResultXORkey[45]), .B0_f (new_AGEMA_signal_5661), .B1_t (new_AGEMA_signal_5662), .B1_f (new_AGEMA_signal_5663), .Z0_t (Midori_rounds_round_Result[45]), .Z0_f (new_AGEMA_signal_6308), .Z1_t (new_AGEMA_signal_6309), .Z1_f (new_AGEMA_signal_6310) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_46_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[46]), .A0_f (new_AGEMA_signal_5827), .A1_t (new_AGEMA_signal_5828), .A1_f (new_AGEMA_signal_5829), .B0_t (Midori_rounds_SR_Inv_Result[46]), .B0_f (new_AGEMA_signal_5755), .B1_t (new_AGEMA_signal_5756), .B1_f (new_AGEMA_signal_5757), .Z0_t (Midori_rounds_Res_Inst_mux_inst_46_U1_X), .Z0_f (new_AGEMA_signal_6125), .Z1_t (new_AGEMA_signal_6126), .Z1_f (new_AGEMA_signal_6127) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_46_U1_X), .B0_f (new_AGEMA_signal_6125), .B1_t (new_AGEMA_signal_6126), .B1_f (new_AGEMA_signal_6127), .Z0_t (Midori_rounds_Res_Inst_mux_inst_46_U1_Y), .Z0_f (new_AGEMA_signal_6311), .Z1_t (new_AGEMA_signal_6312), .Z1_f (new_AGEMA_signal_6313) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_46_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_46_U1_Y), .A0_f (new_AGEMA_signal_6311), .A1_t (new_AGEMA_signal_6312), .A1_f (new_AGEMA_signal_6313), .B0_t (Midori_rounds_mul_ResultXORkey[46]), .B0_f (new_AGEMA_signal_5827), .B1_t (new_AGEMA_signal_5828), .B1_f (new_AGEMA_signal_5829), .Z0_t (Midori_rounds_round_Result[46]), .Z0_f (new_AGEMA_signal_6518), .Z1_t (new_AGEMA_signal_6519), .Z1_f (new_AGEMA_signal_6520) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_47_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[47]), .A0_f (new_AGEMA_signal_5658), .A1_t (new_AGEMA_signal_5659), .A1_f (new_AGEMA_signal_5660), .B0_t (Midori_rounds_SR_Inv_Result[47]), .B0_f (new_AGEMA_signal_5517), .B1_t (new_AGEMA_signal_5518), .B1_f (new_AGEMA_signal_5519), .Z0_t (Midori_rounds_Res_Inst_mux_inst_47_U1_X), .Z0_f (new_AGEMA_signal_5951), .Z1_t (new_AGEMA_signal_5952), .Z1_f (new_AGEMA_signal_5953) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_47_U1_X), .B0_f (new_AGEMA_signal_5951), .B1_t (new_AGEMA_signal_5952), .B1_f (new_AGEMA_signal_5953), .Z0_t (Midori_rounds_Res_Inst_mux_inst_47_U1_Y), .Z0_f (new_AGEMA_signal_6128), .Z1_t (new_AGEMA_signal_6129), .Z1_f (new_AGEMA_signal_6130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_47_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_47_U1_Y), .A0_f (new_AGEMA_signal_6128), .A1_t (new_AGEMA_signal_6129), .A1_f (new_AGEMA_signal_6130), .B0_t (Midori_rounds_mul_ResultXORkey[47]), .B0_f (new_AGEMA_signal_5658), .B1_t (new_AGEMA_signal_5659), .B1_f (new_AGEMA_signal_5660), .Z0_t (Midori_rounds_round_Result[47]), .Z0_f (new_AGEMA_signal_6314), .Z1_t (new_AGEMA_signal_6315), .Z1_f (new_AGEMA_signal_6316) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_48_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[48]), .A0_f (new_AGEMA_signal_6701), .A1_t (new_AGEMA_signal_6702), .A1_f (new_AGEMA_signal_6703), .B0_t (Midori_rounds_SR_Inv_Result[48]), .B0_f (new_AGEMA_signal_6812), .B1_t (new_AGEMA_signal_6813), .B1_f (new_AGEMA_signal_6814), .Z0_t (Midori_rounds_Res_Inst_mux_inst_48_U1_X), .Z0_f (new_AGEMA_signal_6860), .Z1_t (new_AGEMA_signal_6861), .Z1_f (new_AGEMA_signal_6862) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_48_U1_X), .B0_f (new_AGEMA_signal_6860), .B1_t (new_AGEMA_signal_6861), .B1_f (new_AGEMA_signal_6862), .Z0_t (Midori_rounds_Res_Inst_mux_inst_48_U1_Y), .Z0_f (new_AGEMA_signal_6902), .Z1_t (new_AGEMA_signal_6903), .Z1_f (new_AGEMA_signal_6904) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_48_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_48_U1_Y), .A0_f (new_AGEMA_signal_6902), .A1_t (new_AGEMA_signal_6903), .A1_f (new_AGEMA_signal_6904), .B0_t (Midori_rounds_mul_ResultXORkey[48]), .B0_f (new_AGEMA_signal_6701), .B1_t (new_AGEMA_signal_6702), .B1_f (new_AGEMA_signal_6703), .Z0_t (Midori_rounds_round_Result[48]), .Z0_f (new_AGEMA_signal_6950), .Z1_t (new_AGEMA_signal_6951), .Z1_f (new_AGEMA_signal_6952) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_49_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[49]), .A0_f (new_AGEMA_signal_5655), .A1_t (new_AGEMA_signal_5656), .A1_f (new_AGEMA_signal_5657), .B0_t (Midori_rounds_SR_Inv_Result[49]), .B0_f (new_AGEMA_signal_5562), .B1_t (new_AGEMA_signal_5563), .B1_f (new_AGEMA_signal_5564), .Z0_t (Midori_rounds_Res_Inst_mux_inst_49_U1_X), .Z0_f (new_AGEMA_signal_5954), .Z1_t (new_AGEMA_signal_5955), .Z1_f (new_AGEMA_signal_5956) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_49_U1_X), .B0_f (new_AGEMA_signal_5954), .B1_t (new_AGEMA_signal_5955), .B1_f (new_AGEMA_signal_5956), .Z0_t (Midori_rounds_Res_Inst_mux_inst_49_U1_Y), .Z0_f (new_AGEMA_signal_6131), .Z1_t (new_AGEMA_signal_6132), .Z1_f (new_AGEMA_signal_6133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_49_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_49_U1_Y), .A0_f (new_AGEMA_signal_6131), .A1_t (new_AGEMA_signal_6132), .A1_f (new_AGEMA_signal_6133), .B0_t (Midori_rounds_mul_ResultXORkey[49]), .B0_f (new_AGEMA_signal_5655), .B1_t (new_AGEMA_signal_5656), .B1_f (new_AGEMA_signal_5657), .Z0_t (Midori_rounds_round_Result[49]), .Z0_f (new_AGEMA_signal_6317), .Z1_t (new_AGEMA_signal_6318), .Z1_f (new_AGEMA_signal_6319) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_50_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[50]), .A0_f (new_AGEMA_signal_5824), .A1_t (new_AGEMA_signal_5825), .A1_f (new_AGEMA_signal_5826), .B0_t (Midori_rounds_SR_Inv_Result[50]), .B0_f (new_AGEMA_signal_5767), .B1_t (new_AGEMA_signal_5768), .B1_f (new_AGEMA_signal_5769), .Z0_t (Midori_rounds_Res_Inst_mux_inst_50_U1_X), .Z0_f (new_AGEMA_signal_6134), .Z1_t (new_AGEMA_signal_6135), .Z1_f (new_AGEMA_signal_6136) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_50_U1_X), .B0_f (new_AGEMA_signal_6134), .B1_t (new_AGEMA_signal_6135), .B1_f (new_AGEMA_signal_6136), .Z0_t (Midori_rounds_Res_Inst_mux_inst_50_U1_Y), .Z0_f (new_AGEMA_signal_6320), .Z1_t (new_AGEMA_signal_6321), .Z1_f (new_AGEMA_signal_6322) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_50_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_50_U1_Y), .A0_f (new_AGEMA_signal_6320), .A1_t (new_AGEMA_signal_6321), .A1_f (new_AGEMA_signal_6322), .B0_t (Midori_rounds_mul_ResultXORkey[50]), .B0_f (new_AGEMA_signal_5824), .B1_t (new_AGEMA_signal_5825), .B1_f (new_AGEMA_signal_5826), .Z0_t (Midori_rounds_round_Result[50]), .Z0_f (new_AGEMA_signal_6521), .Z1_t (new_AGEMA_signal_6522), .Z1_f (new_AGEMA_signal_6523) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_51_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[51]), .A0_f (new_AGEMA_signal_5652), .A1_t (new_AGEMA_signal_5653), .A1_f (new_AGEMA_signal_5654), .B0_t (Midori_rounds_SR_Inv_Result[51]), .B0_f (new_AGEMA_signal_5547), .B1_t (new_AGEMA_signal_5548), .B1_f (new_AGEMA_signal_5549), .Z0_t (Midori_rounds_Res_Inst_mux_inst_51_U1_X), .Z0_f (new_AGEMA_signal_5957), .Z1_t (new_AGEMA_signal_5958), .Z1_f (new_AGEMA_signal_5959) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_51_U1_X), .B0_f (new_AGEMA_signal_5957), .B1_t (new_AGEMA_signal_5958), .B1_f (new_AGEMA_signal_5959), .Z0_t (Midori_rounds_Res_Inst_mux_inst_51_U1_Y), .Z0_f (new_AGEMA_signal_6137), .Z1_t (new_AGEMA_signal_6138), .Z1_f (new_AGEMA_signal_6139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_51_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_51_U1_Y), .A0_f (new_AGEMA_signal_6137), .A1_t (new_AGEMA_signal_6138), .A1_f (new_AGEMA_signal_6139), .B0_t (Midori_rounds_mul_ResultXORkey[51]), .B0_f (new_AGEMA_signal_5652), .B1_t (new_AGEMA_signal_5653), .B1_f (new_AGEMA_signal_5654), .Z0_t (Midori_rounds_round_Result[51]), .Z0_f (new_AGEMA_signal_6323), .Z1_t (new_AGEMA_signal_6324), .Z1_f (new_AGEMA_signal_6325) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_52_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[52]), .A0_f (new_AGEMA_signal_6785), .A1_t (new_AGEMA_signal_6786), .A1_f (new_AGEMA_signal_6787), .B0_t (Midori_rounds_SR_Inv_Result[52]), .B0_f (new_AGEMA_signal_6779), .B1_t (new_AGEMA_signal_6780), .B1_f (new_AGEMA_signal_6781), .Z0_t (Midori_rounds_Res_Inst_mux_inst_52_U1_X), .Z0_f (new_AGEMA_signal_6863), .Z1_t (new_AGEMA_signal_6864), .Z1_f (new_AGEMA_signal_6865) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_52_U1_X), .B0_f (new_AGEMA_signal_6863), .B1_t (new_AGEMA_signal_6864), .B1_f (new_AGEMA_signal_6865), .Z0_t (Midori_rounds_Res_Inst_mux_inst_52_U1_Y), .Z0_f (new_AGEMA_signal_6905), .Z1_t (new_AGEMA_signal_6906), .Z1_f (new_AGEMA_signal_6907) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_52_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_52_U1_Y), .A0_f (new_AGEMA_signal_6905), .A1_t (new_AGEMA_signal_6906), .A1_f (new_AGEMA_signal_6907), .B0_t (Midori_rounds_mul_ResultXORkey[52]), .B0_f (new_AGEMA_signal_6785), .B1_t (new_AGEMA_signal_6786), .B1_f (new_AGEMA_signal_6787), .Z0_t (Midori_rounds_round_Result[52]), .Z0_f (new_AGEMA_signal_6953), .Z1_t (new_AGEMA_signal_6954), .Z1_f (new_AGEMA_signal_6955) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_53_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[53]), .A0_f (new_AGEMA_signal_5649), .A1_t (new_AGEMA_signal_5650), .A1_f (new_AGEMA_signal_5651), .B0_t (Midori_rounds_SR_Inv_Result[53]), .B0_f (new_AGEMA_signal_5598), .B1_t (new_AGEMA_signal_5599), .B1_f (new_AGEMA_signal_5600), .Z0_t (Midori_rounds_Res_Inst_mux_inst_53_U1_X), .Z0_f (new_AGEMA_signal_5960), .Z1_t (new_AGEMA_signal_5961), .Z1_f (new_AGEMA_signal_5962) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_53_U1_X), .B0_f (new_AGEMA_signal_5960), .B1_t (new_AGEMA_signal_5961), .B1_f (new_AGEMA_signal_5962), .Z0_t (Midori_rounds_Res_Inst_mux_inst_53_U1_Y), .Z0_f (new_AGEMA_signal_6140), .Z1_t (new_AGEMA_signal_6141), .Z1_f (new_AGEMA_signal_6142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_53_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_53_U1_Y), .A0_f (new_AGEMA_signal_6140), .A1_t (new_AGEMA_signal_6141), .A1_f (new_AGEMA_signal_6142), .B0_t (Midori_rounds_mul_ResultXORkey[53]), .B0_f (new_AGEMA_signal_5649), .B1_t (new_AGEMA_signal_5650), .B1_f (new_AGEMA_signal_5651), .Z0_t (Midori_rounds_round_Result[53]), .Z0_f (new_AGEMA_signal_6326), .Z1_t (new_AGEMA_signal_6327), .Z1_f (new_AGEMA_signal_6328) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_54_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[54]), .A0_f (new_AGEMA_signal_5821), .A1_t (new_AGEMA_signal_5822), .A1_f (new_AGEMA_signal_5823), .B0_t (Midori_rounds_SR_Inv_Result[54]), .B0_f (new_AGEMA_signal_5782), .B1_t (new_AGEMA_signal_5783), .B1_f (new_AGEMA_signal_5784), .Z0_t (Midori_rounds_Res_Inst_mux_inst_54_U1_X), .Z0_f (new_AGEMA_signal_6143), .Z1_t (new_AGEMA_signal_6144), .Z1_f (new_AGEMA_signal_6145) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_54_U1_X), .B0_f (new_AGEMA_signal_6143), .B1_t (new_AGEMA_signal_6144), .B1_f (new_AGEMA_signal_6145), .Z0_t (Midori_rounds_Res_Inst_mux_inst_54_U1_Y), .Z0_f (new_AGEMA_signal_6329), .Z1_t (new_AGEMA_signal_6330), .Z1_f (new_AGEMA_signal_6331) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_54_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_54_U1_Y), .A0_f (new_AGEMA_signal_6329), .A1_t (new_AGEMA_signal_6330), .A1_f (new_AGEMA_signal_6331), .B0_t (Midori_rounds_mul_ResultXORkey[54]), .B0_f (new_AGEMA_signal_5821), .B1_t (new_AGEMA_signal_5822), .B1_f (new_AGEMA_signal_5823), .Z0_t (Midori_rounds_round_Result[54]), .Z0_f (new_AGEMA_signal_6524), .Z1_t (new_AGEMA_signal_6525), .Z1_f (new_AGEMA_signal_6526) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_55_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[55]), .A0_f (new_AGEMA_signal_5646), .A1_t (new_AGEMA_signal_5647), .A1_f (new_AGEMA_signal_5648), .B0_t (Midori_rounds_SR_Inv_Result[55]), .B0_f (new_AGEMA_signal_5583), .B1_t (new_AGEMA_signal_5584), .B1_f (new_AGEMA_signal_5585), .Z0_t (Midori_rounds_Res_Inst_mux_inst_55_U1_X), .Z0_f (new_AGEMA_signal_5963), .Z1_t (new_AGEMA_signal_5964), .Z1_f (new_AGEMA_signal_5965) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_55_U1_X), .B0_f (new_AGEMA_signal_5963), .B1_t (new_AGEMA_signal_5964), .B1_f (new_AGEMA_signal_5965), .Z0_t (Midori_rounds_Res_Inst_mux_inst_55_U1_Y), .Z0_f (new_AGEMA_signal_6146), .Z1_t (new_AGEMA_signal_6147), .Z1_f (new_AGEMA_signal_6148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_55_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_55_U1_Y), .A0_f (new_AGEMA_signal_6146), .A1_t (new_AGEMA_signal_6147), .A1_f (new_AGEMA_signal_6148), .B0_t (Midori_rounds_mul_ResultXORkey[55]), .B0_f (new_AGEMA_signal_5646), .B1_t (new_AGEMA_signal_5647), .B1_f (new_AGEMA_signal_5648), .Z0_t (Midori_rounds_round_Result[55]), .Z0_f (new_AGEMA_signal_6332), .Z1_t (new_AGEMA_signal_6333), .Z1_f (new_AGEMA_signal_6334) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_56_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[56]), .A0_f (new_AGEMA_signal_6824), .A1_t (new_AGEMA_signal_6825), .A1_f (new_AGEMA_signal_6826), .B0_t (Midori_rounds_SR_Inv_Result[56]), .B0_f (new_AGEMA_signal_6692), .B1_t (new_AGEMA_signal_6693), .B1_f (new_AGEMA_signal_6694), .Z0_t (Midori_rounds_Res_Inst_mux_inst_56_U1_X), .Z0_f (new_AGEMA_signal_6908), .Z1_t (new_AGEMA_signal_6909), .Z1_f (new_AGEMA_signal_6910) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_56_U1_X), .B0_f (new_AGEMA_signal_6908), .B1_t (new_AGEMA_signal_6909), .B1_f (new_AGEMA_signal_6910), .Z0_t (Midori_rounds_Res_Inst_mux_inst_56_U1_Y), .Z0_f (new_AGEMA_signal_6956), .Z1_t (new_AGEMA_signal_6957), .Z1_f (new_AGEMA_signal_6958) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_56_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_56_U1_Y), .A0_f (new_AGEMA_signal_6956), .A1_t (new_AGEMA_signal_6957), .A1_f (new_AGEMA_signal_6958), .B0_t (Midori_rounds_mul_ResultXORkey[56]), .B0_f (new_AGEMA_signal_6824), .B1_t (new_AGEMA_signal_6825), .B1_f (new_AGEMA_signal_6826), .Z0_t (Midori_rounds_round_Result[56]), .Z0_f (new_AGEMA_signal_7004), .Z1_t (new_AGEMA_signal_7005), .Z1_f (new_AGEMA_signal_7006) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_57_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[57]), .A0_f (new_AGEMA_signal_5643), .A1_t (new_AGEMA_signal_5644), .A1_f (new_AGEMA_signal_5645), .B0_t (Midori_rounds_SR_Inv_Result[57]), .B0_f (new_AGEMA_signal_5541), .B1_t (new_AGEMA_signal_5542), .B1_f (new_AGEMA_signal_5543), .Z0_t (Midori_rounds_Res_Inst_mux_inst_57_U1_X), .Z0_f (new_AGEMA_signal_5966), .Z1_t (new_AGEMA_signal_5967), .Z1_f (new_AGEMA_signal_5968) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_57_U1_X), .B0_f (new_AGEMA_signal_5966), .B1_t (new_AGEMA_signal_5967), .B1_f (new_AGEMA_signal_5968), .Z0_t (Midori_rounds_Res_Inst_mux_inst_57_U1_Y), .Z0_f (new_AGEMA_signal_6149), .Z1_t (new_AGEMA_signal_6150), .Z1_f (new_AGEMA_signal_6151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_57_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_57_U1_Y), .A0_f (new_AGEMA_signal_6149), .A1_t (new_AGEMA_signal_6150), .A1_f (new_AGEMA_signal_6151), .B0_t (Midori_rounds_mul_ResultXORkey[57]), .B0_f (new_AGEMA_signal_5643), .B1_t (new_AGEMA_signal_5644), .B1_f (new_AGEMA_signal_5645), .Z0_t (Midori_rounds_round_Result[57]), .Z0_f (new_AGEMA_signal_6335), .Z1_t (new_AGEMA_signal_6336), .Z1_f (new_AGEMA_signal_6337) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_58_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[58]), .A0_f (new_AGEMA_signal_5818), .A1_t (new_AGEMA_signal_5819), .A1_f (new_AGEMA_signal_5820), .B0_t (Midori_rounds_SR_Inv_Result[58]), .B0_f (new_AGEMA_signal_5761), .B1_t (new_AGEMA_signal_5762), .B1_f (new_AGEMA_signal_5763), .Z0_t (Midori_rounds_Res_Inst_mux_inst_58_U1_X), .Z0_f (new_AGEMA_signal_6152), .Z1_t (new_AGEMA_signal_6153), .Z1_f (new_AGEMA_signal_6154) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_58_U1_X), .B0_f (new_AGEMA_signal_6152), .B1_t (new_AGEMA_signal_6153), .B1_f (new_AGEMA_signal_6154), .Z0_t (Midori_rounds_Res_Inst_mux_inst_58_U1_Y), .Z0_f (new_AGEMA_signal_6338), .Z1_t (new_AGEMA_signal_6339), .Z1_f (new_AGEMA_signal_6340) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_58_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_58_U1_Y), .A0_f (new_AGEMA_signal_6338), .A1_t (new_AGEMA_signal_6339), .A1_f (new_AGEMA_signal_6340), .B0_t (Midori_rounds_mul_ResultXORkey[58]), .B0_f (new_AGEMA_signal_5818), .B1_t (new_AGEMA_signal_5819), .B1_f (new_AGEMA_signal_5820), .Z0_t (Midori_rounds_round_Result[58]), .Z0_f (new_AGEMA_signal_6527), .Z1_t (new_AGEMA_signal_6528), .Z1_f (new_AGEMA_signal_6529) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_59_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[59]), .A0_f (new_AGEMA_signal_5640), .A1_t (new_AGEMA_signal_5641), .A1_f (new_AGEMA_signal_5642), .B0_t (Midori_rounds_SR_Inv_Result[59]), .B0_f (new_AGEMA_signal_5526), .B1_t (new_AGEMA_signal_5527), .B1_f (new_AGEMA_signal_5528), .Z0_t (Midori_rounds_Res_Inst_mux_inst_59_U1_X), .Z0_f (new_AGEMA_signal_5969), .Z1_t (new_AGEMA_signal_5970), .Z1_f (new_AGEMA_signal_5971) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_59_U1_X), .B0_f (new_AGEMA_signal_5969), .B1_t (new_AGEMA_signal_5970), .B1_f (new_AGEMA_signal_5971), .Z0_t (Midori_rounds_Res_Inst_mux_inst_59_U1_Y), .Z0_f (new_AGEMA_signal_6155), .Z1_t (new_AGEMA_signal_6156), .Z1_f (new_AGEMA_signal_6157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_59_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_59_U1_Y), .A0_f (new_AGEMA_signal_6155), .A1_t (new_AGEMA_signal_6156), .A1_f (new_AGEMA_signal_6157), .B0_t (Midori_rounds_mul_ResultXORkey[59]), .B0_f (new_AGEMA_signal_5640), .B1_t (new_AGEMA_signal_5641), .B1_f (new_AGEMA_signal_5642), .Z0_t (Midori_rounds_round_Result[59]), .Z0_f (new_AGEMA_signal_6341), .Z1_t (new_AGEMA_signal_6342), .Z1_f (new_AGEMA_signal_6343) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_60_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[60]), .A0_f (new_AGEMA_signal_6821), .A1_t (new_AGEMA_signal_6822), .A1_f (new_AGEMA_signal_6823), .B0_t (Midori_rounds_SR_Inv_Result[60]), .B0_f (new_AGEMA_signal_6797), .B1_t (new_AGEMA_signal_6798), .B1_f (new_AGEMA_signal_6799), .Z0_t (Midori_rounds_Res_Inst_mux_inst_60_U1_X), .Z0_f (new_AGEMA_signal_6911), .Z1_t (new_AGEMA_signal_6912), .Z1_f (new_AGEMA_signal_6913) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_60_U1_X), .B0_f (new_AGEMA_signal_6911), .B1_t (new_AGEMA_signal_6912), .B1_f (new_AGEMA_signal_6913), .Z0_t (Midori_rounds_Res_Inst_mux_inst_60_U1_Y), .Z0_f (new_AGEMA_signal_6959), .Z1_t (new_AGEMA_signal_6960), .Z1_f (new_AGEMA_signal_6961) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_60_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_60_U1_Y), .A0_f (new_AGEMA_signal_6959), .A1_t (new_AGEMA_signal_6960), .A1_f (new_AGEMA_signal_6961), .B0_t (Midori_rounds_mul_ResultXORkey[60]), .B0_f (new_AGEMA_signal_6821), .B1_t (new_AGEMA_signal_6822), .B1_f (new_AGEMA_signal_6823), .Z0_t (Midori_rounds_round_Result[60]), .Z0_f (new_AGEMA_signal_7007), .Z1_t (new_AGEMA_signal_7008), .Z1_f (new_AGEMA_signal_7009) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_61_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[61]), .A0_f (new_AGEMA_signal_5637), .A1_t (new_AGEMA_signal_5638), .A1_f (new_AGEMA_signal_5639), .B0_t (Midori_rounds_SR_Inv_Result[61]), .B0_f (new_AGEMA_signal_5499), .B1_t (new_AGEMA_signal_5500), .B1_f (new_AGEMA_signal_5501), .Z0_t (Midori_rounds_Res_Inst_mux_inst_61_U1_X), .Z0_f (new_AGEMA_signal_5972), .Z1_t (new_AGEMA_signal_5973), .Z1_f (new_AGEMA_signal_5974) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_61_U1_X), .B0_f (new_AGEMA_signal_5972), .B1_t (new_AGEMA_signal_5973), .B1_f (new_AGEMA_signal_5974), .Z0_t (Midori_rounds_Res_Inst_mux_inst_61_U1_Y), .Z0_f (new_AGEMA_signal_6158), .Z1_t (new_AGEMA_signal_6159), .Z1_f (new_AGEMA_signal_6160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_61_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_61_U1_Y), .A0_f (new_AGEMA_signal_6158), .A1_t (new_AGEMA_signal_6159), .A1_f (new_AGEMA_signal_6160), .B0_t (Midori_rounds_mul_ResultXORkey[61]), .B0_f (new_AGEMA_signal_5637), .B1_t (new_AGEMA_signal_5638), .B1_f (new_AGEMA_signal_5639), .Z0_t (Midori_rounds_round_Result[61]), .Z0_f (new_AGEMA_signal_6344), .Z1_t (new_AGEMA_signal_6345), .Z1_f (new_AGEMA_signal_6346) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_62_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[62]), .A0_f (new_AGEMA_signal_5815), .A1_t (new_AGEMA_signal_5816), .A1_f (new_AGEMA_signal_5817), .B0_t (Midori_rounds_SR_Inv_Result[62]), .B0_f (new_AGEMA_signal_5740), .B1_t (new_AGEMA_signal_5741), .B1_f (new_AGEMA_signal_5742), .Z0_t (Midori_rounds_Res_Inst_mux_inst_62_U1_X), .Z0_f (new_AGEMA_signal_6161), .Z1_t (new_AGEMA_signal_6162), .Z1_f (new_AGEMA_signal_6163) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_62_U1_X), .B0_f (new_AGEMA_signal_6161), .B1_t (new_AGEMA_signal_6162), .B1_f (new_AGEMA_signal_6163), .Z0_t (Midori_rounds_Res_Inst_mux_inst_62_U1_Y), .Z0_f (new_AGEMA_signal_6347), .Z1_t (new_AGEMA_signal_6348), .Z1_f (new_AGEMA_signal_6349) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_62_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_62_U1_Y), .A0_f (new_AGEMA_signal_6347), .A1_t (new_AGEMA_signal_6348), .A1_f (new_AGEMA_signal_6349), .B0_t (Midori_rounds_mul_ResultXORkey[62]), .B0_f (new_AGEMA_signal_5815), .B1_t (new_AGEMA_signal_5816), .B1_f (new_AGEMA_signal_5817), .Z0_t (Midori_rounds_round_Result[62]), .Z0_f (new_AGEMA_signal_6530), .Z1_t (new_AGEMA_signal_6531), .Z1_f (new_AGEMA_signal_6532) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_63_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[63]), .A0_f (new_AGEMA_signal_5634), .A1_t (new_AGEMA_signal_5635), .A1_f (new_AGEMA_signal_5636), .B0_t (Midori_rounds_SR_Inv_Result[63]), .B0_f (new_AGEMA_signal_5484), .B1_t (new_AGEMA_signal_5485), .B1_f (new_AGEMA_signal_5486), .Z0_t (Midori_rounds_Res_Inst_mux_inst_63_U1_X), .Z0_f (new_AGEMA_signal_5975), .Z1_t (new_AGEMA_signal_5976), .Z1_f (new_AGEMA_signal_5977) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enc_dec_t), .A1_f (enc_dec_f), .B0_t (Midori_rounds_Res_Inst_mux_inst_63_U1_X), .B0_f (new_AGEMA_signal_5975), .B1_t (new_AGEMA_signal_5976), .B1_f (new_AGEMA_signal_5977), .Z0_t (Midori_rounds_Res_Inst_mux_inst_63_U1_Y), .Z0_f (new_AGEMA_signal_6164), .Z1_t (new_AGEMA_signal_6165), .Z1_f (new_AGEMA_signal_6166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_63_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_63_U1_Y), .A0_f (new_AGEMA_signal_6164), .A1_t (new_AGEMA_signal_6165), .A1_f (new_AGEMA_signal_6166), .B0_t (Midori_rounds_mul_ResultXORkey[63]), .B0_f (new_AGEMA_signal_5634), .B1_t (new_AGEMA_signal_5635), .B1_f (new_AGEMA_signal_5636), .Z0_t (Midori_rounds_round_Result[63]), .Z0_f (new_AGEMA_signal_6350), .Z1_t (new_AGEMA_signal_6351), .Z1_f (new_AGEMA_signal_6352) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_1804 ( .A0_t (controller_roundCounter_N7), .A0_f (new_AGEMA_signal_2591), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (round_Signal[0]), .Z0_f (new_AGEMA_signal_2582) ) ;

    /* register cells */
endmodule
