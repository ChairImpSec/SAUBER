/* modified netlist. Source: module AES in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/5-AES_EncRoundBased_PortParallel/4-AGEMA/AES.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module AES_SAUBER_Pipeline_d1 (plaintext, key, start, ciphertext, done);
    input [127:0] plaintext ;
    input [127:0] key ;
    input start ;
    output [127:0] ciphertext ;
    output done ;
    wire n283 ;
    wire n285 ;
    wire n577 ;
    wire n585 ;
    wire n586 ;
    wire n588 ;
    wire n589 ;
    wire n591 ;
    wire n592 ;
    wire n593 ;
    wire n594 ;
    wire n595 ;
    wire n596 ;
    wire n597 ;
    wire n598 ;
    wire n599 ;
    wire n600 ;
    wire n601 ;
    wire n602 ;
    wire n603 ;
    wire n604 ;
    wire n605 ;
    wire n606 ;
    wire n607 ;
    wire n608 ;
    wire n609 ;
    wire n610 ;
    wire n611 ;
    wire n612 ;
    wire n613 ;
    wire n614 ;
    wire n615 ;
    wire n616 ;
    wire n617 ;
    wire n618 ;
    wire n619 ;
    wire n620 ;
    wire n621 ;
    wire n622 ;
    wire n623 ;
    wire n624 ;
    wire n625 ;
    wire n626 ;
    wire n627 ;
    wire n628 ;
    wire n629 ;
    wire n630 ;
    wire n631 ;
    wire n632 ;
    wire n633 ;
    wire n634 ;
    wire n635 ;
    wire n636 ;
    wire n637 ;
    wire n638 ;
    wire n639 ;
    wire n640 ;
    wire n641 ;
    wire n642 ;
    wire n643 ;
    wire n644 ;
    wire n645 ;
    wire n646 ;
    wire n647 ;
    wire n648 ;
    wire n649 ;
    wire n650 ;
    wire n651 ;
    wire n652 ;
    wire n653 ;
    wire n654 ;
    wire n655 ;
    wire n656 ;
    wire n657 ;
    wire n658 ;
    wire n659 ;
    wire n660 ;
    wire n661 ;
    wire n662 ;
    wire n663 ;
    wire n664 ;
    wire n665 ;
    wire n666 ;
    wire n667 ;
    wire n668 ;
    wire n669 ;
    wire n670 ;
    wire n671 ;
    wire n672 ;
    wire n673 ;
    wire n674 ;
    wire n675 ;
    wire n676 ;
    wire n677 ;
    wire n678 ;
    wire n679 ;
    wire n680 ;
    wire n681 ;
    wire n682 ;
    wire n683 ;
    wire n684 ;
    wire n685 ;
    wire n686 ;
    wire n687 ;
    wire n688 ;
    wire n689 ;
    wire n690 ;
    wire n691 ;
    wire n692 ;
    wire n693 ;
    wire n694 ;
    wire n695 ;
    wire n696 ;
    wire n697 ;
    wire n698 ;
    wire n699 ;
    wire n700 ;
    wire n701 ;
    wire n702 ;
    wire n703 ;
    wire n704 ;
    wire n705 ;
    wire n706 ;
    wire n707 ;
    wire n708 ;
    wire n709 ;
    wire n710 ;
    wire n711 ;
    wire n712 ;
    wire n713 ;
    wire n714 ;
    wire n715 ;
    wire n716 ;
    wire n717 ;
    wire n718 ;
    wire n719 ;
    wire n720 ;
    wire n721 ;
    wire n722 ;
    wire n723 ;
    wire n724 ;
    wire n725 ;
    wire n726 ;
    wire n727 ;
    wire n728 ;
    wire n729 ;
    wire n730 ;
    wire n731 ;
    wire n732 ;
    wire n733 ;
    wire n734 ;
    wire n735 ;
    wire n736 ;
    wire n737 ;
    wire n738 ;
    wire n739 ;
    wire n740 ;
    wire n741 ;
    wire n742 ;
    wire n743 ;
    wire n744 ;
    wire n745 ;
    wire n746 ;
    wire n747 ;
    wire n748 ;
    wire n749 ;
    wire n750 ;
    wire n751 ;
    wire n752 ;
    wire n753 ;
    wire n754 ;
    wire n755 ;
    wire n756 ;
    wire n757 ;
    wire n758 ;
    wire n759 ;
    wire n760 ;
    wire n761 ;
    wire n762 ;
    wire n763 ;
    wire n764 ;
    wire n765 ;
    wire n766 ;
    wire n767 ;
    wire n768 ;
    wire n769 ;
    wire n770 ;
    wire n771 ;
    wire n772 ;
    wire n773 ;
    wire n774 ;
    wire n775 ;
    wire n776 ;
    wire n777 ;
    wire n778 ;
    wire n779 ;
    wire n780 ;
    wire n781 ;
    wire n782 ;
    wire n783 ;
    wire n784 ;
    wire n785 ;
    wire n786 ;
    wire n787 ;
    wire n788 ;
    wire n789 ;
    wire n790 ;
    wire n791 ;
    wire n792 ;
    wire n793 ;
    wire n794 ;
    wire n795 ;
    wire n796 ;
    wire n797 ;
    wire n798 ;
    wire n799 ;
    wire n800 ;
    wire n801 ;
    wire n802 ;
    wire n803 ;
    wire n804 ;
    wire n805 ;
    wire n806 ;
    wire n807 ;
    wire n808 ;
    wire n809 ;
    wire n810 ;
    wire n811 ;
    wire n812 ;
    wire n813 ;
    wire n814 ;
    wire n815 ;
    wire n816 ;
    wire n817 ;
    wire n818 ;
    wire n819 ;
    wire n820 ;
    wire n821 ;
    wire n822 ;
    wire n823 ;
    wire n824 ;
    wire n825 ;
    wire n826 ;
    wire n827 ;
    wire n828 ;
    wire n829 ;
    wire n830 ;
    wire n831 ;
    wire n832 ;
    wire n833 ;
    wire n834 ;
    wire n835 ;
    wire n836 ;
    wire n837 ;
    wire n838 ;
    wire n839 ;
    wire n840 ;
    wire n841 ;
    wire n842 ;
    wire n843 ;
    wire n844 ;
    wire n845 ;
    wire n846 ;
    wire n847 ;
    wire n848 ;
    wire n849 ;
    wire n850 ;
    wire n851 ;
    wire n852 ;
    wire n853 ;
    wire n855 ;
    wire n856 ;
    wire RoundReg_Inst_ff_SDE_0_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_0_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_1_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_1_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_2_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_2_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_3_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_3_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_4_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_4_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_5_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_5_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_6_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_6_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_7_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_7_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_8_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_8_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_9_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_9_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_10_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_10_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_11_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_11_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_12_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_12_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_13_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_13_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_14_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_14_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_15_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_15_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_16_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_16_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_17_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_17_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_18_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_18_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_19_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_19_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_20_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_20_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_21_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_21_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_22_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_22_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_23_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_23_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_24_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_24_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_25_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_25_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_26_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_26_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_27_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_27_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_28_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_28_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_29_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_29_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_30_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_30_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_31_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_31_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_32_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_32_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_33_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_33_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_34_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_34_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_35_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_35_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_36_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_36_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_37_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_37_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_38_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_38_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_39_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_39_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_40_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_40_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_41_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_41_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_42_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_42_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_43_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_43_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_44_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_44_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_45_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_45_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_46_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_46_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_47_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_47_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_48_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_48_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_49_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_49_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_50_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_50_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_51_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_51_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_52_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_52_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_53_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_53_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_54_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_54_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_55_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_55_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_56_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_56_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_57_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_57_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_58_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_58_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_59_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_59_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_60_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_60_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_61_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_61_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_62_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_62_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_63_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_63_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_64_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_64_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_65_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_65_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_66_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_66_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_67_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_67_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_68_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_68_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_69_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_69_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_70_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_70_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_71_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_71_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_72_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_72_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_73_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_73_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_74_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_74_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_75_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_75_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_76_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_76_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_77_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_77_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_78_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_78_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_79_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_79_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_80_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_80_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_81_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_81_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_82_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_82_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_83_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_83_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_84_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_84_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_85_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_85_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_86_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_86_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_87_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_87_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_88_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_88_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_89_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_89_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_90_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_90_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_91_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_91_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_92_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_92_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_93_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_93_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_94_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_94_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_95_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_95_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_96_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_96_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_97_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_97_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_98_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_98_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_99_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_99_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_100_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_100_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_101_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_101_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_102_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_102_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_103_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_103_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_104_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_104_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_105_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_105_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_106_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_106_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_107_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_107_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_108_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_108_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_109_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_109_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_110_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_110_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_111_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_111_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_112_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_112_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_113_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_113_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_114_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_114_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_115_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_115_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_116_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_116_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_117_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_117_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_118_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_118_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_119_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_119_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_120_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_120_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_121_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_121_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_122_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_122_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_123_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_123_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_124_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_124_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_125_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_125_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_126_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_126_MUX_inst_X ;
    wire RoundReg_Inst_ff_SDE_127_MUX_inst_Y ;
    wire RoundReg_Inst_ff_SDE_127_MUX_inst_X ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire SubBytesIns_Inst_Sbox_4_L29 ;
    wire SubBytesIns_Inst_Sbox_4_L28 ;
    wire SubBytesIns_Inst_Sbox_4_L27 ;
    wire SubBytesIns_Inst_Sbox_4_L26 ;
    wire SubBytesIns_Inst_Sbox_4_L25 ;
    wire SubBytesIns_Inst_Sbox_4_L24 ;
    wire SubBytesIns_Inst_Sbox_4_L23 ;
    wire SubBytesIns_Inst_Sbox_4_L22 ;
    wire SubBytesIns_Inst_Sbox_4_L21 ;
    wire SubBytesIns_Inst_Sbox_4_L20 ;
    wire SubBytesIns_Inst_Sbox_4_L19 ;
    wire SubBytesIns_Inst_Sbox_4_L18 ;
    wire SubBytesIns_Inst_Sbox_4_L17 ;
    wire SubBytesIns_Inst_Sbox_4_L16 ;
    wire SubBytesIns_Inst_Sbox_4_L15 ;
    wire SubBytesIns_Inst_Sbox_4_L14 ;
    wire SubBytesIns_Inst_Sbox_4_L13 ;
    wire SubBytesIns_Inst_Sbox_4_L12 ;
    wire SubBytesIns_Inst_Sbox_4_L11 ;
    wire SubBytesIns_Inst_Sbox_4_L10 ;
    wire SubBytesIns_Inst_Sbox_4_L9 ;
    wire SubBytesIns_Inst_Sbox_4_L8 ;
    wire SubBytesIns_Inst_Sbox_4_L7 ;
    wire SubBytesIns_Inst_Sbox_4_L6 ;
    wire SubBytesIns_Inst_Sbox_4_L5 ;
    wire SubBytesIns_Inst_Sbox_4_L4 ;
    wire SubBytesIns_Inst_Sbox_4_L3 ;
    wire SubBytesIns_Inst_Sbox_4_L2 ;
    wire SubBytesIns_Inst_Sbox_4_L1 ;
    wire SubBytesIns_Inst_Sbox_4_L0 ;
    wire SubBytesIns_Inst_Sbox_4_M63 ;
    wire SubBytesIns_Inst_Sbox_4_M62 ;
    wire SubBytesIns_Inst_Sbox_4_M61 ;
    wire SubBytesIns_Inst_Sbox_4_M60 ;
    wire SubBytesIns_Inst_Sbox_4_M59 ;
    wire SubBytesIns_Inst_Sbox_4_M58 ;
    wire SubBytesIns_Inst_Sbox_4_M57 ;
    wire SubBytesIns_Inst_Sbox_4_M56 ;
    wire SubBytesIns_Inst_Sbox_4_M55 ;
    wire SubBytesIns_Inst_Sbox_4_M54 ;
    wire SubBytesIns_Inst_Sbox_4_M53 ;
    wire SubBytesIns_Inst_Sbox_4_M52 ;
    wire SubBytesIns_Inst_Sbox_4_M51 ;
    wire SubBytesIns_Inst_Sbox_4_M50 ;
    wire SubBytesIns_Inst_Sbox_4_M49 ;
    wire SubBytesIns_Inst_Sbox_4_M48 ;
    wire SubBytesIns_Inst_Sbox_4_M47 ;
    wire SubBytesIns_Inst_Sbox_4_M46 ;
    wire SubBytesIns_Inst_Sbox_4_M45 ;
    wire SubBytesIns_Inst_Sbox_4_M44 ;
    wire SubBytesIns_Inst_Sbox_4_M43 ;
    wire SubBytesIns_Inst_Sbox_4_M42 ;
    wire SubBytesIns_Inst_Sbox_4_M41 ;
    wire SubBytesIns_Inst_Sbox_4_M40 ;
    wire SubBytesIns_Inst_Sbox_4_M39 ;
    wire SubBytesIns_Inst_Sbox_4_M38 ;
    wire SubBytesIns_Inst_Sbox_4_M37 ;
    wire SubBytesIns_Inst_Sbox_4_M36 ;
    wire SubBytesIns_Inst_Sbox_4_M35 ;
    wire SubBytesIns_Inst_Sbox_4_M34 ;
    wire SubBytesIns_Inst_Sbox_4_M33 ;
    wire SubBytesIns_Inst_Sbox_4_M32 ;
    wire SubBytesIns_Inst_Sbox_4_M31 ;
    wire SubBytesIns_Inst_Sbox_4_M30 ;
    wire SubBytesIns_Inst_Sbox_4_M29 ;
    wire SubBytesIns_Inst_Sbox_4_M28 ;
    wire SubBytesIns_Inst_Sbox_4_M27 ;
    wire SubBytesIns_Inst_Sbox_4_M26 ;
    wire SubBytesIns_Inst_Sbox_4_M25 ;
    wire SubBytesIns_Inst_Sbox_4_M24 ;
    wire SubBytesIns_Inst_Sbox_4_M23 ;
    wire SubBytesIns_Inst_Sbox_4_M22 ;
    wire SubBytesIns_Inst_Sbox_4_M21 ;
    wire SubBytesIns_Inst_Sbox_4_M20 ;
    wire SubBytesIns_Inst_Sbox_4_M19 ;
    wire SubBytesIns_Inst_Sbox_4_M18 ;
    wire SubBytesIns_Inst_Sbox_4_M17 ;
    wire SubBytesIns_Inst_Sbox_4_M16 ;
    wire SubBytesIns_Inst_Sbox_4_M15 ;
    wire SubBytesIns_Inst_Sbox_4_M14 ;
    wire SubBytesIns_Inst_Sbox_4_M13 ;
    wire SubBytesIns_Inst_Sbox_4_M12 ;
    wire SubBytesIns_Inst_Sbox_4_M11 ;
    wire SubBytesIns_Inst_Sbox_4_M10 ;
    wire SubBytesIns_Inst_Sbox_4_M9 ;
    wire SubBytesIns_Inst_Sbox_4_M8 ;
    wire SubBytesIns_Inst_Sbox_4_M7 ;
    wire SubBytesIns_Inst_Sbox_4_M6 ;
    wire SubBytesIns_Inst_Sbox_4_M5 ;
    wire SubBytesIns_Inst_Sbox_4_M4 ;
    wire SubBytesIns_Inst_Sbox_4_M3 ;
    wire SubBytesIns_Inst_Sbox_4_M2 ;
    wire SubBytesIns_Inst_Sbox_4_M1 ;
    wire SubBytesIns_Inst_Sbox_4_T27 ;
    wire SubBytesIns_Inst_Sbox_4_T26 ;
    wire SubBytesIns_Inst_Sbox_4_T25 ;
    wire SubBytesIns_Inst_Sbox_4_T24 ;
    wire SubBytesIns_Inst_Sbox_4_T23 ;
    wire SubBytesIns_Inst_Sbox_4_T22 ;
    wire SubBytesIns_Inst_Sbox_4_T21 ;
    wire SubBytesIns_Inst_Sbox_4_T20 ;
    wire SubBytesIns_Inst_Sbox_4_T19 ;
    wire SubBytesIns_Inst_Sbox_4_T18 ;
    wire SubBytesIns_Inst_Sbox_4_T17 ;
    wire SubBytesIns_Inst_Sbox_4_T16 ;
    wire SubBytesIns_Inst_Sbox_4_T15 ;
    wire SubBytesIns_Inst_Sbox_4_T14 ;
    wire SubBytesIns_Inst_Sbox_4_T13 ;
    wire SubBytesIns_Inst_Sbox_4_T12 ;
    wire SubBytesIns_Inst_Sbox_4_T11 ;
    wire SubBytesIns_Inst_Sbox_4_T10 ;
    wire SubBytesIns_Inst_Sbox_4_T9 ;
    wire SubBytesIns_Inst_Sbox_4_T8 ;
    wire SubBytesIns_Inst_Sbox_4_T7 ;
    wire SubBytesIns_Inst_Sbox_4_T6 ;
    wire SubBytesIns_Inst_Sbox_4_T5 ;
    wire SubBytesIns_Inst_Sbox_4_T4 ;
    wire SubBytesIns_Inst_Sbox_4_T3 ;
    wire SubBytesIns_Inst_Sbox_4_T2 ;
    wire SubBytesIns_Inst_Sbox_4_T1 ;
    wire SubBytesIns_Inst_Sbox_5_L29 ;
    wire SubBytesIns_Inst_Sbox_5_L28 ;
    wire SubBytesIns_Inst_Sbox_5_L27 ;
    wire SubBytesIns_Inst_Sbox_5_L26 ;
    wire SubBytesIns_Inst_Sbox_5_L25 ;
    wire SubBytesIns_Inst_Sbox_5_L24 ;
    wire SubBytesIns_Inst_Sbox_5_L23 ;
    wire SubBytesIns_Inst_Sbox_5_L22 ;
    wire SubBytesIns_Inst_Sbox_5_L21 ;
    wire SubBytesIns_Inst_Sbox_5_L20 ;
    wire SubBytesIns_Inst_Sbox_5_L19 ;
    wire SubBytesIns_Inst_Sbox_5_L18 ;
    wire SubBytesIns_Inst_Sbox_5_L17 ;
    wire SubBytesIns_Inst_Sbox_5_L16 ;
    wire SubBytesIns_Inst_Sbox_5_L15 ;
    wire SubBytesIns_Inst_Sbox_5_L14 ;
    wire SubBytesIns_Inst_Sbox_5_L13 ;
    wire SubBytesIns_Inst_Sbox_5_L12 ;
    wire SubBytesIns_Inst_Sbox_5_L11 ;
    wire SubBytesIns_Inst_Sbox_5_L10 ;
    wire SubBytesIns_Inst_Sbox_5_L9 ;
    wire SubBytesIns_Inst_Sbox_5_L8 ;
    wire SubBytesIns_Inst_Sbox_5_L7 ;
    wire SubBytesIns_Inst_Sbox_5_L6 ;
    wire SubBytesIns_Inst_Sbox_5_L5 ;
    wire SubBytesIns_Inst_Sbox_5_L4 ;
    wire SubBytesIns_Inst_Sbox_5_L3 ;
    wire SubBytesIns_Inst_Sbox_5_L2 ;
    wire SubBytesIns_Inst_Sbox_5_L1 ;
    wire SubBytesIns_Inst_Sbox_5_L0 ;
    wire SubBytesIns_Inst_Sbox_5_M63 ;
    wire SubBytesIns_Inst_Sbox_5_M62 ;
    wire SubBytesIns_Inst_Sbox_5_M61 ;
    wire SubBytesIns_Inst_Sbox_5_M60 ;
    wire SubBytesIns_Inst_Sbox_5_M59 ;
    wire SubBytesIns_Inst_Sbox_5_M58 ;
    wire SubBytesIns_Inst_Sbox_5_M57 ;
    wire SubBytesIns_Inst_Sbox_5_M56 ;
    wire SubBytesIns_Inst_Sbox_5_M55 ;
    wire SubBytesIns_Inst_Sbox_5_M54 ;
    wire SubBytesIns_Inst_Sbox_5_M53 ;
    wire SubBytesIns_Inst_Sbox_5_M52 ;
    wire SubBytesIns_Inst_Sbox_5_M51 ;
    wire SubBytesIns_Inst_Sbox_5_M50 ;
    wire SubBytesIns_Inst_Sbox_5_M49 ;
    wire SubBytesIns_Inst_Sbox_5_M48 ;
    wire SubBytesIns_Inst_Sbox_5_M47 ;
    wire SubBytesIns_Inst_Sbox_5_M46 ;
    wire SubBytesIns_Inst_Sbox_5_M45 ;
    wire SubBytesIns_Inst_Sbox_5_M44 ;
    wire SubBytesIns_Inst_Sbox_5_M43 ;
    wire SubBytesIns_Inst_Sbox_5_M42 ;
    wire SubBytesIns_Inst_Sbox_5_M41 ;
    wire SubBytesIns_Inst_Sbox_5_M40 ;
    wire SubBytesIns_Inst_Sbox_5_M39 ;
    wire SubBytesIns_Inst_Sbox_5_M38 ;
    wire SubBytesIns_Inst_Sbox_5_M37 ;
    wire SubBytesIns_Inst_Sbox_5_M36 ;
    wire SubBytesIns_Inst_Sbox_5_M35 ;
    wire SubBytesIns_Inst_Sbox_5_M34 ;
    wire SubBytesIns_Inst_Sbox_5_M33 ;
    wire SubBytesIns_Inst_Sbox_5_M32 ;
    wire SubBytesIns_Inst_Sbox_5_M31 ;
    wire SubBytesIns_Inst_Sbox_5_M30 ;
    wire SubBytesIns_Inst_Sbox_5_M29 ;
    wire SubBytesIns_Inst_Sbox_5_M28 ;
    wire SubBytesIns_Inst_Sbox_5_M27 ;
    wire SubBytesIns_Inst_Sbox_5_M26 ;
    wire SubBytesIns_Inst_Sbox_5_M25 ;
    wire SubBytesIns_Inst_Sbox_5_M24 ;
    wire SubBytesIns_Inst_Sbox_5_M23 ;
    wire SubBytesIns_Inst_Sbox_5_M22 ;
    wire SubBytesIns_Inst_Sbox_5_M21 ;
    wire SubBytesIns_Inst_Sbox_5_M20 ;
    wire SubBytesIns_Inst_Sbox_5_M19 ;
    wire SubBytesIns_Inst_Sbox_5_M18 ;
    wire SubBytesIns_Inst_Sbox_5_M17 ;
    wire SubBytesIns_Inst_Sbox_5_M16 ;
    wire SubBytesIns_Inst_Sbox_5_M15 ;
    wire SubBytesIns_Inst_Sbox_5_M14 ;
    wire SubBytesIns_Inst_Sbox_5_M13 ;
    wire SubBytesIns_Inst_Sbox_5_M12 ;
    wire SubBytesIns_Inst_Sbox_5_M11 ;
    wire SubBytesIns_Inst_Sbox_5_M10 ;
    wire SubBytesIns_Inst_Sbox_5_M9 ;
    wire SubBytesIns_Inst_Sbox_5_M8 ;
    wire SubBytesIns_Inst_Sbox_5_M7 ;
    wire SubBytesIns_Inst_Sbox_5_M6 ;
    wire SubBytesIns_Inst_Sbox_5_M5 ;
    wire SubBytesIns_Inst_Sbox_5_M4 ;
    wire SubBytesIns_Inst_Sbox_5_M3 ;
    wire SubBytesIns_Inst_Sbox_5_M2 ;
    wire SubBytesIns_Inst_Sbox_5_M1 ;
    wire SubBytesIns_Inst_Sbox_5_T27 ;
    wire SubBytesIns_Inst_Sbox_5_T26 ;
    wire SubBytesIns_Inst_Sbox_5_T25 ;
    wire SubBytesIns_Inst_Sbox_5_T24 ;
    wire SubBytesIns_Inst_Sbox_5_T23 ;
    wire SubBytesIns_Inst_Sbox_5_T22 ;
    wire SubBytesIns_Inst_Sbox_5_T21 ;
    wire SubBytesIns_Inst_Sbox_5_T20 ;
    wire SubBytesIns_Inst_Sbox_5_T19 ;
    wire SubBytesIns_Inst_Sbox_5_T18 ;
    wire SubBytesIns_Inst_Sbox_5_T17 ;
    wire SubBytesIns_Inst_Sbox_5_T16 ;
    wire SubBytesIns_Inst_Sbox_5_T15 ;
    wire SubBytesIns_Inst_Sbox_5_T14 ;
    wire SubBytesIns_Inst_Sbox_5_T13 ;
    wire SubBytesIns_Inst_Sbox_5_T12 ;
    wire SubBytesIns_Inst_Sbox_5_T11 ;
    wire SubBytesIns_Inst_Sbox_5_T10 ;
    wire SubBytesIns_Inst_Sbox_5_T9 ;
    wire SubBytesIns_Inst_Sbox_5_T8 ;
    wire SubBytesIns_Inst_Sbox_5_T7 ;
    wire SubBytesIns_Inst_Sbox_5_T6 ;
    wire SubBytesIns_Inst_Sbox_5_T5 ;
    wire SubBytesIns_Inst_Sbox_5_T4 ;
    wire SubBytesIns_Inst_Sbox_5_T3 ;
    wire SubBytesIns_Inst_Sbox_5_T2 ;
    wire SubBytesIns_Inst_Sbox_5_T1 ;
    wire SubBytesIns_Inst_Sbox_6_L29 ;
    wire SubBytesIns_Inst_Sbox_6_L28 ;
    wire SubBytesIns_Inst_Sbox_6_L27 ;
    wire SubBytesIns_Inst_Sbox_6_L26 ;
    wire SubBytesIns_Inst_Sbox_6_L25 ;
    wire SubBytesIns_Inst_Sbox_6_L24 ;
    wire SubBytesIns_Inst_Sbox_6_L23 ;
    wire SubBytesIns_Inst_Sbox_6_L22 ;
    wire SubBytesIns_Inst_Sbox_6_L21 ;
    wire SubBytesIns_Inst_Sbox_6_L20 ;
    wire SubBytesIns_Inst_Sbox_6_L19 ;
    wire SubBytesIns_Inst_Sbox_6_L18 ;
    wire SubBytesIns_Inst_Sbox_6_L17 ;
    wire SubBytesIns_Inst_Sbox_6_L16 ;
    wire SubBytesIns_Inst_Sbox_6_L15 ;
    wire SubBytesIns_Inst_Sbox_6_L14 ;
    wire SubBytesIns_Inst_Sbox_6_L13 ;
    wire SubBytesIns_Inst_Sbox_6_L12 ;
    wire SubBytesIns_Inst_Sbox_6_L11 ;
    wire SubBytesIns_Inst_Sbox_6_L10 ;
    wire SubBytesIns_Inst_Sbox_6_L9 ;
    wire SubBytesIns_Inst_Sbox_6_L8 ;
    wire SubBytesIns_Inst_Sbox_6_L7 ;
    wire SubBytesIns_Inst_Sbox_6_L6 ;
    wire SubBytesIns_Inst_Sbox_6_L5 ;
    wire SubBytesIns_Inst_Sbox_6_L4 ;
    wire SubBytesIns_Inst_Sbox_6_L3 ;
    wire SubBytesIns_Inst_Sbox_6_L2 ;
    wire SubBytesIns_Inst_Sbox_6_L1 ;
    wire SubBytesIns_Inst_Sbox_6_L0 ;
    wire SubBytesIns_Inst_Sbox_6_M63 ;
    wire SubBytesIns_Inst_Sbox_6_M62 ;
    wire SubBytesIns_Inst_Sbox_6_M61 ;
    wire SubBytesIns_Inst_Sbox_6_M60 ;
    wire SubBytesIns_Inst_Sbox_6_M59 ;
    wire SubBytesIns_Inst_Sbox_6_M58 ;
    wire SubBytesIns_Inst_Sbox_6_M57 ;
    wire SubBytesIns_Inst_Sbox_6_M56 ;
    wire SubBytesIns_Inst_Sbox_6_M55 ;
    wire SubBytesIns_Inst_Sbox_6_M54 ;
    wire SubBytesIns_Inst_Sbox_6_M53 ;
    wire SubBytesIns_Inst_Sbox_6_M52 ;
    wire SubBytesIns_Inst_Sbox_6_M51 ;
    wire SubBytesIns_Inst_Sbox_6_M50 ;
    wire SubBytesIns_Inst_Sbox_6_M49 ;
    wire SubBytesIns_Inst_Sbox_6_M48 ;
    wire SubBytesIns_Inst_Sbox_6_M47 ;
    wire SubBytesIns_Inst_Sbox_6_M46 ;
    wire SubBytesIns_Inst_Sbox_6_M45 ;
    wire SubBytesIns_Inst_Sbox_6_M44 ;
    wire SubBytesIns_Inst_Sbox_6_M43 ;
    wire SubBytesIns_Inst_Sbox_6_M42 ;
    wire SubBytesIns_Inst_Sbox_6_M41 ;
    wire SubBytesIns_Inst_Sbox_6_M40 ;
    wire SubBytesIns_Inst_Sbox_6_M39 ;
    wire SubBytesIns_Inst_Sbox_6_M38 ;
    wire SubBytesIns_Inst_Sbox_6_M37 ;
    wire SubBytesIns_Inst_Sbox_6_M36 ;
    wire SubBytesIns_Inst_Sbox_6_M35 ;
    wire SubBytesIns_Inst_Sbox_6_M34 ;
    wire SubBytesIns_Inst_Sbox_6_M33 ;
    wire SubBytesIns_Inst_Sbox_6_M32 ;
    wire SubBytesIns_Inst_Sbox_6_M31 ;
    wire SubBytesIns_Inst_Sbox_6_M30 ;
    wire SubBytesIns_Inst_Sbox_6_M29 ;
    wire SubBytesIns_Inst_Sbox_6_M28 ;
    wire SubBytesIns_Inst_Sbox_6_M27 ;
    wire SubBytesIns_Inst_Sbox_6_M26 ;
    wire SubBytesIns_Inst_Sbox_6_M25 ;
    wire SubBytesIns_Inst_Sbox_6_M24 ;
    wire SubBytesIns_Inst_Sbox_6_M23 ;
    wire SubBytesIns_Inst_Sbox_6_M22 ;
    wire SubBytesIns_Inst_Sbox_6_M21 ;
    wire SubBytesIns_Inst_Sbox_6_M20 ;
    wire SubBytesIns_Inst_Sbox_6_M19 ;
    wire SubBytesIns_Inst_Sbox_6_M18 ;
    wire SubBytesIns_Inst_Sbox_6_M17 ;
    wire SubBytesIns_Inst_Sbox_6_M16 ;
    wire SubBytesIns_Inst_Sbox_6_M15 ;
    wire SubBytesIns_Inst_Sbox_6_M14 ;
    wire SubBytesIns_Inst_Sbox_6_M13 ;
    wire SubBytesIns_Inst_Sbox_6_M12 ;
    wire SubBytesIns_Inst_Sbox_6_M11 ;
    wire SubBytesIns_Inst_Sbox_6_M10 ;
    wire SubBytesIns_Inst_Sbox_6_M9 ;
    wire SubBytesIns_Inst_Sbox_6_M8 ;
    wire SubBytesIns_Inst_Sbox_6_M7 ;
    wire SubBytesIns_Inst_Sbox_6_M6 ;
    wire SubBytesIns_Inst_Sbox_6_M5 ;
    wire SubBytesIns_Inst_Sbox_6_M4 ;
    wire SubBytesIns_Inst_Sbox_6_M3 ;
    wire SubBytesIns_Inst_Sbox_6_M2 ;
    wire SubBytesIns_Inst_Sbox_6_M1 ;
    wire SubBytesIns_Inst_Sbox_6_T27 ;
    wire SubBytesIns_Inst_Sbox_6_T26 ;
    wire SubBytesIns_Inst_Sbox_6_T25 ;
    wire SubBytesIns_Inst_Sbox_6_T24 ;
    wire SubBytesIns_Inst_Sbox_6_T23 ;
    wire SubBytesIns_Inst_Sbox_6_T22 ;
    wire SubBytesIns_Inst_Sbox_6_T21 ;
    wire SubBytesIns_Inst_Sbox_6_T20 ;
    wire SubBytesIns_Inst_Sbox_6_T19 ;
    wire SubBytesIns_Inst_Sbox_6_T18 ;
    wire SubBytesIns_Inst_Sbox_6_T17 ;
    wire SubBytesIns_Inst_Sbox_6_T16 ;
    wire SubBytesIns_Inst_Sbox_6_T15 ;
    wire SubBytesIns_Inst_Sbox_6_T14 ;
    wire SubBytesIns_Inst_Sbox_6_T13 ;
    wire SubBytesIns_Inst_Sbox_6_T12 ;
    wire SubBytesIns_Inst_Sbox_6_T11 ;
    wire SubBytesIns_Inst_Sbox_6_T10 ;
    wire SubBytesIns_Inst_Sbox_6_T9 ;
    wire SubBytesIns_Inst_Sbox_6_T8 ;
    wire SubBytesIns_Inst_Sbox_6_T7 ;
    wire SubBytesIns_Inst_Sbox_6_T6 ;
    wire SubBytesIns_Inst_Sbox_6_T5 ;
    wire SubBytesIns_Inst_Sbox_6_T4 ;
    wire SubBytesIns_Inst_Sbox_6_T3 ;
    wire SubBytesIns_Inst_Sbox_6_T2 ;
    wire SubBytesIns_Inst_Sbox_6_T1 ;
    wire SubBytesIns_Inst_Sbox_7_L29 ;
    wire SubBytesIns_Inst_Sbox_7_L28 ;
    wire SubBytesIns_Inst_Sbox_7_L27 ;
    wire SubBytesIns_Inst_Sbox_7_L26 ;
    wire SubBytesIns_Inst_Sbox_7_L25 ;
    wire SubBytesIns_Inst_Sbox_7_L24 ;
    wire SubBytesIns_Inst_Sbox_7_L23 ;
    wire SubBytesIns_Inst_Sbox_7_L22 ;
    wire SubBytesIns_Inst_Sbox_7_L21 ;
    wire SubBytesIns_Inst_Sbox_7_L20 ;
    wire SubBytesIns_Inst_Sbox_7_L19 ;
    wire SubBytesIns_Inst_Sbox_7_L18 ;
    wire SubBytesIns_Inst_Sbox_7_L17 ;
    wire SubBytesIns_Inst_Sbox_7_L16 ;
    wire SubBytesIns_Inst_Sbox_7_L15 ;
    wire SubBytesIns_Inst_Sbox_7_L14 ;
    wire SubBytesIns_Inst_Sbox_7_L13 ;
    wire SubBytesIns_Inst_Sbox_7_L12 ;
    wire SubBytesIns_Inst_Sbox_7_L11 ;
    wire SubBytesIns_Inst_Sbox_7_L10 ;
    wire SubBytesIns_Inst_Sbox_7_L9 ;
    wire SubBytesIns_Inst_Sbox_7_L8 ;
    wire SubBytesIns_Inst_Sbox_7_L7 ;
    wire SubBytesIns_Inst_Sbox_7_L6 ;
    wire SubBytesIns_Inst_Sbox_7_L5 ;
    wire SubBytesIns_Inst_Sbox_7_L4 ;
    wire SubBytesIns_Inst_Sbox_7_L3 ;
    wire SubBytesIns_Inst_Sbox_7_L2 ;
    wire SubBytesIns_Inst_Sbox_7_L1 ;
    wire SubBytesIns_Inst_Sbox_7_L0 ;
    wire SubBytesIns_Inst_Sbox_7_M63 ;
    wire SubBytesIns_Inst_Sbox_7_M62 ;
    wire SubBytesIns_Inst_Sbox_7_M61 ;
    wire SubBytesIns_Inst_Sbox_7_M60 ;
    wire SubBytesIns_Inst_Sbox_7_M59 ;
    wire SubBytesIns_Inst_Sbox_7_M58 ;
    wire SubBytesIns_Inst_Sbox_7_M57 ;
    wire SubBytesIns_Inst_Sbox_7_M56 ;
    wire SubBytesIns_Inst_Sbox_7_M55 ;
    wire SubBytesIns_Inst_Sbox_7_M54 ;
    wire SubBytesIns_Inst_Sbox_7_M53 ;
    wire SubBytesIns_Inst_Sbox_7_M52 ;
    wire SubBytesIns_Inst_Sbox_7_M51 ;
    wire SubBytesIns_Inst_Sbox_7_M50 ;
    wire SubBytesIns_Inst_Sbox_7_M49 ;
    wire SubBytesIns_Inst_Sbox_7_M48 ;
    wire SubBytesIns_Inst_Sbox_7_M47 ;
    wire SubBytesIns_Inst_Sbox_7_M46 ;
    wire SubBytesIns_Inst_Sbox_7_M45 ;
    wire SubBytesIns_Inst_Sbox_7_M44 ;
    wire SubBytesIns_Inst_Sbox_7_M43 ;
    wire SubBytesIns_Inst_Sbox_7_M42 ;
    wire SubBytesIns_Inst_Sbox_7_M41 ;
    wire SubBytesIns_Inst_Sbox_7_M40 ;
    wire SubBytesIns_Inst_Sbox_7_M39 ;
    wire SubBytesIns_Inst_Sbox_7_M38 ;
    wire SubBytesIns_Inst_Sbox_7_M37 ;
    wire SubBytesIns_Inst_Sbox_7_M36 ;
    wire SubBytesIns_Inst_Sbox_7_M35 ;
    wire SubBytesIns_Inst_Sbox_7_M34 ;
    wire SubBytesIns_Inst_Sbox_7_M33 ;
    wire SubBytesIns_Inst_Sbox_7_M32 ;
    wire SubBytesIns_Inst_Sbox_7_M31 ;
    wire SubBytesIns_Inst_Sbox_7_M30 ;
    wire SubBytesIns_Inst_Sbox_7_M29 ;
    wire SubBytesIns_Inst_Sbox_7_M28 ;
    wire SubBytesIns_Inst_Sbox_7_M27 ;
    wire SubBytesIns_Inst_Sbox_7_M26 ;
    wire SubBytesIns_Inst_Sbox_7_M25 ;
    wire SubBytesIns_Inst_Sbox_7_M24 ;
    wire SubBytesIns_Inst_Sbox_7_M23 ;
    wire SubBytesIns_Inst_Sbox_7_M22 ;
    wire SubBytesIns_Inst_Sbox_7_M21 ;
    wire SubBytesIns_Inst_Sbox_7_M20 ;
    wire SubBytesIns_Inst_Sbox_7_M19 ;
    wire SubBytesIns_Inst_Sbox_7_M18 ;
    wire SubBytesIns_Inst_Sbox_7_M17 ;
    wire SubBytesIns_Inst_Sbox_7_M16 ;
    wire SubBytesIns_Inst_Sbox_7_M15 ;
    wire SubBytesIns_Inst_Sbox_7_M14 ;
    wire SubBytesIns_Inst_Sbox_7_M13 ;
    wire SubBytesIns_Inst_Sbox_7_M12 ;
    wire SubBytesIns_Inst_Sbox_7_M11 ;
    wire SubBytesIns_Inst_Sbox_7_M10 ;
    wire SubBytesIns_Inst_Sbox_7_M9 ;
    wire SubBytesIns_Inst_Sbox_7_M8 ;
    wire SubBytesIns_Inst_Sbox_7_M7 ;
    wire SubBytesIns_Inst_Sbox_7_M6 ;
    wire SubBytesIns_Inst_Sbox_7_M5 ;
    wire SubBytesIns_Inst_Sbox_7_M4 ;
    wire SubBytesIns_Inst_Sbox_7_M3 ;
    wire SubBytesIns_Inst_Sbox_7_M2 ;
    wire SubBytesIns_Inst_Sbox_7_M1 ;
    wire SubBytesIns_Inst_Sbox_7_T27 ;
    wire SubBytesIns_Inst_Sbox_7_T26 ;
    wire SubBytesIns_Inst_Sbox_7_T25 ;
    wire SubBytesIns_Inst_Sbox_7_T24 ;
    wire SubBytesIns_Inst_Sbox_7_T23 ;
    wire SubBytesIns_Inst_Sbox_7_T22 ;
    wire SubBytesIns_Inst_Sbox_7_T21 ;
    wire SubBytesIns_Inst_Sbox_7_T20 ;
    wire SubBytesIns_Inst_Sbox_7_T19 ;
    wire SubBytesIns_Inst_Sbox_7_T18 ;
    wire SubBytesIns_Inst_Sbox_7_T17 ;
    wire SubBytesIns_Inst_Sbox_7_T16 ;
    wire SubBytesIns_Inst_Sbox_7_T15 ;
    wire SubBytesIns_Inst_Sbox_7_T14 ;
    wire SubBytesIns_Inst_Sbox_7_T13 ;
    wire SubBytesIns_Inst_Sbox_7_T12 ;
    wire SubBytesIns_Inst_Sbox_7_T11 ;
    wire SubBytesIns_Inst_Sbox_7_T10 ;
    wire SubBytesIns_Inst_Sbox_7_T9 ;
    wire SubBytesIns_Inst_Sbox_7_T8 ;
    wire SubBytesIns_Inst_Sbox_7_T7 ;
    wire SubBytesIns_Inst_Sbox_7_T6 ;
    wire SubBytesIns_Inst_Sbox_7_T5 ;
    wire SubBytesIns_Inst_Sbox_7_T4 ;
    wire SubBytesIns_Inst_Sbox_7_T3 ;
    wire SubBytesIns_Inst_Sbox_7_T2 ;
    wire SubBytesIns_Inst_Sbox_7_T1 ;
    wire SubBytesIns_Inst_Sbox_8_L29 ;
    wire SubBytesIns_Inst_Sbox_8_L28 ;
    wire SubBytesIns_Inst_Sbox_8_L27 ;
    wire SubBytesIns_Inst_Sbox_8_L26 ;
    wire SubBytesIns_Inst_Sbox_8_L25 ;
    wire SubBytesIns_Inst_Sbox_8_L24 ;
    wire SubBytesIns_Inst_Sbox_8_L23 ;
    wire SubBytesIns_Inst_Sbox_8_L22 ;
    wire SubBytesIns_Inst_Sbox_8_L21 ;
    wire SubBytesIns_Inst_Sbox_8_L20 ;
    wire SubBytesIns_Inst_Sbox_8_L19 ;
    wire SubBytesIns_Inst_Sbox_8_L18 ;
    wire SubBytesIns_Inst_Sbox_8_L17 ;
    wire SubBytesIns_Inst_Sbox_8_L16 ;
    wire SubBytesIns_Inst_Sbox_8_L15 ;
    wire SubBytesIns_Inst_Sbox_8_L14 ;
    wire SubBytesIns_Inst_Sbox_8_L13 ;
    wire SubBytesIns_Inst_Sbox_8_L12 ;
    wire SubBytesIns_Inst_Sbox_8_L11 ;
    wire SubBytesIns_Inst_Sbox_8_L10 ;
    wire SubBytesIns_Inst_Sbox_8_L9 ;
    wire SubBytesIns_Inst_Sbox_8_L8 ;
    wire SubBytesIns_Inst_Sbox_8_L7 ;
    wire SubBytesIns_Inst_Sbox_8_L6 ;
    wire SubBytesIns_Inst_Sbox_8_L5 ;
    wire SubBytesIns_Inst_Sbox_8_L4 ;
    wire SubBytesIns_Inst_Sbox_8_L3 ;
    wire SubBytesIns_Inst_Sbox_8_L2 ;
    wire SubBytesIns_Inst_Sbox_8_L1 ;
    wire SubBytesIns_Inst_Sbox_8_L0 ;
    wire SubBytesIns_Inst_Sbox_8_M63 ;
    wire SubBytesIns_Inst_Sbox_8_M62 ;
    wire SubBytesIns_Inst_Sbox_8_M61 ;
    wire SubBytesIns_Inst_Sbox_8_M60 ;
    wire SubBytesIns_Inst_Sbox_8_M59 ;
    wire SubBytesIns_Inst_Sbox_8_M58 ;
    wire SubBytesIns_Inst_Sbox_8_M57 ;
    wire SubBytesIns_Inst_Sbox_8_M56 ;
    wire SubBytesIns_Inst_Sbox_8_M55 ;
    wire SubBytesIns_Inst_Sbox_8_M54 ;
    wire SubBytesIns_Inst_Sbox_8_M53 ;
    wire SubBytesIns_Inst_Sbox_8_M52 ;
    wire SubBytesIns_Inst_Sbox_8_M51 ;
    wire SubBytesIns_Inst_Sbox_8_M50 ;
    wire SubBytesIns_Inst_Sbox_8_M49 ;
    wire SubBytesIns_Inst_Sbox_8_M48 ;
    wire SubBytesIns_Inst_Sbox_8_M47 ;
    wire SubBytesIns_Inst_Sbox_8_M46 ;
    wire SubBytesIns_Inst_Sbox_8_M45 ;
    wire SubBytesIns_Inst_Sbox_8_M44 ;
    wire SubBytesIns_Inst_Sbox_8_M43 ;
    wire SubBytesIns_Inst_Sbox_8_M42 ;
    wire SubBytesIns_Inst_Sbox_8_M41 ;
    wire SubBytesIns_Inst_Sbox_8_M40 ;
    wire SubBytesIns_Inst_Sbox_8_M39 ;
    wire SubBytesIns_Inst_Sbox_8_M38 ;
    wire SubBytesIns_Inst_Sbox_8_M37 ;
    wire SubBytesIns_Inst_Sbox_8_M36 ;
    wire SubBytesIns_Inst_Sbox_8_M35 ;
    wire SubBytesIns_Inst_Sbox_8_M34 ;
    wire SubBytesIns_Inst_Sbox_8_M33 ;
    wire SubBytesIns_Inst_Sbox_8_M32 ;
    wire SubBytesIns_Inst_Sbox_8_M31 ;
    wire SubBytesIns_Inst_Sbox_8_M30 ;
    wire SubBytesIns_Inst_Sbox_8_M29 ;
    wire SubBytesIns_Inst_Sbox_8_M28 ;
    wire SubBytesIns_Inst_Sbox_8_M27 ;
    wire SubBytesIns_Inst_Sbox_8_M26 ;
    wire SubBytesIns_Inst_Sbox_8_M25 ;
    wire SubBytesIns_Inst_Sbox_8_M24 ;
    wire SubBytesIns_Inst_Sbox_8_M23 ;
    wire SubBytesIns_Inst_Sbox_8_M22 ;
    wire SubBytesIns_Inst_Sbox_8_M21 ;
    wire SubBytesIns_Inst_Sbox_8_M20 ;
    wire SubBytesIns_Inst_Sbox_8_M19 ;
    wire SubBytesIns_Inst_Sbox_8_M18 ;
    wire SubBytesIns_Inst_Sbox_8_M17 ;
    wire SubBytesIns_Inst_Sbox_8_M16 ;
    wire SubBytesIns_Inst_Sbox_8_M15 ;
    wire SubBytesIns_Inst_Sbox_8_M14 ;
    wire SubBytesIns_Inst_Sbox_8_M13 ;
    wire SubBytesIns_Inst_Sbox_8_M12 ;
    wire SubBytesIns_Inst_Sbox_8_M11 ;
    wire SubBytesIns_Inst_Sbox_8_M10 ;
    wire SubBytesIns_Inst_Sbox_8_M9 ;
    wire SubBytesIns_Inst_Sbox_8_M8 ;
    wire SubBytesIns_Inst_Sbox_8_M7 ;
    wire SubBytesIns_Inst_Sbox_8_M6 ;
    wire SubBytesIns_Inst_Sbox_8_M5 ;
    wire SubBytesIns_Inst_Sbox_8_M4 ;
    wire SubBytesIns_Inst_Sbox_8_M3 ;
    wire SubBytesIns_Inst_Sbox_8_M2 ;
    wire SubBytesIns_Inst_Sbox_8_M1 ;
    wire SubBytesIns_Inst_Sbox_8_T27 ;
    wire SubBytesIns_Inst_Sbox_8_T26 ;
    wire SubBytesIns_Inst_Sbox_8_T25 ;
    wire SubBytesIns_Inst_Sbox_8_T24 ;
    wire SubBytesIns_Inst_Sbox_8_T23 ;
    wire SubBytesIns_Inst_Sbox_8_T22 ;
    wire SubBytesIns_Inst_Sbox_8_T21 ;
    wire SubBytesIns_Inst_Sbox_8_T20 ;
    wire SubBytesIns_Inst_Sbox_8_T19 ;
    wire SubBytesIns_Inst_Sbox_8_T18 ;
    wire SubBytesIns_Inst_Sbox_8_T17 ;
    wire SubBytesIns_Inst_Sbox_8_T16 ;
    wire SubBytesIns_Inst_Sbox_8_T15 ;
    wire SubBytesIns_Inst_Sbox_8_T14 ;
    wire SubBytesIns_Inst_Sbox_8_T13 ;
    wire SubBytesIns_Inst_Sbox_8_T12 ;
    wire SubBytesIns_Inst_Sbox_8_T11 ;
    wire SubBytesIns_Inst_Sbox_8_T10 ;
    wire SubBytesIns_Inst_Sbox_8_T9 ;
    wire SubBytesIns_Inst_Sbox_8_T8 ;
    wire SubBytesIns_Inst_Sbox_8_T7 ;
    wire SubBytesIns_Inst_Sbox_8_T6 ;
    wire SubBytesIns_Inst_Sbox_8_T5 ;
    wire SubBytesIns_Inst_Sbox_8_T4 ;
    wire SubBytesIns_Inst_Sbox_8_T3 ;
    wire SubBytesIns_Inst_Sbox_8_T2 ;
    wire SubBytesIns_Inst_Sbox_8_T1 ;
    wire SubBytesIns_Inst_Sbox_9_L29 ;
    wire SubBytesIns_Inst_Sbox_9_L28 ;
    wire SubBytesIns_Inst_Sbox_9_L27 ;
    wire SubBytesIns_Inst_Sbox_9_L26 ;
    wire SubBytesIns_Inst_Sbox_9_L25 ;
    wire SubBytesIns_Inst_Sbox_9_L24 ;
    wire SubBytesIns_Inst_Sbox_9_L23 ;
    wire SubBytesIns_Inst_Sbox_9_L22 ;
    wire SubBytesIns_Inst_Sbox_9_L21 ;
    wire SubBytesIns_Inst_Sbox_9_L20 ;
    wire SubBytesIns_Inst_Sbox_9_L19 ;
    wire SubBytesIns_Inst_Sbox_9_L18 ;
    wire SubBytesIns_Inst_Sbox_9_L17 ;
    wire SubBytesIns_Inst_Sbox_9_L16 ;
    wire SubBytesIns_Inst_Sbox_9_L15 ;
    wire SubBytesIns_Inst_Sbox_9_L14 ;
    wire SubBytesIns_Inst_Sbox_9_L13 ;
    wire SubBytesIns_Inst_Sbox_9_L12 ;
    wire SubBytesIns_Inst_Sbox_9_L11 ;
    wire SubBytesIns_Inst_Sbox_9_L10 ;
    wire SubBytesIns_Inst_Sbox_9_L9 ;
    wire SubBytesIns_Inst_Sbox_9_L8 ;
    wire SubBytesIns_Inst_Sbox_9_L7 ;
    wire SubBytesIns_Inst_Sbox_9_L6 ;
    wire SubBytesIns_Inst_Sbox_9_L5 ;
    wire SubBytesIns_Inst_Sbox_9_L4 ;
    wire SubBytesIns_Inst_Sbox_9_L3 ;
    wire SubBytesIns_Inst_Sbox_9_L2 ;
    wire SubBytesIns_Inst_Sbox_9_L1 ;
    wire SubBytesIns_Inst_Sbox_9_L0 ;
    wire SubBytesIns_Inst_Sbox_9_M63 ;
    wire SubBytesIns_Inst_Sbox_9_M62 ;
    wire SubBytesIns_Inst_Sbox_9_M61 ;
    wire SubBytesIns_Inst_Sbox_9_M60 ;
    wire SubBytesIns_Inst_Sbox_9_M59 ;
    wire SubBytesIns_Inst_Sbox_9_M58 ;
    wire SubBytesIns_Inst_Sbox_9_M57 ;
    wire SubBytesIns_Inst_Sbox_9_M56 ;
    wire SubBytesIns_Inst_Sbox_9_M55 ;
    wire SubBytesIns_Inst_Sbox_9_M54 ;
    wire SubBytesIns_Inst_Sbox_9_M53 ;
    wire SubBytesIns_Inst_Sbox_9_M52 ;
    wire SubBytesIns_Inst_Sbox_9_M51 ;
    wire SubBytesIns_Inst_Sbox_9_M50 ;
    wire SubBytesIns_Inst_Sbox_9_M49 ;
    wire SubBytesIns_Inst_Sbox_9_M48 ;
    wire SubBytesIns_Inst_Sbox_9_M47 ;
    wire SubBytesIns_Inst_Sbox_9_M46 ;
    wire SubBytesIns_Inst_Sbox_9_M45 ;
    wire SubBytesIns_Inst_Sbox_9_M44 ;
    wire SubBytesIns_Inst_Sbox_9_M43 ;
    wire SubBytesIns_Inst_Sbox_9_M42 ;
    wire SubBytesIns_Inst_Sbox_9_M41 ;
    wire SubBytesIns_Inst_Sbox_9_M40 ;
    wire SubBytesIns_Inst_Sbox_9_M39 ;
    wire SubBytesIns_Inst_Sbox_9_M38 ;
    wire SubBytesIns_Inst_Sbox_9_M37 ;
    wire SubBytesIns_Inst_Sbox_9_M36 ;
    wire SubBytesIns_Inst_Sbox_9_M35 ;
    wire SubBytesIns_Inst_Sbox_9_M34 ;
    wire SubBytesIns_Inst_Sbox_9_M33 ;
    wire SubBytesIns_Inst_Sbox_9_M32 ;
    wire SubBytesIns_Inst_Sbox_9_M31 ;
    wire SubBytesIns_Inst_Sbox_9_M30 ;
    wire SubBytesIns_Inst_Sbox_9_M29 ;
    wire SubBytesIns_Inst_Sbox_9_M28 ;
    wire SubBytesIns_Inst_Sbox_9_M27 ;
    wire SubBytesIns_Inst_Sbox_9_M26 ;
    wire SubBytesIns_Inst_Sbox_9_M25 ;
    wire SubBytesIns_Inst_Sbox_9_M24 ;
    wire SubBytesIns_Inst_Sbox_9_M23 ;
    wire SubBytesIns_Inst_Sbox_9_M22 ;
    wire SubBytesIns_Inst_Sbox_9_M21 ;
    wire SubBytesIns_Inst_Sbox_9_M20 ;
    wire SubBytesIns_Inst_Sbox_9_M19 ;
    wire SubBytesIns_Inst_Sbox_9_M18 ;
    wire SubBytesIns_Inst_Sbox_9_M17 ;
    wire SubBytesIns_Inst_Sbox_9_M16 ;
    wire SubBytesIns_Inst_Sbox_9_M15 ;
    wire SubBytesIns_Inst_Sbox_9_M14 ;
    wire SubBytesIns_Inst_Sbox_9_M13 ;
    wire SubBytesIns_Inst_Sbox_9_M12 ;
    wire SubBytesIns_Inst_Sbox_9_M11 ;
    wire SubBytesIns_Inst_Sbox_9_M10 ;
    wire SubBytesIns_Inst_Sbox_9_M9 ;
    wire SubBytesIns_Inst_Sbox_9_M8 ;
    wire SubBytesIns_Inst_Sbox_9_M7 ;
    wire SubBytesIns_Inst_Sbox_9_M6 ;
    wire SubBytesIns_Inst_Sbox_9_M5 ;
    wire SubBytesIns_Inst_Sbox_9_M4 ;
    wire SubBytesIns_Inst_Sbox_9_M3 ;
    wire SubBytesIns_Inst_Sbox_9_M2 ;
    wire SubBytesIns_Inst_Sbox_9_M1 ;
    wire SubBytesIns_Inst_Sbox_9_T27 ;
    wire SubBytesIns_Inst_Sbox_9_T26 ;
    wire SubBytesIns_Inst_Sbox_9_T25 ;
    wire SubBytesIns_Inst_Sbox_9_T24 ;
    wire SubBytesIns_Inst_Sbox_9_T23 ;
    wire SubBytesIns_Inst_Sbox_9_T22 ;
    wire SubBytesIns_Inst_Sbox_9_T21 ;
    wire SubBytesIns_Inst_Sbox_9_T20 ;
    wire SubBytesIns_Inst_Sbox_9_T19 ;
    wire SubBytesIns_Inst_Sbox_9_T18 ;
    wire SubBytesIns_Inst_Sbox_9_T17 ;
    wire SubBytesIns_Inst_Sbox_9_T16 ;
    wire SubBytesIns_Inst_Sbox_9_T15 ;
    wire SubBytesIns_Inst_Sbox_9_T14 ;
    wire SubBytesIns_Inst_Sbox_9_T13 ;
    wire SubBytesIns_Inst_Sbox_9_T12 ;
    wire SubBytesIns_Inst_Sbox_9_T11 ;
    wire SubBytesIns_Inst_Sbox_9_T10 ;
    wire SubBytesIns_Inst_Sbox_9_T9 ;
    wire SubBytesIns_Inst_Sbox_9_T8 ;
    wire SubBytesIns_Inst_Sbox_9_T7 ;
    wire SubBytesIns_Inst_Sbox_9_T6 ;
    wire SubBytesIns_Inst_Sbox_9_T5 ;
    wire SubBytesIns_Inst_Sbox_9_T4 ;
    wire SubBytesIns_Inst_Sbox_9_T3 ;
    wire SubBytesIns_Inst_Sbox_9_T2 ;
    wire SubBytesIns_Inst_Sbox_9_T1 ;
    wire SubBytesIns_Inst_Sbox_10_L29 ;
    wire SubBytesIns_Inst_Sbox_10_L28 ;
    wire SubBytesIns_Inst_Sbox_10_L27 ;
    wire SubBytesIns_Inst_Sbox_10_L26 ;
    wire SubBytesIns_Inst_Sbox_10_L25 ;
    wire SubBytesIns_Inst_Sbox_10_L24 ;
    wire SubBytesIns_Inst_Sbox_10_L23 ;
    wire SubBytesIns_Inst_Sbox_10_L22 ;
    wire SubBytesIns_Inst_Sbox_10_L21 ;
    wire SubBytesIns_Inst_Sbox_10_L20 ;
    wire SubBytesIns_Inst_Sbox_10_L19 ;
    wire SubBytesIns_Inst_Sbox_10_L18 ;
    wire SubBytesIns_Inst_Sbox_10_L17 ;
    wire SubBytesIns_Inst_Sbox_10_L16 ;
    wire SubBytesIns_Inst_Sbox_10_L15 ;
    wire SubBytesIns_Inst_Sbox_10_L14 ;
    wire SubBytesIns_Inst_Sbox_10_L13 ;
    wire SubBytesIns_Inst_Sbox_10_L12 ;
    wire SubBytesIns_Inst_Sbox_10_L11 ;
    wire SubBytesIns_Inst_Sbox_10_L10 ;
    wire SubBytesIns_Inst_Sbox_10_L9 ;
    wire SubBytesIns_Inst_Sbox_10_L8 ;
    wire SubBytesIns_Inst_Sbox_10_L7 ;
    wire SubBytesIns_Inst_Sbox_10_L6 ;
    wire SubBytesIns_Inst_Sbox_10_L5 ;
    wire SubBytesIns_Inst_Sbox_10_L4 ;
    wire SubBytesIns_Inst_Sbox_10_L3 ;
    wire SubBytesIns_Inst_Sbox_10_L2 ;
    wire SubBytesIns_Inst_Sbox_10_L1 ;
    wire SubBytesIns_Inst_Sbox_10_L0 ;
    wire SubBytesIns_Inst_Sbox_10_M63 ;
    wire SubBytesIns_Inst_Sbox_10_M62 ;
    wire SubBytesIns_Inst_Sbox_10_M61 ;
    wire SubBytesIns_Inst_Sbox_10_M60 ;
    wire SubBytesIns_Inst_Sbox_10_M59 ;
    wire SubBytesIns_Inst_Sbox_10_M58 ;
    wire SubBytesIns_Inst_Sbox_10_M57 ;
    wire SubBytesIns_Inst_Sbox_10_M56 ;
    wire SubBytesIns_Inst_Sbox_10_M55 ;
    wire SubBytesIns_Inst_Sbox_10_M54 ;
    wire SubBytesIns_Inst_Sbox_10_M53 ;
    wire SubBytesIns_Inst_Sbox_10_M52 ;
    wire SubBytesIns_Inst_Sbox_10_M51 ;
    wire SubBytesIns_Inst_Sbox_10_M50 ;
    wire SubBytesIns_Inst_Sbox_10_M49 ;
    wire SubBytesIns_Inst_Sbox_10_M48 ;
    wire SubBytesIns_Inst_Sbox_10_M47 ;
    wire SubBytesIns_Inst_Sbox_10_M46 ;
    wire SubBytesIns_Inst_Sbox_10_M45 ;
    wire SubBytesIns_Inst_Sbox_10_M44 ;
    wire SubBytesIns_Inst_Sbox_10_M43 ;
    wire SubBytesIns_Inst_Sbox_10_M42 ;
    wire SubBytesIns_Inst_Sbox_10_M41 ;
    wire SubBytesIns_Inst_Sbox_10_M40 ;
    wire SubBytesIns_Inst_Sbox_10_M39 ;
    wire SubBytesIns_Inst_Sbox_10_M38 ;
    wire SubBytesIns_Inst_Sbox_10_M37 ;
    wire SubBytesIns_Inst_Sbox_10_M36 ;
    wire SubBytesIns_Inst_Sbox_10_M35 ;
    wire SubBytesIns_Inst_Sbox_10_M34 ;
    wire SubBytesIns_Inst_Sbox_10_M33 ;
    wire SubBytesIns_Inst_Sbox_10_M32 ;
    wire SubBytesIns_Inst_Sbox_10_M31 ;
    wire SubBytesIns_Inst_Sbox_10_M30 ;
    wire SubBytesIns_Inst_Sbox_10_M29 ;
    wire SubBytesIns_Inst_Sbox_10_M28 ;
    wire SubBytesIns_Inst_Sbox_10_M27 ;
    wire SubBytesIns_Inst_Sbox_10_M26 ;
    wire SubBytesIns_Inst_Sbox_10_M25 ;
    wire SubBytesIns_Inst_Sbox_10_M24 ;
    wire SubBytesIns_Inst_Sbox_10_M23 ;
    wire SubBytesIns_Inst_Sbox_10_M22 ;
    wire SubBytesIns_Inst_Sbox_10_M21 ;
    wire SubBytesIns_Inst_Sbox_10_M20 ;
    wire SubBytesIns_Inst_Sbox_10_M19 ;
    wire SubBytesIns_Inst_Sbox_10_M18 ;
    wire SubBytesIns_Inst_Sbox_10_M17 ;
    wire SubBytesIns_Inst_Sbox_10_M16 ;
    wire SubBytesIns_Inst_Sbox_10_M15 ;
    wire SubBytesIns_Inst_Sbox_10_M14 ;
    wire SubBytesIns_Inst_Sbox_10_M13 ;
    wire SubBytesIns_Inst_Sbox_10_M12 ;
    wire SubBytesIns_Inst_Sbox_10_M11 ;
    wire SubBytesIns_Inst_Sbox_10_M10 ;
    wire SubBytesIns_Inst_Sbox_10_M9 ;
    wire SubBytesIns_Inst_Sbox_10_M8 ;
    wire SubBytesIns_Inst_Sbox_10_M7 ;
    wire SubBytesIns_Inst_Sbox_10_M6 ;
    wire SubBytesIns_Inst_Sbox_10_M5 ;
    wire SubBytesIns_Inst_Sbox_10_M4 ;
    wire SubBytesIns_Inst_Sbox_10_M3 ;
    wire SubBytesIns_Inst_Sbox_10_M2 ;
    wire SubBytesIns_Inst_Sbox_10_M1 ;
    wire SubBytesIns_Inst_Sbox_10_T27 ;
    wire SubBytesIns_Inst_Sbox_10_T26 ;
    wire SubBytesIns_Inst_Sbox_10_T25 ;
    wire SubBytesIns_Inst_Sbox_10_T24 ;
    wire SubBytesIns_Inst_Sbox_10_T23 ;
    wire SubBytesIns_Inst_Sbox_10_T22 ;
    wire SubBytesIns_Inst_Sbox_10_T21 ;
    wire SubBytesIns_Inst_Sbox_10_T20 ;
    wire SubBytesIns_Inst_Sbox_10_T19 ;
    wire SubBytesIns_Inst_Sbox_10_T18 ;
    wire SubBytesIns_Inst_Sbox_10_T17 ;
    wire SubBytesIns_Inst_Sbox_10_T16 ;
    wire SubBytesIns_Inst_Sbox_10_T15 ;
    wire SubBytesIns_Inst_Sbox_10_T14 ;
    wire SubBytesIns_Inst_Sbox_10_T13 ;
    wire SubBytesIns_Inst_Sbox_10_T12 ;
    wire SubBytesIns_Inst_Sbox_10_T11 ;
    wire SubBytesIns_Inst_Sbox_10_T10 ;
    wire SubBytesIns_Inst_Sbox_10_T9 ;
    wire SubBytesIns_Inst_Sbox_10_T8 ;
    wire SubBytesIns_Inst_Sbox_10_T7 ;
    wire SubBytesIns_Inst_Sbox_10_T6 ;
    wire SubBytesIns_Inst_Sbox_10_T5 ;
    wire SubBytesIns_Inst_Sbox_10_T4 ;
    wire SubBytesIns_Inst_Sbox_10_T3 ;
    wire SubBytesIns_Inst_Sbox_10_T2 ;
    wire SubBytesIns_Inst_Sbox_10_T1 ;
    wire SubBytesIns_Inst_Sbox_11_L29 ;
    wire SubBytesIns_Inst_Sbox_11_L28 ;
    wire SubBytesIns_Inst_Sbox_11_L27 ;
    wire SubBytesIns_Inst_Sbox_11_L26 ;
    wire SubBytesIns_Inst_Sbox_11_L25 ;
    wire SubBytesIns_Inst_Sbox_11_L24 ;
    wire SubBytesIns_Inst_Sbox_11_L23 ;
    wire SubBytesIns_Inst_Sbox_11_L22 ;
    wire SubBytesIns_Inst_Sbox_11_L21 ;
    wire SubBytesIns_Inst_Sbox_11_L20 ;
    wire SubBytesIns_Inst_Sbox_11_L19 ;
    wire SubBytesIns_Inst_Sbox_11_L18 ;
    wire SubBytesIns_Inst_Sbox_11_L17 ;
    wire SubBytesIns_Inst_Sbox_11_L16 ;
    wire SubBytesIns_Inst_Sbox_11_L15 ;
    wire SubBytesIns_Inst_Sbox_11_L14 ;
    wire SubBytesIns_Inst_Sbox_11_L13 ;
    wire SubBytesIns_Inst_Sbox_11_L12 ;
    wire SubBytesIns_Inst_Sbox_11_L11 ;
    wire SubBytesIns_Inst_Sbox_11_L10 ;
    wire SubBytesIns_Inst_Sbox_11_L9 ;
    wire SubBytesIns_Inst_Sbox_11_L8 ;
    wire SubBytesIns_Inst_Sbox_11_L7 ;
    wire SubBytesIns_Inst_Sbox_11_L6 ;
    wire SubBytesIns_Inst_Sbox_11_L5 ;
    wire SubBytesIns_Inst_Sbox_11_L4 ;
    wire SubBytesIns_Inst_Sbox_11_L3 ;
    wire SubBytesIns_Inst_Sbox_11_L2 ;
    wire SubBytesIns_Inst_Sbox_11_L1 ;
    wire SubBytesIns_Inst_Sbox_11_L0 ;
    wire SubBytesIns_Inst_Sbox_11_M63 ;
    wire SubBytesIns_Inst_Sbox_11_M62 ;
    wire SubBytesIns_Inst_Sbox_11_M61 ;
    wire SubBytesIns_Inst_Sbox_11_M60 ;
    wire SubBytesIns_Inst_Sbox_11_M59 ;
    wire SubBytesIns_Inst_Sbox_11_M58 ;
    wire SubBytesIns_Inst_Sbox_11_M57 ;
    wire SubBytesIns_Inst_Sbox_11_M56 ;
    wire SubBytesIns_Inst_Sbox_11_M55 ;
    wire SubBytesIns_Inst_Sbox_11_M54 ;
    wire SubBytesIns_Inst_Sbox_11_M53 ;
    wire SubBytesIns_Inst_Sbox_11_M52 ;
    wire SubBytesIns_Inst_Sbox_11_M51 ;
    wire SubBytesIns_Inst_Sbox_11_M50 ;
    wire SubBytesIns_Inst_Sbox_11_M49 ;
    wire SubBytesIns_Inst_Sbox_11_M48 ;
    wire SubBytesIns_Inst_Sbox_11_M47 ;
    wire SubBytesIns_Inst_Sbox_11_M46 ;
    wire SubBytesIns_Inst_Sbox_11_M45 ;
    wire SubBytesIns_Inst_Sbox_11_M44 ;
    wire SubBytesIns_Inst_Sbox_11_M43 ;
    wire SubBytesIns_Inst_Sbox_11_M42 ;
    wire SubBytesIns_Inst_Sbox_11_M41 ;
    wire SubBytesIns_Inst_Sbox_11_M40 ;
    wire SubBytesIns_Inst_Sbox_11_M39 ;
    wire SubBytesIns_Inst_Sbox_11_M38 ;
    wire SubBytesIns_Inst_Sbox_11_M37 ;
    wire SubBytesIns_Inst_Sbox_11_M36 ;
    wire SubBytesIns_Inst_Sbox_11_M35 ;
    wire SubBytesIns_Inst_Sbox_11_M34 ;
    wire SubBytesIns_Inst_Sbox_11_M33 ;
    wire SubBytesIns_Inst_Sbox_11_M32 ;
    wire SubBytesIns_Inst_Sbox_11_M31 ;
    wire SubBytesIns_Inst_Sbox_11_M30 ;
    wire SubBytesIns_Inst_Sbox_11_M29 ;
    wire SubBytesIns_Inst_Sbox_11_M28 ;
    wire SubBytesIns_Inst_Sbox_11_M27 ;
    wire SubBytesIns_Inst_Sbox_11_M26 ;
    wire SubBytesIns_Inst_Sbox_11_M25 ;
    wire SubBytesIns_Inst_Sbox_11_M24 ;
    wire SubBytesIns_Inst_Sbox_11_M23 ;
    wire SubBytesIns_Inst_Sbox_11_M22 ;
    wire SubBytesIns_Inst_Sbox_11_M21 ;
    wire SubBytesIns_Inst_Sbox_11_M20 ;
    wire SubBytesIns_Inst_Sbox_11_M19 ;
    wire SubBytesIns_Inst_Sbox_11_M18 ;
    wire SubBytesIns_Inst_Sbox_11_M17 ;
    wire SubBytesIns_Inst_Sbox_11_M16 ;
    wire SubBytesIns_Inst_Sbox_11_M15 ;
    wire SubBytesIns_Inst_Sbox_11_M14 ;
    wire SubBytesIns_Inst_Sbox_11_M13 ;
    wire SubBytesIns_Inst_Sbox_11_M12 ;
    wire SubBytesIns_Inst_Sbox_11_M11 ;
    wire SubBytesIns_Inst_Sbox_11_M10 ;
    wire SubBytesIns_Inst_Sbox_11_M9 ;
    wire SubBytesIns_Inst_Sbox_11_M8 ;
    wire SubBytesIns_Inst_Sbox_11_M7 ;
    wire SubBytesIns_Inst_Sbox_11_M6 ;
    wire SubBytesIns_Inst_Sbox_11_M5 ;
    wire SubBytesIns_Inst_Sbox_11_M4 ;
    wire SubBytesIns_Inst_Sbox_11_M3 ;
    wire SubBytesIns_Inst_Sbox_11_M2 ;
    wire SubBytesIns_Inst_Sbox_11_M1 ;
    wire SubBytesIns_Inst_Sbox_11_T27 ;
    wire SubBytesIns_Inst_Sbox_11_T26 ;
    wire SubBytesIns_Inst_Sbox_11_T25 ;
    wire SubBytesIns_Inst_Sbox_11_T24 ;
    wire SubBytesIns_Inst_Sbox_11_T23 ;
    wire SubBytesIns_Inst_Sbox_11_T22 ;
    wire SubBytesIns_Inst_Sbox_11_T21 ;
    wire SubBytesIns_Inst_Sbox_11_T20 ;
    wire SubBytesIns_Inst_Sbox_11_T19 ;
    wire SubBytesIns_Inst_Sbox_11_T18 ;
    wire SubBytesIns_Inst_Sbox_11_T17 ;
    wire SubBytesIns_Inst_Sbox_11_T16 ;
    wire SubBytesIns_Inst_Sbox_11_T15 ;
    wire SubBytesIns_Inst_Sbox_11_T14 ;
    wire SubBytesIns_Inst_Sbox_11_T13 ;
    wire SubBytesIns_Inst_Sbox_11_T12 ;
    wire SubBytesIns_Inst_Sbox_11_T11 ;
    wire SubBytesIns_Inst_Sbox_11_T10 ;
    wire SubBytesIns_Inst_Sbox_11_T9 ;
    wire SubBytesIns_Inst_Sbox_11_T8 ;
    wire SubBytesIns_Inst_Sbox_11_T7 ;
    wire SubBytesIns_Inst_Sbox_11_T6 ;
    wire SubBytesIns_Inst_Sbox_11_T5 ;
    wire SubBytesIns_Inst_Sbox_11_T4 ;
    wire SubBytesIns_Inst_Sbox_11_T3 ;
    wire SubBytesIns_Inst_Sbox_11_T2 ;
    wire SubBytesIns_Inst_Sbox_11_T1 ;
    wire SubBytesIns_Inst_Sbox_12_L29 ;
    wire SubBytesIns_Inst_Sbox_12_L28 ;
    wire SubBytesIns_Inst_Sbox_12_L27 ;
    wire SubBytesIns_Inst_Sbox_12_L26 ;
    wire SubBytesIns_Inst_Sbox_12_L25 ;
    wire SubBytesIns_Inst_Sbox_12_L24 ;
    wire SubBytesIns_Inst_Sbox_12_L23 ;
    wire SubBytesIns_Inst_Sbox_12_L22 ;
    wire SubBytesIns_Inst_Sbox_12_L21 ;
    wire SubBytesIns_Inst_Sbox_12_L20 ;
    wire SubBytesIns_Inst_Sbox_12_L19 ;
    wire SubBytesIns_Inst_Sbox_12_L18 ;
    wire SubBytesIns_Inst_Sbox_12_L17 ;
    wire SubBytesIns_Inst_Sbox_12_L16 ;
    wire SubBytesIns_Inst_Sbox_12_L15 ;
    wire SubBytesIns_Inst_Sbox_12_L14 ;
    wire SubBytesIns_Inst_Sbox_12_L13 ;
    wire SubBytesIns_Inst_Sbox_12_L12 ;
    wire SubBytesIns_Inst_Sbox_12_L11 ;
    wire SubBytesIns_Inst_Sbox_12_L10 ;
    wire SubBytesIns_Inst_Sbox_12_L9 ;
    wire SubBytesIns_Inst_Sbox_12_L8 ;
    wire SubBytesIns_Inst_Sbox_12_L7 ;
    wire SubBytesIns_Inst_Sbox_12_L6 ;
    wire SubBytesIns_Inst_Sbox_12_L5 ;
    wire SubBytesIns_Inst_Sbox_12_L4 ;
    wire SubBytesIns_Inst_Sbox_12_L3 ;
    wire SubBytesIns_Inst_Sbox_12_L2 ;
    wire SubBytesIns_Inst_Sbox_12_L1 ;
    wire SubBytesIns_Inst_Sbox_12_L0 ;
    wire SubBytesIns_Inst_Sbox_12_M63 ;
    wire SubBytesIns_Inst_Sbox_12_M62 ;
    wire SubBytesIns_Inst_Sbox_12_M61 ;
    wire SubBytesIns_Inst_Sbox_12_M60 ;
    wire SubBytesIns_Inst_Sbox_12_M59 ;
    wire SubBytesIns_Inst_Sbox_12_M58 ;
    wire SubBytesIns_Inst_Sbox_12_M57 ;
    wire SubBytesIns_Inst_Sbox_12_M56 ;
    wire SubBytesIns_Inst_Sbox_12_M55 ;
    wire SubBytesIns_Inst_Sbox_12_M54 ;
    wire SubBytesIns_Inst_Sbox_12_M53 ;
    wire SubBytesIns_Inst_Sbox_12_M52 ;
    wire SubBytesIns_Inst_Sbox_12_M51 ;
    wire SubBytesIns_Inst_Sbox_12_M50 ;
    wire SubBytesIns_Inst_Sbox_12_M49 ;
    wire SubBytesIns_Inst_Sbox_12_M48 ;
    wire SubBytesIns_Inst_Sbox_12_M47 ;
    wire SubBytesIns_Inst_Sbox_12_M46 ;
    wire SubBytesIns_Inst_Sbox_12_M45 ;
    wire SubBytesIns_Inst_Sbox_12_M44 ;
    wire SubBytesIns_Inst_Sbox_12_M43 ;
    wire SubBytesIns_Inst_Sbox_12_M42 ;
    wire SubBytesIns_Inst_Sbox_12_M41 ;
    wire SubBytesIns_Inst_Sbox_12_M40 ;
    wire SubBytesIns_Inst_Sbox_12_M39 ;
    wire SubBytesIns_Inst_Sbox_12_M38 ;
    wire SubBytesIns_Inst_Sbox_12_M37 ;
    wire SubBytesIns_Inst_Sbox_12_M36 ;
    wire SubBytesIns_Inst_Sbox_12_M35 ;
    wire SubBytesIns_Inst_Sbox_12_M34 ;
    wire SubBytesIns_Inst_Sbox_12_M33 ;
    wire SubBytesIns_Inst_Sbox_12_M32 ;
    wire SubBytesIns_Inst_Sbox_12_M31 ;
    wire SubBytesIns_Inst_Sbox_12_M30 ;
    wire SubBytesIns_Inst_Sbox_12_M29 ;
    wire SubBytesIns_Inst_Sbox_12_M28 ;
    wire SubBytesIns_Inst_Sbox_12_M27 ;
    wire SubBytesIns_Inst_Sbox_12_M26 ;
    wire SubBytesIns_Inst_Sbox_12_M25 ;
    wire SubBytesIns_Inst_Sbox_12_M24 ;
    wire SubBytesIns_Inst_Sbox_12_M23 ;
    wire SubBytesIns_Inst_Sbox_12_M22 ;
    wire SubBytesIns_Inst_Sbox_12_M21 ;
    wire SubBytesIns_Inst_Sbox_12_M20 ;
    wire SubBytesIns_Inst_Sbox_12_M19 ;
    wire SubBytesIns_Inst_Sbox_12_M18 ;
    wire SubBytesIns_Inst_Sbox_12_M17 ;
    wire SubBytesIns_Inst_Sbox_12_M16 ;
    wire SubBytesIns_Inst_Sbox_12_M15 ;
    wire SubBytesIns_Inst_Sbox_12_M14 ;
    wire SubBytesIns_Inst_Sbox_12_M13 ;
    wire SubBytesIns_Inst_Sbox_12_M12 ;
    wire SubBytesIns_Inst_Sbox_12_M11 ;
    wire SubBytesIns_Inst_Sbox_12_M10 ;
    wire SubBytesIns_Inst_Sbox_12_M9 ;
    wire SubBytesIns_Inst_Sbox_12_M8 ;
    wire SubBytesIns_Inst_Sbox_12_M7 ;
    wire SubBytesIns_Inst_Sbox_12_M6 ;
    wire SubBytesIns_Inst_Sbox_12_M5 ;
    wire SubBytesIns_Inst_Sbox_12_M4 ;
    wire SubBytesIns_Inst_Sbox_12_M3 ;
    wire SubBytesIns_Inst_Sbox_12_M2 ;
    wire SubBytesIns_Inst_Sbox_12_M1 ;
    wire SubBytesIns_Inst_Sbox_12_T27 ;
    wire SubBytesIns_Inst_Sbox_12_T26 ;
    wire SubBytesIns_Inst_Sbox_12_T25 ;
    wire SubBytesIns_Inst_Sbox_12_T24 ;
    wire SubBytesIns_Inst_Sbox_12_T23 ;
    wire SubBytesIns_Inst_Sbox_12_T22 ;
    wire SubBytesIns_Inst_Sbox_12_T21 ;
    wire SubBytesIns_Inst_Sbox_12_T20 ;
    wire SubBytesIns_Inst_Sbox_12_T19 ;
    wire SubBytesIns_Inst_Sbox_12_T18 ;
    wire SubBytesIns_Inst_Sbox_12_T17 ;
    wire SubBytesIns_Inst_Sbox_12_T16 ;
    wire SubBytesIns_Inst_Sbox_12_T15 ;
    wire SubBytesIns_Inst_Sbox_12_T14 ;
    wire SubBytesIns_Inst_Sbox_12_T13 ;
    wire SubBytesIns_Inst_Sbox_12_T12 ;
    wire SubBytesIns_Inst_Sbox_12_T11 ;
    wire SubBytesIns_Inst_Sbox_12_T10 ;
    wire SubBytesIns_Inst_Sbox_12_T9 ;
    wire SubBytesIns_Inst_Sbox_12_T8 ;
    wire SubBytesIns_Inst_Sbox_12_T7 ;
    wire SubBytesIns_Inst_Sbox_12_T6 ;
    wire SubBytesIns_Inst_Sbox_12_T5 ;
    wire SubBytesIns_Inst_Sbox_12_T4 ;
    wire SubBytesIns_Inst_Sbox_12_T3 ;
    wire SubBytesIns_Inst_Sbox_12_T2 ;
    wire SubBytesIns_Inst_Sbox_12_T1 ;
    wire SubBytesIns_Inst_Sbox_13_L29 ;
    wire SubBytesIns_Inst_Sbox_13_L28 ;
    wire SubBytesIns_Inst_Sbox_13_L27 ;
    wire SubBytesIns_Inst_Sbox_13_L26 ;
    wire SubBytesIns_Inst_Sbox_13_L25 ;
    wire SubBytesIns_Inst_Sbox_13_L24 ;
    wire SubBytesIns_Inst_Sbox_13_L23 ;
    wire SubBytesIns_Inst_Sbox_13_L22 ;
    wire SubBytesIns_Inst_Sbox_13_L21 ;
    wire SubBytesIns_Inst_Sbox_13_L20 ;
    wire SubBytesIns_Inst_Sbox_13_L19 ;
    wire SubBytesIns_Inst_Sbox_13_L18 ;
    wire SubBytesIns_Inst_Sbox_13_L17 ;
    wire SubBytesIns_Inst_Sbox_13_L16 ;
    wire SubBytesIns_Inst_Sbox_13_L15 ;
    wire SubBytesIns_Inst_Sbox_13_L14 ;
    wire SubBytesIns_Inst_Sbox_13_L13 ;
    wire SubBytesIns_Inst_Sbox_13_L12 ;
    wire SubBytesIns_Inst_Sbox_13_L11 ;
    wire SubBytesIns_Inst_Sbox_13_L10 ;
    wire SubBytesIns_Inst_Sbox_13_L9 ;
    wire SubBytesIns_Inst_Sbox_13_L8 ;
    wire SubBytesIns_Inst_Sbox_13_L7 ;
    wire SubBytesIns_Inst_Sbox_13_L6 ;
    wire SubBytesIns_Inst_Sbox_13_L5 ;
    wire SubBytesIns_Inst_Sbox_13_L4 ;
    wire SubBytesIns_Inst_Sbox_13_L3 ;
    wire SubBytesIns_Inst_Sbox_13_L2 ;
    wire SubBytesIns_Inst_Sbox_13_L1 ;
    wire SubBytesIns_Inst_Sbox_13_L0 ;
    wire SubBytesIns_Inst_Sbox_13_M63 ;
    wire SubBytesIns_Inst_Sbox_13_M62 ;
    wire SubBytesIns_Inst_Sbox_13_M61 ;
    wire SubBytesIns_Inst_Sbox_13_M60 ;
    wire SubBytesIns_Inst_Sbox_13_M59 ;
    wire SubBytesIns_Inst_Sbox_13_M58 ;
    wire SubBytesIns_Inst_Sbox_13_M57 ;
    wire SubBytesIns_Inst_Sbox_13_M56 ;
    wire SubBytesIns_Inst_Sbox_13_M55 ;
    wire SubBytesIns_Inst_Sbox_13_M54 ;
    wire SubBytesIns_Inst_Sbox_13_M53 ;
    wire SubBytesIns_Inst_Sbox_13_M52 ;
    wire SubBytesIns_Inst_Sbox_13_M51 ;
    wire SubBytesIns_Inst_Sbox_13_M50 ;
    wire SubBytesIns_Inst_Sbox_13_M49 ;
    wire SubBytesIns_Inst_Sbox_13_M48 ;
    wire SubBytesIns_Inst_Sbox_13_M47 ;
    wire SubBytesIns_Inst_Sbox_13_M46 ;
    wire SubBytesIns_Inst_Sbox_13_M45 ;
    wire SubBytesIns_Inst_Sbox_13_M44 ;
    wire SubBytesIns_Inst_Sbox_13_M43 ;
    wire SubBytesIns_Inst_Sbox_13_M42 ;
    wire SubBytesIns_Inst_Sbox_13_M41 ;
    wire SubBytesIns_Inst_Sbox_13_M40 ;
    wire SubBytesIns_Inst_Sbox_13_M39 ;
    wire SubBytesIns_Inst_Sbox_13_M38 ;
    wire SubBytesIns_Inst_Sbox_13_M37 ;
    wire SubBytesIns_Inst_Sbox_13_M36 ;
    wire SubBytesIns_Inst_Sbox_13_M35 ;
    wire SubBytesIns_Inst_Sbox_13_M34 ;
    wire SubBytesIns_Inst_Sbox_13_M33 ;
    wire SubBytesIns_Inst_Sbox_13_M32 ;
    wire SubBytesIns_Inst_Sbox_13_M31 ;
    wire SubBytesIns_Inst_Sbox_13_M30 ;
    wire SubBytesIns_Inst_Sbox_13_M29 ;
    wire SubBytesIns_Inst_Sbox_13_M28 ;
    wire SubBytesIns_Inst_Sbox_13_M27 ;
    wire SubBytesIns_Inst_Sbox_13_M26 ;
    wire SubBytesIns_Inst_Sbox_13_M25 ;
    wire SubBytesIns_Inst_Sbox_13_M24 ;
    wire SubBytesIns_Inst_Sbox_13_M23 ;
    wire SubBytesIns_Inst_Sbox_13_M22 ;
    wire SubBytesIns_Inst_Sbox_13_M21 ;
    wire SubBytesIns_Inst_Sbox_13_M20 ;
    wire SubBytesIns_Inst_Sbox_13_M19 ;
    wire SubBytesIns_Inst_Sbox_13_M18 ;
    wire SubBytesIns_Inst_Sbox_13_M17 ;
    wire SubBytesIns_Inst_Sbox_13_M16 ;
    wire SubBytesIns_Inst_Sbox_13_M15 ;
    wire SubBytesIns_Inst_Sbox_13_M14 ;
    wire SubBytesIns_Inst_Sbox_13_M13 ;
    wire SubBytesIns_Inst_Sbox_13_M12 ;
    wire SubBytesIns_Inst_Sbox_13_M11 ;
    wire SubBytesIns_Inst_Sbox_13_M10 ;
    wire SubBytesIns_Inst_Sbox_13_M9 ;
    wire SubBytesIns_Inst_Sbox_13_M8 ;
    wire SubBytesIns_Inst_Sbox_13_M7 ;
    wire SubBytesIns_Inst_Sbox_13_M6 ;
    wire SubBytesIns_Inst_Sbox_13_M5 ;
    wire SubBytesIns_Inst_Sbox_13_M4 ;
    wire SubBytesIns_Inst_Sbox_13_M3 ;
    wire SubBytesIns_Inst_Sbox_13_M2 ;
    wire SubBytesIns_Inst_Sbox_13_M1 ;
    wire SubBytesIns_Inst_Sbox_13_T27 ;
    wire SubBytesIns_Inst_Sbox_13_T26 ;
    wire SubBytesIns_Inst_Sbox_13_T25 ;
    wire SubBytesIns_Inst_Sbox_13_T24 ;
    wire SubBytesIns_Inst_Sbox_13_T23 ;
    wire SubBytesIns_Inst_Sbox_13_T22 ;
    wire SubBytesIns_Inst_Sbox_13_T21 ;
    wire SubBytesIns_Inst_Sbox_13_T20 ;
    wire SubBytesIns_Inst_Sbox_13_T19 ;
    wire SubBytesIns_Inst_Sbox_13_T18 ;
    wire SubBytesIns_Inst_Sbox_13_T17 ;
    wire SubBytesIns_Inst_Sbox_13_T16 ;
    wire SubBytesIns_Inst_Sbox_13_T15 ;
    wire SubBytesIns_Inst_Sbox_13_T14 ;
    wire SubBytesIns_Inst_Sbox_13_T13 ;
    wire SubBytesIns_Inst_Sbox_13_T12 ;
    wire SubBytesIns_Inst_Sbox_13_T11 ;
    wire SubBytesIns_Inst_Sbox_13_T10 ;
    wire SubBytesIns_Inst_Sbox_13_T9 ;
    wire SubBytesIns_Inst_Sbox_13_T8 ;
    wire SubBytesIns_Inst_Sbox_13_T7 ;
    wire SubBytesIns_Inst_Sbox_13_T6 ;
    wire SubBytesIns_Inst_Sbox_13_T5 ;
    wire SubBytesIns_Inst_Sbox_13_T4 ;
    wire SubBytesIns_Inst_Sbox_13_T3 ;
    wire SubBytesIns_Inst_Sbox_13_T2 ;
    wire SubBytesIns_Inst_Sbox_13_T1 ;
    wire SubBytesIns_Inst_Sbox_14_L29 ;
    wire SubBytesIns_Inst_Sbox_14_L28 ;
    wire SubBytesIns_Inst_Sbox_14_L27 ;
    wire SubBytesIns_Inst_Sbox_14_L26 ;
    wire SubBytesIns_Inst_Sbox_14_L25 ;
    wire SubBytesIns_Inst_Sbox_14_L24 ;
    wire SubBytesIns_Inst_Sbox_14_L23 ;
    wire SubBytesIns_Inst_Sbox_14_L22 ;
    wire SubBytesIns_Inst_Sbox_14_L21 ;
    wire SubBytesIns_Inst_Sbox_14_L20 ;
    wire SubBytesIns_Inst_Sbox_14_L19 ;
    wire SubBytesIns_Inst_Sbox_14_L18 ;
    wire SubBytesIns_Inst_Sbox_14_L17 ;
    wire SubBytesIns_Inst_Sbox_14_L16 ;
    wire SubBytesIns_Inst_Sbox_14_L15 ;
    wire SubBytesIns_Inst_Sbox_14_L14 ;
    wire SubBytesIns_Inst_Sbox_14_L13 ;
    wire SubBytesIns_Inst_Sbox_14_L12 ;
    wire SubBytesIns_Inst_Sbox_14_L11 ;
    wire SubBytesIns_Inst_Sbox_14_L10 ;
    wire SubBytesIns_Inst_Sbox_14_L9 ;
    wire SubBytesIns_Inst_Sbox_14_L8 ;
    wire SubBytesIns_Inst_Sbox_14_L7 ;
    wire SubBytesIns_Inst_Sbox_14_L6 ;
    wire SubBytesIns_Inst_Sbox_14_L5 ;
    wire SubBytesIns_Inst_Sbox_14_L4 ;
    wire SubBytesIns_Inst_Sbox_14_L3 ;
    wire SubBytesIns_Inst_Sbox_14_L2 ;
    wire SubBytesIns_Inst_Sbox_14_L1 ;
    wire SubBytesIns_Inst_Sbox_14_L0 ;
    wire SubBytesIns_Inst_Sbox_14_M63 ;
    wire SubBytesIns_Inst_Sbox_14_M62 ;
    wire SubBytesIns_Inst_Sbox_14_M61 ;
    wire SubBytesIns_Inst_Sbox_14_M60 ;
    wire SubBytesIns_Inst_Sbox_14_M59 ;
    wire SubBytesIns_Inst_Sbox_14_M58 ;
    wire SubBytesIns_Inst_Sbox_14_M57 ;
    wire SubBytesIns_Inst_Sbox_14_M56 ;
    wire SubBytesIns_Inst_Sbox_14_M55 ;
    wire SubBytesIns_Inst_Sbox_14_M54 ;
    wire SubBytesIns_Inst_Sbox_14_M53 ;
    wire SubBytesIns_Inst_Sbox_14_M52 ;
    wire SubBytesIns_Inst_Sbox_14_M51 ;
    wire SubBytesIns_Inst_Sbox_14_M50 ;
    wire SubBytesIns_Inst_Sbox_14_M49 ;
    wire SubBytesIns_Inst_Sbox_14_M48 ;
    wire SubBytesIns_Inst_Sbox_14_M47 ;
    wire SubBytesIns_Inst_Sbox_14_M46 ;
    wire SubBytesIns_Inst_Sbox_14_M45 ;
    wire SubBytesIns_Inst_Sbox_14_M44 ;
    wire SubBytesIns_Inst_Sbox_14_M43 ;
    wire SubBytesIns_Inst_Sbox_14_M42 ;
    wire SubBytesIns_Inst_Sbox_14_M41 ;
    wire SubBytesIns_Inst_Sbox_14_M40 ;
    wire SubBytesIns_Inst_Sbox_14_M39 ;
    wire SubBytesIns_Inst_Sbox_14_M38 ;
    wire SubBytesIns_Inst_Sbox_14_M37 ;
    wire SubBytesIns_Inst_Sbox_14_M36 ;
    wire SubBytesIns_Inst_Sbox_14_M35 ;
    wire SubBytesIns_Inst_Sbox_14_M34 ;
    wire SubBytesIns_Inst_Sbox_14_M33 ;
    wire SubBytesIns_Inst_Sbox_14_M32 ;
    wire SubBytesIns_Inst_Sbox_14_M31 ;
    wire SubBytesIns_Inst_Sbox_14_M30 ;
    wire SubBytesIns_Inst_Sbox_14_M29 ;
    wire SubBytesIns_Inst_Sbox_14_M28 ;
    wire SubBytesIns_Inst_Sbox_14_M27 ;
    wire SubBytesIns_Inst_Sbox_14_M26 ;
    wire SubBytesIns_Inst_Sbox_14_M25 ;
    wire SubBytesIns_Inst_Sbox_14_M24 ;
    wire SubBytesIns_Inst_Sbox_14_M23 ;
    wire SubBytesIns_Inst_Sbox_14_M22 ;
    wire SubBytesIns_Inst_Sbox_14_M21 ;
    wire SubBytesIns_Inst_Sbox_14_M20 ;
    wire SubBytesIns_Inst_Sbox_14_M19 ;
    wire SubBytesIns_Inst_Sbox_14_M18 ;
    wire SubBytesIns_Inst_Sbox_14_M17 ;
    wire SubBytesIns_Inst_Sbox_14_M16 ;
    wire SubBytesIns_Inst_Sbox_14_M15 ;
    wire SubBytesIns_Inst_Sbox_14_M14 ;
    wire SubBytesIns_Inst_Sbox_14_M13 ;
    wire SubBytesIns_Inst_Sbox_14_M12 ;
    wire SubBytesIns_Inst_Sbox_14_M11 ;
    wire SubBytesIns_Inst_Sbox_14_M10 ;
    wire SubBytesIns_Inst_Sbox_14_M9 ;
    wire SubBytesIns_Inst_Sbox_14_M8 ;
    wire SubBytesIns_Inst_Sbox_14_M7 ;
    wire SubBytesIns_Inst_Sbox_14_M6 ;
    wire SubBytesIns_Inst_Sbox_14_M5 ;
    wire SubBytesIns_Inst_Sbox_14_M4 ;
    wire SubBytesIns_Inst_Sbox_14_M3 ;
    wire SubBytesIns_Inst_Sbox_14_M2 ;
    wire SubBytesIns_Inst_Sbox_14_M1 ;
    wire SubBytesIns_Inst_Sbox_14_T27 ;
    wire SubBytesIns_Inst_Sbox_14_T26 ;
    wire SubBytesIns_Inst_Sbox_14_T25 ;
    wire SubBytesIns_Inst_Sbox_14_T24 ;
    wire SubBytesIns_Inst_Sbox_14_T23 ;
    wire SubBytesIns_Inst_Sbox_14_T22 ;
    wire SubBytesIns_Inst_Sbox_14_T21 ;
    wire SubBytesIns_Inst_Sbox_14_T20 ;
    wire SubBytesIns_Inst_Sbox_14_T19 ;
    wire SubBytesIns_Inst_Sbox_14_T18 ;
    wire SubBytesIns_Inst_Sbox_14_T17 ;
    wire SubBytesIns_Inst_Sbox_14_T16 ;
    wire SubBytesIns_Inst_Sbox_14_T15 ;
    wire SubBytesIns_Inst_Sbox_14_T14 ;
    wire SubBytesIns_Inst_Sbox_14_T13 ;
    wire SubBytesIns_Inst_Sbox_14_T12 ;
    wire SubBytesIns_Inst_Sbox_14_T11 ;
    wire SubBytesIns_Inst_Sbox_14_T10 ;
    wire SubBytesIns_Inst_Sbox_14_T9 ;
    wire SubBytesIns_Inst_Sbox_14_T8 ;
    wire SubBytesIns_Inst_Sbox_14_T7 ;
    wire SubBytesIns_Inst_Sbox_14_T6 ;
    wire SubBytesIns_Inst_Sbox_14_T5 ;
    wire SubBytesIns_Inst_Sbox_14_T4 ;
    wire SubBytesIns_Inst_Sbox_14_T3 ;
    wire SubBytesIns_Inst_Sbox_14_T2 ;
    wire SubBytesIns_Inst_Sbox_14_T1 ;
    wire SubBytesIns_Inst_Sbox_15_L29 ;
    wire SubBytesIns_Inst_Sbox_15_L28 ;
    wire SubBytesIns_Inst_Sbox_15_L27 ;
    wire SubBytesIns_Inst_Sbox_15_L26 ;
    wire SubBytesIns_Inst_Sbox_15_L25 ;
    wire SubBytesIns_Inst_Sbox_15_L24 ;
    wire SubBytesIns_Inst_Sbox_15_L23 ;
    wire SubBytesIns_Inst_Sbox_15_L22 ;
    wire SubBytesIns_Inst_Sbox_15_L21 ;
    wire SubBytesIns_Inst_Sbox_15_L20 ;
    wire SubBytesIns_Inst_Sbox_15_L19 ;
    wire SubBytesIns_Inst_Sbox_15_L18 ;
    wire SubBytesIns_Inst_Sbox_15_L17 ;
    wire SubBytesIns_Inst_Sbox_15_L16 ;
    wire SubBytesIns_Inst_Sbox_15_L15 ;
    wire SubBytesIns_Inst_Sbox_15_L14 ;
    wire SubBytesIns_Inst_Sbox_15_L13 ;
    wire SubBytesIns_Inst_Sbox_15_L12 ;
    wire SubBytesIns_Inst_Sbox_15_L11 ;
    wire SubBytesIns_Inst_Sbox_15_L10 ;
    wire SubBytesIns_Inst_Sbox_15_L9 ;
    wire SubBytesIns_Inst_Sbox_15_L8 ;
    wire SubBytesIns_Inst_Sbox_15_L7 ;
    wire SubBytesIns_Inst_Sbox_15_L6 ;
    wire SubBytesIns_Inst_Sbox_15_L5 ;
    wire SubBytesIns_Inst_Sbox_15_L4 ;
    wire SubBytesIns_Inst_Sbox_15_L3 ;
    wire SubBytesIns_Inst_Sbox_15_L2 ;
    wire SubBytesIns_Inst_Sbox_15_L1 ;
    wire SubBytesIns_Inst_Sbox_15_L0 ;
    wire SubBytesIns_Inst_Sbox_15_M63 ;
    wire SubBytesIns_Inst_Sbox_15_M62 ;
    wire SubBytesIns_Inst_Sbox_15_M61 ;
    wire SubBytesIns_Inst_Sbox_15_M60 ;
    wire SubBytesIns_Inst_Sbox_15_M59 ;
    wire SubBytesIns_Inst_Sbox_15_M58 ;
    wire SubBytesIns_Inst_Sbox_15_M57 ;
    wire SubBytesIns_Inst_Sbox_15_M56 ;
    wire SubBytesIns_Inst_Sbox_15_M55 ;
    wire SubBytesIns_Inst_Sbox_15_M54 ;
    wire SubBytesIns_Inst_Sbox_15_M53 ;
    wire SubBytesIns_Inst_Sbox_15_M52 ;
    wire SubBytesIns_Inst_Sbox_15_M51 ;
    wire SubBytesIns_Inst_Sbox_15_M50 ;
    wire SubBytesIns_Inst_Sbox_15_M49 ;
    wire SubBytesIns_Inst_Sbox_15_M48 ;
    wire SubBytesIns_Inst_Sbox_15_M47 ;
    wire SubBytesIns_Inst_Sbox_15_M46 ;
    wire SubBytesIns_Inst_Sbox_15_M45 ;
    wire SubBytesIns_Inst_Sbox_15_M44 ;
    wire SubBytesIns_Inst_Sbox_15_M43 ;
    wire SubBytesIns_Inst_Sbox_15_M42 ;
    wire SubBytesIns_Inst_Sbox_15_M41 ;
    wire SubBytesIns_Inst_Sbox_15_M40 ;
    wire SubBytesIns_Inst_Sbox_15_M39 ;
    wire SubBytesIns_Inst_Sbox_15_M38 ;
    wire SubBytesIns_Inst_Sbox_15_M37 ;
    wire SubBytesIns_Inst_Sbox_15_M36 ;
    wire SubBytesIns_Inst_Sbox_15_M35 ;
    wire SubBytesIns_Inst_Sbox_15_M34 ;
    wire SubBytesIns_Inst_Sbox_15_M33 ;
    wire SubBytesIns_Inst_Sbox_15_M32 ;
    wire SubBytesIns_Inst_Sbox_15_M31 ;
    wire SubBytesIns_Inst_Sbox_15_M30 ;
    wire SubBytesIns_Inst_Sbox_15_M29 ;
    wire SubBytesIns_Inst_Sbox_15_M28 ;
    wire SubBytesIns_Inst_Sbox_15_M27 ;
    wire SubBytesIns_Inst_Sbox_15_M26 ;
    wire SubBytesIns_Inst_Sbox_15_M25 ;
    wire SubBytesIns_Inst_Sbox_15_M24 ;
    wire SubBytesIns_Inst_Sbox_15_M23 ;
    wire SubBytesIns_Inst_Sbox_15_M22 ;
    wire SubBytesIns_Inst_Sbox_15_M21 ;
    wire SubBytesIns_Inst_Sbox_15_M20 ;
    wire SubBytesIns_Inst_Sbox_15_M19 ;
    wire SubBytesIns_Inst_Sbox_15_M18 ;
    wire SubBytesIns_Inst_Sbox_15_M17 ;
    wire SubBytesIns_Inst_Sbox_15_M16 ;
    wire SubBytesIns_Inst_Sbox_15_M15 ;
    wire SubBytesIns_Inst_Sbox_15_M14 ;
    wire SubBytesIns_Inst_Sbox_15_M13 ;
    wire SubBytesIns_Inst_Sbox_15_M12 ;
    wire SubBytesIns_Inst_Sbox_15_M11 ;
    wire SubBytesIns_Inst_Sbox_15_M10 ;
    wire SubBytesIns_Inst_Sbox_15_M9 ;
    wire SubBytesIns_Inst_Sbox_15_M8 ;
    wire SubBytesIns_Inst_Sbox_15_M7 ;
    wire SubBytesIns_Inst_Sbox_15_M6 ;
    wire SubBytesIns_Inst_Sbox_15_M5 ;
    wire SubBytesIns_Inst_Sbox_15_M4 ;
    wire SubBytesIns_Inst_Sbox_15_M3 ;
    wire SubBytesIns_Inst_Sbox_15_M2 ;
    wire SubBytesIns_Inst_Sbox_15_M1 ;
    wire SubBytesIns_Inst_Sbox_15_T27 ;
    wire SubBytesIns_Inst_Sbox_15_T26 ;
    wire SubBytesIns_Inst_Sbox_15_T25 ;
    wire SubBytesIns_Inst_Sbox_15_T24 ;
    wire SubBytesIns_Inst_Sbox_15_T23 ;
    wire SubBytesIns_Inst_Sbox_15_T22 ;
    wire SubBytesIns_Inst_Sbox_15_T21 ;
    wire SubBytesIns_Inst_Sbox_15_T20 ;
    wire SubBytesIns_Inst_Sbox_15_T19 ;
    wire SubBytesIns_Inst_Sbox_15_T18 ;
    wire SubBytesIns_Inst_Sbox_15_T17 ;
    wire SubBytesIns_Inst_Sbox_15_T16 ;
    wire SubBytesIns_Inst_Sbox_15_T15 ;
    wire SubBytesIns_Inst_Sbox_15_T14 ;
    wire SubBytesIns_Inst_Sbox_15_T13 ;
    wire SubBytesIns_Inst_Sbox_15_T12 ;
    wire SubBytesIns_Inst_Sbox_15_T11 ;
    wire SubBytesIns_Inst_Sbox_15_T10 ;
    wire SubBytesIns_Inst_Sbox_15_T9 ;
    wire SubBytesIns_Inst_Sbox_15_T8 ;
    wire SubBytesIns_Inst_Sbox_15_T7 ;
    wire SubBytesIns_Inst_Sbox_15_T6 ;
    wire SubBytesIns_Inst_Sbox_15_T5 ;
    wire SubBytesIns_Inst_Sbox_15_T4 ;
    wire SubBytesIns_Inst_Sbox_15_T3 ;
    wire SubBytesIns_Inst_Sbox_15_T2 ;
    wire SubBytesIns_Inst_Sbox_15_T1 ;
    wire MixColumnsIns_MixOneColumnInst_0_n192 ;
    wire MixColumnsIns_MixOneColumnInst_0_n191 ;
    wire MixColumnsIns_MixOneColumnInst_0_n190 ;
    wire MixColumnsIns_MixOneColumnInst_0_n189 ;
    wire MixColumnsIns_MixOneColumnInst_0_n188 ;
    wire MixColumnsIns_MixOneColumnInst_0_n187 ;
    wire MixColumnsIns_MixOneColumnInst_0_n186 ;
    wire MixColumnsIns_MixOneColumnInst_0_n185 ;
    wire MixColumnsIns_MixOneColumnInst_0_n184 ;
    wire MixColumnsIns_MixOneColumnInst_0_n183 ;
    wire MixColumnsIns_MixOneColumnInst_0_n182 ;
    wire MixColumnsIns_MixOneColumnInst_0_n181 ;
    wire MixColumnsIns_MixOneColumnInst_0_n180 ;
    wire MixColumnsIns_MixOneColumnInst_0_n179 ;
    wire MixColumnsIns_MixOneColumnInst_0_n178 ;
    wire MixColumnsIns_MixOneColumnInst_0_n177 ;
    wire MixColumnsIns_MixOneColumnInst_0_n176 ;
    wire MixColumnsIns_MixOneColumnInst_0_n175 ;
    wire MixColumnsIns_MixOneColumnInst_0_n174 ;
    wire MixColumnsIns_MixOneColumnInst_0_n173 ;
    wire MixColumnsIns_MixOneColumnInst_0_n172 ;
    wire MixColumnsIns_MixOneColumnInst_0_n171 ;
    wire MixColumnsIns_MixOneColumnInst_0_n170 ;
    wire MixColumnsIns_MixOneColumnInst_0_n169 ;
    wire MixColumnsIns_MixOneColumnInst_0_n168 ;
    wire MixColumnsIns_MixOneColumnInst_0_n167 ;
    wire MixColumnsIns_MixOneColumnInst_0_n166 ;
    wire MixColumnsIns_MixOneColumnInst_0_n165 ;
    wire MixColumnsIns_MixOneColumnInst_0_n164 ;
    wire MixColumnsIns_MixOneColumnInst_0_n163 ;
    wire MixColumnsIns_MixOneColumnInst_0_n162 ;
    wire MixColumnsIns_MixOneColumnInst_0_n161 ;
    wire MixColumnsIns_MixOneColumnInst_0_n160 ;
    wire MixColumnsIns_MixOneColumnInst_0_n159 ;
    wire MixColumnsIns_MixOneColumnInst_0_n158 ;
    wire MixColumnsIns_MixOneColumnInst_0_n157 ;
    wire MixColumnsIns_MixOneColumnInst_0_n156 ;
    wire MixColumnsIns_MixOneColumnInst_0_n155 ;
    wire MixColumnsIns_MixOneColumnInst_0_n154 ;
    wire MixColumnsIns_MixOneColumnInst_0_n153 ;
    wire MixColumnsIns_MixOneColumnInst_0_n152 ;
    wire MixColumnsIns_MixOneColumnInst_0_n151 ;
    wire MixColumnsIns_MixOneColumnInst_0_n150 ;
    wire MixColumnsIns_MixOneColumnInst_0_n149 ;
    wire MixColumnsIns_MixOneColumnInst_0_n148 ;
    wire MixColumnsIns_MixOneColumnInst_0_n147 ;
    wire MixColumnsIns_MixOneColumnInst_0_n146 ;
    wire MixColumnsIns_MixOneColumnInst_0_n145 ;
    wire MixColumnsIns_MixOneColumnInst_0_n144 ;
    wire MixColumnsIns_MixOneColumnInst_0_n143 ;
    wire MixColumnsIns_MixOneColumnInst_0_n142 ;
    wire MixColumnsIns_MixOneColumnInst_0_n141 ;
    wire MixColumnsIns_MixOneColumnInst_0_n140 ;
    wire MixColumnsIns_MixOneColumnInst_0_n139 ;
    wire MixColumnsIns_MixOneColumnInst_0_n138 ;
    wire MixColumnsIns_MixOneColumnInst_0_n137 ;
    wire MixColumnsIns_MixOneColumnInst_0_n136 ;
    wire MixColumnsIns_MixOneColumnInst_0_n135 ;
    wire MixColumnsIns_MixOneColumnInst_0_n134 ;
    wire MixColumnsIns_MixOneColumnInst_0_n133 ;
    wire MixColumnsIns_MixOneColumnInst_0_n132 ;
    wire MixColumnsIns_MixOneColumnInst_0_n131 ;
    wire MixColumnsIns_MixOneColumnInst_0_n130 ;
    wire MixColumnsIns_MixOneColumnInst_0_n129 ;
    wire MixColumnsIns_MixOneColumnInst_1_n192 ;
    wire MixColumnsIns_MixOneColumnInst_1_n191 ;
    wire MixColumnsIns_MixOneColumnInst_1_n190 ;
    wire MixColumnsIns_MixOneColumnInst_1_n189 ;
    wire MixColumnsIns_MixOneColumnInst_1_n188 ;
    wire MixColumnsIns_MixOneColumnInst_1_n187 ;
    wire MixColumnsIns_MixOneColumnInst_1_n186 ;
    wire MixColumnsIns_MixOneColumnInst_1_n185 ;
    wire MixColumnsIns_MixOneColumnInst_1_n184 ;
    wire MixColumnsIns_MixOneColumnInst_1_n183 ;
    wire MixColumnsIns_MixOneColumnInst_1_n182 ;
    wire MixColumnsIns_MixOneColumnInst_1_n181 ;
    wire MixColumnsIns_MixOneColumnInst_1_n180 ;
    wire MixColumnsIns_MixOneColumnInst_1_n179 ;
    wire MixColumnsIns_MixOneColumnInst_1_n178 ;
    wire MixColumnsIns_MixOneColumnInst_1_n177 ;
    wire MixColumnsIns_MixOneColumnInst_1_n176 ;
    wire MixColumnsIns_MixOneColumnInst_1_n175 ;
    wire MixColumnsIns_MixOneColumnInst_1_n174 ;
    wire MixColumnsIns_MixOneColumnInst_1_n173 ;
    wire MixColumnsIns_MixOneColumnInst_1_n172 ;
    wire MixColumnsIns_MixOneColumnInst_1_n171 ;
    wire MixColumnsIns_MixOneColumnInst_1_n170 ;
    wire MixColumnsIns_MixOneColumnInst_1_n169 ;
    wire MixColumnsIns_MixOneColumnInst_1_n168 ;
    wire MixColumnsIns_MixOneColumnInst_1_n167 ;
    wire MixColumnsIns_MixOneColumnInst_1_n166 ;
    wire MixColumnsIns_MixOneColumnInst_1_n165 ;
    wire MixColumnsIns_MixOneColumnInst_1_n164 ;
    wire MixColumnsIns_MixOneColumnInst_1_n163 ;
    wire MixColumnsIns_MixOneColumnInst_1_n162 ;
    wire MixColumnsIns_MixOneColumnInst_1_n161 ;
    wire MixColumnsIns_MixOneColumnInst_1_n160 ;
    wire MixColumnsIns_MixOneColumnInst_1_n159 ;
    wire MixColumnsIns_MixOneColumnInst_1_n158 ;
    wire MixColumnsIns_MixOneColumnInst_1_n157 ;
    wire MixColumnsIns_MixOneColumnInst_1_n156 ;
    wire MixColumnsIns_MixOneColumnInst_1_n155 ;
    wire MixColumnsIns_MixOneColumnInst_1_n154 ;
    wire MixColumnsIns_MixOneColumnInst_1_n153 ;
    wire MixColumnsIns_MixOneColumnInst_1_n152 ;
    wire MixColumnsIns_MixOneColumnInst_1_n151 ;
    wire MixColumnsIns_MixOneColumnInst_1_n150 ;
    wire MixColumnsIns_MixOneColumnInst_1_n149 ;
    wire MixColumnsIns_MixOneColumnInst_1_n148 ;
    wire MixColumnsIns_MixOneColumnInst_1_n147 ;
    wire MixColumnsIns_MixOneColumnInst_1_n146 ;
    wire MixColumnsIns_MixOneColumnInst_1_n145 ;
    wire MixColumnsIns_MixOneColumnInst_1_n144 ;
    wire MixColumnsIns_MixOneColumnInst_1_n143 ;
    wire MixColumnsIns_MixOneColumnInst_1_n142 ;
    wire MixColumnsIns_MixOneColumnInst_1_n141 ;
    wire MixColumnsIns_MixOneColumnInst_1_n140 ;
    wire MixColumnsIns_MixOneColumnInst_1_n139 ;
    wire MixColumnsIns_MixOneColumnInst_1_n138 ;
    wire MixColumnsIns_MixOneColumnInst_1_n137 ;
    wire MixColumnsIns_MixOneColumnInst_1_n136 ;
    wire MixColumnsIns_MixOneColumnInst_1_n135 ;
    wire MixColumnsIns_MixOneColumnInst_1_n134 ;
    wire MixColumnsIns_MixOneColumnInst_1_n133 ;
    wire MixColumnsIns_MixOneColumnInst_1_n132 ;
    wire MixColumnsIns_MixOneColumnInst_1_n131 ;
    wire MixColumnsIns_MixOneColumnInst_1_n130 ;
    wire MixColumnsIns_MixOneColumnInst_1_n129 ;
    wire MixColumnsIns_MixOneColumnInst_2_n192 ;
    wire MixColumnsIns_MixOneColumnInst_2_n191 ;
    wire MixColumnsIns_MixOneColumnInst_2_n190 ;
    wire MixColumnsIns_MixOneColumnInst_2_n189 ;
    wire MixColumnsIns_MixOneColumnInst_2_n188 ;
    wire MixColumnsIns_MixOneColumnInst_2_n187 ;
    wire MixColumnsIns_MixOneColumnInst_2_n186 ;
    wire MixColumnsIns_MixOneColumnInst_2_n185 ;
    wire MixColumnsIns_MixOneColumnInst_2_n184 ;
    wire MixColumnsIns_MixOneColumnInst_2_n183 ;
    wire MixColumnsIns_MixOneColumnInst_2_n182 ;
    wire MixColumnsIns_MixOneColumnInst_2_n181 ;
    wire MixColumnsIns_MixOneColumnInst_2_n180 ;
    wire MixColumnsIns_MixOneColumnInst_2_n179 ;
    wire MixColumnsIns_MixOneColumnInst_2_n178 ;
    wire MixColumnsIns_MixOneColumnInst_2_n177 ;
    wire MixColumnsIns_MixOneColumnInst_2_n176 ;
    wire MixColumnsIns_MixOneColumnInst_2_n175 ;
    wire MixColumnsIns_MixOneColumnInst_2_n174 ;
    wire MixColumnsIns_MixOneColumnInst_2_n173 ;
    wire MixColumnsIns_MixOneColumnInst_2_n172 ;
    wire MixColumnsIns_MixOneColumnInst_2_n171 ;
    wire MixColumnsIns_MixOneColumnInst_2_n170 ;
    wire MixColumnsIns_MixOneColumnInst_2_n169 ;
    wire MixColumnsIns_MixOneColumnInst_2_n168 ;
    wire MixColumnsIns_MixOneColumnInst_2_n167 ;
    wire MixColumnsIns_MixOneColumnInst_2_n166 ;
    wire MixColumnsIns_MixOneColumnInst_2_n165 ;
    wire MixColumnsIns_MixOneColumnInst_2_n164 ;
    wire MixColumnsIns_MixOneColumnInst_2_n163 ;
    wire MixColumnsIns_MixOneColumnInst_2_n162 ;
    wire MixColumnsIns_MixOneColumnInst_2_n161 ;
    wire MixColumnsIns_MixOneColumnInst_2_n160 ;
    wire MixColumnsIns_MixOneColumnInst_2_n159 ;
    wire MixColumnsIns_MixOneColumnInst_2_n158 ;
    wire MixColumnsIns_MixOneColumnInst_2_n157 ;
    wire MixColumnsIns_MixOneColumnInst_2_n156 ;
    wire MixColumnsIns_MixOneColumnInst_2_n155 ;
    wire MixColumnsIns_MixOneColumnInst_2_n154 ;
    wire MixColumnsIns_MixOneColumnInst_2_n153 ;
    wire MixColumnsIns_MixOneColumnInst_2_n152 ;
    wire MixColumnsIns_MixOneColumnInst_2_n151 ;
    wire MixColumnsIns_MixOneColumnInst_2_n150 ;
    wire MixColumnsIns_MixOneColumnInst_2_n149 ;
    wire MixColumnsIns_MixOneColumnInst_2_n148 ;
    wire MixColumnsIns_MixOneColumnInst_2_n147 ;
    wire MixColumnsIns_MixOneColumnInst_2_n146 ;
    wire MixColumnsIns_MixOneColumnInst_2_n145 ;
    wire MixColumnsIns_MixOneColumnInst_2_n144 ;
    wire MixColumnsIns_MixOneColumnInst_2_n143 ;
    wire MixColumnsIns_MixOneColumnInst_2_n142 ;
    wire MixColumnsIns_MixOneColumnInst_2_n141 ;
    wire MixColumnsIns_MixOneColumnInst_2_n140 ;
    wire MixColumnsIns_MixOneColumnInst_2_n139 ;
    wire MixColumnsIns_MixOneColumnInst_2_n138 ;
    wire MixColumnsIns_MixOneColumnInst_2_n137 ;
    wire MixColumnsIns_MixOneColumnInst_2_n136 ;
    wire MixColumnsIns_MixOneColumnInst_2_n135 ;
    wire MixColumnsIns_MixOneColumnInst_2_n134 ;
    wire MixColumnsIns_MixOneColumnInst_2_n133 ;
    wire MixColumnsIns_MixOneColumnInst_2_n132 ;
    wire MixColumnsIns_MixOneColumnInst_2_n131 ;
    wire MixColumnsIns_MixOneColumnInst_2_n130 ;
    wire MixColumnsIns_MixOneColumnInst_2_n129 ;
    wire MixColumnsIns_MixOneColumnInst_3_n192 ;
    wire MixColumnsIns_MixOneColumnInst_3_n191 ;
    wire MixColumnsIns_MixOneColumnInst_3_n190 ;
    wire MixColumnsIns_MixOneColumnInst_3_n189 ;
    wire MixColumnsIns_MixOneColumnInst_3_n188 ;
    wire MixColumnsIns_MixOneColumnInst_3_n187 ;
    wire MixColumnsIns_MixOneColumnInst_3_n186 ;
    wire MixColumnsIns_MixOneColumnInst_3_n185 ;
    wire MixColumnsIns_MixOneColumnInst_3_n184 ;
    wire MixColumnsIns_MixOneColumnInst_3_n183 ;
    wire MixColumnsIns_MixOneColumnInst_3_n182 ;
    wire MixColumnsIns_MixOneColumnInst_3_n181 ;
    wire MixColumnsIns_MixOneColumnInst_3_n180 ;
    wire MixColumnsIns_MixOneColumnInst_3_n179 ;
    wire MixColumnsIns_MixOneColumnInst_3_n178 ;
    wire MixColumnsIns_MixOneColumnInst_3_n177 ;
    wire MixColumnsIns_MixOneColumnInst_3_n176 ;
    wire MixColumnsIns_MixOneColumnInst_3_n175 ;
    wire MixColumnsIns_MixOneColumnInst_3_n174 ;
    wire MixColumnsIns_MixOneColumnInst_3_n173 ;
    wire MixColumnsIns_MixOneColumnInst_3_n172 ;
    wire MixColumnsIns_MixOneColumnInst_3_n171 ;
    wire MixColumnsIns_MixOneColumnInst_3_n170 ;
    wire MixColumnsIns_MixOneColumnInst_3_n169 ;
    wire MixColumnsIns_MixOneColumnInst_3_n168 ;
    wire MixColumnsIns_MixOneColumnInst_3_n167 ;
    wire MixColumnsIns_MixOneColumnInst_3_n166 ;
    wire MixColumnsIns_MixOneColumnInst_3_n165 ;
    wire MixColumnsIns_MixOneColumnInst_3_n164 ;
    wire MixColumnsIns_MixOneColumnInst_3_n163 ;
    wire MixColumnsIns_MixOneColumnInst_3_n162 ;
    wire MixColumnsIns_MixOneColumnInst_3_n161 ;
    wire MixColumnsIns_MixOneColumnInst_3_n160 ;
    wire MixColumnsIns_MixOneColumnInst_3_n159 ;
    wire MixColumnsIns_MixOneColumnInst_3_n158 ;
    wire MixColumnsIns_MixOneColumnInst_3_n157 ;
    wire MixColumnsIns_MixOneColumnInst_3_n156 ;
    wire MixColumnsIns_MixOneColumnInst_3_n155 ;
    wire MixColumnsIns_MixOneColumnInst_3_n154 ;
    wire MixColumnsIns_MixOneColumnInst_3_n153 ;
    wire MixColumnsIns_MixOneColumnInst_3_n152 ;
    wire MixColumnsIns_MixOneColumnInst_3_n151 ;
    wire MixColumnsIns_MixOneColumnInst_3_n150 ;
    wire MixColumnsIns_MixOneColumnInst_3_n149 ;
    wire MixColumnsIns_MixOneColumnInst_3_n148 ;
    wire MixColumnsIns_MixOneColumnInst_3_n147 ;
    wire MixColumnsIns_MixOneColumnInst_3_n146 ;
    wire MixColumnsIns_MixOneColumnInst_3_n145 ;
    wire MixColumnsIns_MixOneColumnInst_3_n144 ;
    wire MixColumnsIns_MixOneColumnInst_3_n143 ;
    wire MixColumnsIns_MixOneColumnInst_3_n142 ;
    wire MixColumnsIns_MixOneColumnInst_3_n141 ;
    wire MixColumnsIns_MixOneColumnInst_3_n140 ;
    wire MixColumnsIns_MixOneColumnInst_3_n139 ;
    wire MixColumnsIns_MixOneColumnInst_3_n138 ;
    wire MixColumnsIns_MixOneColumnInst_3_n137 ;
    wire MixColumnsIns_MixOneColumnInst_3_n136 ;
    wire MixColumnsIns_MixOneColumnInst_3_n135 ;
    wire MixColumnsIns_MixOneColumnInst_3_n134 ;
    wire MixColumnsIns_MixOneColumnInst_3_n133 ;
    wire MixColumnsIns_MixOneColumnInst_3_n132 ;
    wire MixColumnsIns_MixOneColumnInst_3_n131 ;
    wire MixColumnsIns_MixOneColumnInst_3_n130 ;
    wire MixColumnsIns_MixOneColumnInst_3_n129 ;
    wire KeyReg_Inst_ff_SDE_0_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_0_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_1_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_1_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_2_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_2_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_3_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_3_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_4_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_4_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_5_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_5_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_6_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_6_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_7_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_7_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_8_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_8_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_9_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_9_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_10_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_10_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_11_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_11_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_12_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_12_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_13_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_13_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_14_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_14_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_15_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_15_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_16_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_16_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_17_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_17_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_18_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_18_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_19_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_19_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_20_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_20_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_21_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_21_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_22_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_22_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_23_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_23_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_24_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_24_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_25_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_25_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_26_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_26_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_27_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_27_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_28_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_28_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_29_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_29_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_30_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_30_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_31_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_31_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_32_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_32_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_33_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_33_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_34_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_34_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_35_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_35_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_36_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_36_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_37_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_37_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_38_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_38_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_39_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_39_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_40_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_40_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_41_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_41_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_42_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_42_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_43_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_43_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_44_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_44_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_45_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_45_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_46_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_46_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_47_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_47_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_48_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_48_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_49_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_49_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_50_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_50_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_51_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_51_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_52_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_52_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_53_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_53_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_54_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_54_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_55_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_55_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_56_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_56_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_57_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_57_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_58_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_58_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_59_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_59_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_60_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_60_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_61_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_61_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_62_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_62_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_63_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_63_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_64_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_64_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_65_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_65_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_66_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_66_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_67_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_67_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_68_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_68_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_69_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_69_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_70_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_70_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_71_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_71_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_72_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_72_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_73_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_73_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_74_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_74_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_75_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_75_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_76_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_76_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_77_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_77_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_78_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_78_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_79_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_79_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_80_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_80_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_81_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_81_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_82_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_82_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_83_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_83_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_84_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_84_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_85_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_85_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_86_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_86_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_87_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_87_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_88_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_88_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_89_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_89_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_90_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_90_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_91_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_91_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_92_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_92_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_93_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_93_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_94_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_94_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_95_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_95_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_96_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_96_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_97_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_97_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_98_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_98_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_99_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_99_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_100_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_100_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_101_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_101_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_102_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_102_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_103_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_103_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_104_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_104_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_105_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_105_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_106_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_106_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_107_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_107_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_108_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_108_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_109_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_109_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_110_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_110_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_111_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_111_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_112_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_112_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_113_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_113_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_114_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_114_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_115_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_115_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_116_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_116_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_117_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_117_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_118_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_118_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_119_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_119_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_120_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_120_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_121_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_121_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_122_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_122_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_123_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_123_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_124_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_124_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_125_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_125_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_126_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_126_MUX_inst_X ;
    wire KeyReg_Inst_ff_SDE_127_MUX_inst_Y ;
    wire KeyReg_Inst_ff_SDE_127_MUX_inst_X ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_ ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n3 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n1 ;
    wire [127:0] RoundOutput ;
    wire [127:0] RoundInput ;
    wire [127:0] RoundKey ;
    wire [123:0] MixColumnsInput ;
    wire [127:0] MixColumnsOutput ;
    wire [127:0] KeyExpansionOutput ;
    wire [5:0] Rcon ;
    wire [3:0] RoundCounter ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_0_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_1_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_2_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_3_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;

    /* cells in depth 0 */
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1093 ( .A0_t (RoundCounter[0]), .B0_t (n592), .Z0_t (n577) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1099 ( .A0_t (RoundCounter[3]), .B0_t (n585), .Z0_t (n592) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1100 ( .A0_t (RoundCounter[1]), .B0_t (RoundCounter[2]), .Z0_t (n585) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1103 ( .A0_t (RoundCounter[0]), .B0_t (n585), .Z0_t (Rcon[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1104 ( .A0_t (RoundCounter[0]), .B0_t (RoundCounter[3]), .Z0_t (n855) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1105 ( .A0_t (n855), .B0_t (n585), .Z0_t (Rcon[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1107 ( .A0_t (RoundCounter[2]), .B0_t (RoundCounter[1]), .Z0_t (n851) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1108 ( .A0_t (n855), .B0_t (n851), .Z0_t (n586) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1109 ( .A0_t (n577), .B0_t (n586), .Z0_t (Rcon[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1110 ( .A0_t (RoundCounter[3]), .B0_t (RoundCounter[0]), .Z0_t (n853) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1111 ( .A0_t (n851), .B0_t (n853), .Z0_t (n589) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1112 ( .A0_t (RoundCounter[3]), .B0_t (Rcon[0]), .Z0_t (n588) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1113 ( .A0_t (n589), .B0_t (n588), .Z0_t (Rcon[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1114 ( .A0_t (RoundCounter[1]), .B0_t (RoundCounter[2]), .Z0_t (n593) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1115 ( .A0_t (n855), .B0_t (n593), .Z0_t (n591) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1116 ( .A0_t (n592), .B0_t (n591), .Z0_t (Rcon[4]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1117 ( .A0_t (n853), .B0_t (n593), .Z0_t (n594) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1118 ( .A0_t (n577), .B0_t (n594), .Z0_t (Rcon[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1119 ( .A0_t (MixColumnsOutput[0]), .B0_t (n577), .Z0_t (n596) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1120 ( .A0_t (n577), .B0_t (MixColumnsInput[0]), .Z0_t (n595) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1121 ( .A0_t (n596), .B0_t (n595), .Z0_t (RoundOutput[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1122 ( .A0_t (MixColumnsOutput[100]), .B0_t (n577), .Z0_t (n598) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1123 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .Z0_t (n597) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1124 ( .A0_t (n598), .B0_t (n597), .Z0_t (RoundOutput[100]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1125 ( .A0_t (MixColumnsOutput[101]), .B0_t (n577), .Z0_t (n600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1126 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .Z0_t (n599) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1127 ( .A0_t (n600), .B0_t (n599), .Z0_t (RoundOutput[101]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1128 ( .A0_t (MixColumnsOutput[102]), .B0_t (n577), .Z0_t (n602) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1129 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .Z0_t (n601) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1130 ( .A0_t (n602), .B0_t (n601), .Z0_t (RoundOutput[102]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1131 ( .A0_t (MixColumnsOutput[103]), .B0_t (n577), .Z0_t (n604) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1132 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .Z0_t (n603) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1133 ( .A0_t (n604), .B0_t (n603), .Z0_t (RoundOutput[103]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1134 ( .A0_t (MixColumnsOutput[104]), .B0_t (n577), .Z0_t (n606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1135 ( .A0_t (n577), .B0_t (MixColumnsInput[104]), .Z0_t (n605) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1136 ( .A0_t (n606), .B0_t (n605), .Z0_t (RoundOutput[104]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1137 ( .A0_t (MixColumnsOutput[105]), .B0_t (n577), .Z0_t (n608) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1138 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .Z0_t (n607) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1139 ( .A0_t (n608), .B0_t (n607), .Z0_t (RoundOutput[105]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1140 ( .A0_t (MixColumnsOutput[106]), .B0_t (n577), .Z0_t (n610) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1141 ( .A0_t (n577), .B0_t (MixColumnsInput[106]), .Z0_t (n609) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1142 ( .A0_t (n610), .B0_t (n609), .Z0_t (RoundOutput[106]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1143 ( .A0_t (MixColumnsOutput[107]), .B0_t (n577), .Z0_t (n612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1144 ( .A0_t (n577), .B0_t (MixColumnsInput[107]), .Z0_t (n611) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1145 ( .A0_t (n612), .B0_t (n611), .Z0_t (RoundOutput[107]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1146 ( .A0_t (MixColumnsOutput[108]), .B0_t (n577), .Z0_t (n614) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1147 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .Z0_t (n613) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1148 ( .A0_t (n614), .B0_t (n613), .Z0_t (RoundOutput[108]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1149 ( .A0_t (MixColumnsOutput[109]), .B0_t (n577), .Z0_t (n616) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1150 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .Z0_t (n615) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1151 ( .A0_t (n616), .B0_t (n615), .Z0_t (RoundOutput[109]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1152 ( .A0_t (MixColumnsOutput[10]), .B0_t (n577), .Z0_t (n618) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1153 ( .A0_t (n577), .B0_t (MixColumnsInput[10]), .Z0_t (n617) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1154 ( .A0_t (n618), .B0_t (n617), .Z0_t (RoundOutput[10]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1155 ( .A0_t (MixColumnsOutput[110]), .B0_t (n577), .Z0_t (n620) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1156 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .Z0_t (n619) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1157 ( .A0_t (n620), .B0_t (n619), .Z0_t (RoundOutput[110]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1158 ( .A0_t (MixColumnsOutput[111]), .B0_t (n577), .Z0_t (n622) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1159 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .Z0_t (n621) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1160 ( .A0_t (n622), .B0_t (n621), .Z0_t (RoundOutput[111]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1161 ( .A0_t (MixColumnsOutput[112]), .B0_t (n577), .Z0_t (n624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1162 ( .A0_t (n577), .B0_t (MixColumnsInput[112]), .Z0_t (n623) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1163 ( .A0_t (n624), .B0_t (n623), .Z0_t (RoundOutput[112]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1164 ( .A0_t (MixColumnsOutput[113]), .B0_t (n577), .Z0_t (n626) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1165 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .Z0_t (n625) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1166 ( .A0_t (n626), .B0_t (n625), .Z0_t (RoundOutput[113]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1167 ( .A0_t (MixColumnsOutput[114]), .B0_t (n577), .Z0_t (n628) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1168 ( .A0_t (n577), .B0_t (MixColumnsInput[114]), .Z0_t (n627) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1169 ( .A0_t (n628), .B0_t (n627), .Z0_t (RoundOutput[114]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1170 ( .A0_t (MixColumnsOutput[115]), .B0_t (n577), .Z0_t (n630) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1171 ( .A0_t (n577), .B0_t (MixColumnsInput[115]), .Z0_t (n629) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1172 ( .A0_t (n630), .B0_t (n629), .Z0_t (RoundOutput[115]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1173 ( .A0_t (MixColumnsOutput[116]), .B0_t (n577), .Z0_t (n632) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1174 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .Z0_t (n631) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1175 ( .A0_t (n632), .B0_t (n631), .Z0_t (RoundOutput[116]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1176 ( .A0_t (MixColumnsOutput[117]), .B0_t (n577), .Z0_t (n634) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1177 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .Z0_t (n633) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1178 ( .A0_t (n634), .B0_t (n633), .Z0_t (RoundOutput[117]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1179 ( .A0_t (MixColumnsOutput[118]), .B0_t (n577), .Z0_t (n636) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1180 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .Z0_t (n635) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1181 ( .A0_t (n636), .B0_t (n635), .Z0_t (RoundOutput[118]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1182 ( .A0_t (MixColumnsOutput[119]), .B0_t (n577), .Z0_t (n638) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1183 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .Z0_t (n637) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1184 ( .A0_t (n638), .B0_t (n637), .Z0_t (RoundOutput[119]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1185 ( .A0_t (MixColumnsOutput[11]), .B0_t (n577), .Z0_t (n640) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1186 ( .A0_t (n577), .B0_t (MixColumnsInput[11]), .Z0_t (n639) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1187 ( .A0_t (n640), .B0_t (n639), .Z0_t (RoundOutput[11]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1188 ( .A0_t (MixColumnsOutput[120]), .B0_t (n577), .Z0_t (n642) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1189 ( .A0_t (n577), .B0_t (MixColumnsInput[120]), .Z0_t (n641) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1190 ( .A0_t (n642), .B0_t (n641), .Z0_t (RoundOutput[120]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1191 ( .A0_t (MixColumnsOutput[121]), .B0_t (n577), .Z0_t (n644) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1192 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .Z0_t (n643) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1193 ( .A0_t (n644), .B0_t (n643), .Z0_t (RoundOutput[121]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1194 ( .A0_t (MixColumnsOutput[122]), .B0_t (n577), .Z0_t (n646) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1195 ( .A0_t (n577), .B0_t (MixColumnsInput[122]), .Z0_t (n645) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1196 ( .A0_t (n646), .B0_t (n645), .Z0_t (RoundOutput[122]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1197 ( .A0_t (MixColumnsOutput[123]), .B0_t (n577), .Z0_t (n648) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1198 ( .A0_t (n577), .B0_t (MixColumnsInput[123]), .Z0_t (n647) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1199 ( .A0_t (n648), .B0_t (n647), .Z0_t (RoundOutput[123]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1200 ( .A0_t (MixColumnsOutput[124]), .B0_t (n577), .Z0_t (n650) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1201 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .Z0_t (n649) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1202 ( .A0_t (n650), .B0_t (n649), .Z0_t (RoundOutput[124]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1203 ( .A0_t (MixColumnsOutput[125]), .B0_t (n577), .Z0_t (n652) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1204 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .Z0_t (n651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1205 ( .A0_t (n652), .B0_t (n651), .Z0_t (RoundOutput[125]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1206 ( .A0_t (MixColumnsOutput[126]), .B0_t (n577), .Z0_t (n654) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1207 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .Z0_t (n653) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1208 ( .A0_t (n654), .B0_t (n653), .Z0_t (RoundOutput[126]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1209 ( .A0_t (MixColumnsOutput[127]), .B0_t (n577), .Z0_t (n656) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1210 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .Z0_t (n655) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1211 ( .A0_t (n656), .B0_t (n655), .Z0_t (RoundOutput[127]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1212 ( .A0_t (MixColumnsOutput[12]), .B0_t (n577), .Z0_t (n658) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1213 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .Z0_t (n657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1214 ( .A0_t (n658), .B0_t (n657), .Z0_t (RoundOutput[12]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1215 ( .A0_t (MixColumnsOutput[13]), .B0_t (n577), .Z0_t (n660) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1216 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .Z0_t (n659) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1217 ( .A0_t (n660), .B0_t (n659), .Z0_t (RoundOutput[13]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1218 ( .A0_t (MixColumnsOutput[14]), .B0_t (n577), .Z0_t (n662) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1219 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .Z0_t (n661) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1220 ( .A0_t (n662), .B0_t (n661), .Z0_t (RoundOutput[14]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1221 ( .A0_t (MixColumnsOutput[15]), .B0_t (n577), .Z0_t (n664) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1222 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .Z0_t (n663) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1223 ( .A0_t (n664), .B0_t (n663), .Z0_t (RoundOutput[15]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1224 ( .A0_t (MixColumnsOutput[16]), .B0_t (n577), .Z0_t (n666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1225 ( .A0_t (n577), .B0_t (MixColumnsInput[16]), .Z0_t (n665) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1226 ( .A0_t (n666), .B0_t (n665), .Z0_t (RoundOutput[16]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1227 ( .A0_t (MixColumnsOutput[17]), .B0_t (n577), .Z0_t (n668) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1228 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .Z0_t (n667) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1229 ( .A0_t (n668), .B0_t (n667), .Z0_t (RoundOutput[17]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1230 ( .A0_t (MixColumnsOutput[18]), .B0_t (n577), .Z0_t (n670) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1231 ( .A0_t (n577), .B0_t (MixColumnsInput[18]), .Z0_t (n669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1232 ( .A0_t (n670), .B0_t (n669), .Z0_t (RoundOutput[18]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1233 ( .A0_t (MixColumnsOutput[19]), .B0_t (n577), .Z0_t (n672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1234 ( .A0_t (n577), .B0_t (MixColumnsInput[19]), .Z0_t (n671) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1235 ( .A0_t (n672), .B0_t (n671), .Z0_t (RoundOutput[19]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1236 ( .A0_t (MixColumnsOutput[1]), .B0_t (n577), .Z0_t (n674) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1237 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .Z0_t (n673) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1238 ( .A0_t (n674), .B0_t (n673), .Z0_t (RoundOutput[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1239 ( .A0_t (MixColumnsOutput[20]), .B0_t (n577), .Z0_t (n676) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1240 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .Z0_t (n675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1241 ( .A0_t (n676), .B0_t (n675), .Z0_t (RoundOutput[20]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1242 ( .A0_t (MixColumnsOutput[21]), .B0_t (n577), .Z0_t (n678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1243 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .Z0_t (n677) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1244 ( .A0_t (n678), .B0_t (n677), .Z0_t (RoundOutput[21]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1245 ( .A0_t (MixColumnsOutput[22]), .B0_t (n577), .Z0_t (n680) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1246 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .Z0_t (n679) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1247 ( .A0_t (n680), .B0_t (n679), .Z0_t (RoundOutput[22]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1248 ( .A0_t (MixColumnsOutput[23]), .B0_t (n577), .Z0_t (n682) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1249 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .Z0_t (n681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1250 ( .A0_t (n682), .B0_t (n681), .Z0_t (RoundOutput[23]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1251 ( .A0_t (MixColumnsOutput[24]), .B0_t (n577), .Z0_t (n684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1252 ( .A0_t (n577), .B0_t (MixColumnsInput[24]), .Z0_t (n683) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1253 ( .A0_t (n684), .B0_t (n683), .Z0_t (RoundOutput[24]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1254 ( .A0_t (MixColumnsOutput[25]), .B0_t (n577), .Z0_t (n686) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1255 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .Z0_t (n685) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1256 ( .A0_t (n686), .B0_t (n685), .Z0_t (RoundOutput[25]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1257 ( .A0_t (MixColumnsOutput[26]), .B0_t (n577), .Z0_t (n688) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1258 ( .A0_t (n577), .B0_t (MixColumnsInput[26]), .Z0_t (n687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1259 ( .A0_t (n688), .B0_t (n687), .Z0_t (RoundOutput[26]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1260 ( .A0_t (MixColumnsOutput[27]), .B0_t (n577), .Z0_t (n690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1261 ( .A0_t (n577), .B0_t (MixColumnsInput[27]), .Z0_t (n689) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1262 ( .A0_t (n690), .B0_t (n689), .Z0_t (RoundOutput[27]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1263 ( .A0_t (MixColumnsOutput[28]), .B0_t (n577), .Z0_t (n692) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1264 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .Z0_t (n691) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1265 ( .A0_t (n692), .B0_t (n691), .Z0_t (RoundOutput[28]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1266 ( .A0_t (MixColumnsOutput[29]), .B0_t (n577), .Z0_t (n694) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1267 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .Z0_t (n693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1268 ( .A0_t (n694), .B0_t (n693), .Z0_t (RoundOutput[29]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1269 ( .A0_t (MixColumnsOutput[2]), .B0_t (n577), .Z0_t (n696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1270 ( .A0_t (n577), .B0_t (MixColumnsInput[2]), .Z0_t (n695) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1271 ( .A0_t (n696), .B0_t (n695), .Z0_t (RoundOutput[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1272 ( .A0_t (MixColumnsOutput[30]), .B0_t (n577), .Z0_t (n698) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1273 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .Z0_t (n697) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1274 ( .A0_t (n698), .B0_t (n697), .Z0_t (RoundOutput[30]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1275 ( .A0_t (MixColumnsOutput[31]), .B0_t (n577), .Z0_t (n700) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1276 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .Z0_t (n699) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1277 ( .A0_t (n700), .B0_t (n699), .Z0_t (RoundOutput[31]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1278 ( .A0_t (MixColumnsOutput[32]), .B0_t (n577), .Z0_t (n702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1279 ( .A0_t (n577), .B0_t (MixColumnsInput[32]), .Z0_t (n701) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1280 ( .A0_t (n702), .B0_t (n701), .Z0_t (RoundOutput[32]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1281 ( .A0_t (MixColumnsOutput[33]), .B0_t (n577), .Z0_t (n704) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1282 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .Z0_t (n703) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1283 ( .A0_t (n704), .B0_t (n703), .Z0_t (RoundOutput[33]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1284 ( .A0_t (MixColumnsOutput[34]), .B0_t (n577), .Z0_t (n706) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1285 ( .A0_t (n577), .B0_t (MixColumnsInput[34]), .Z0_t (n705) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1286 ( .A0_t (n706), .B0_t (n705), .Z0_t (RoundOutput[34]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1287 ( .A0_t (MixColumnsOutput[35]), .B0_t (n577), .Z0_t (n708) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1288 ( .A0_t (n577), .B0_t (MixColumnsInput[35]), .Z0_t (n707) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1289 ( .A0_t (n708), .B0_t (n707), .Z0_t (RoundOutput[35]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1290 ( .A0_t (MixColumnsOutput[36]), .B0_t (n577), .Z0_t (n710) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1291 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .Z0_t (n709) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1292 ( .A0_t (n710), .B0_t (n709), .Z0_t (RoundOutput[36]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1293 ( .A0_t (MixColumnsOutput[37]), .B0_t (n577), .Z0_t (n712) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1294 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .Z0_t (n711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1295 ( .A0_t (n712), .B0_t (n711), .Z0_t (RoundOutput[37]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1296 ( .A0_t (MixColumnsOutput[38]), .B0_t (n577), .Z0_t (n714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1297 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .Z0_t (n713) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1298 ( .A0_t (n714), .B0_t (n713), .Z0_t (RoundOutput[38]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1299 ( .A0_t (MixColumnsOutput[39]), .B0_t (n577), .Z0_t (n716) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1300 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .Z0_t (n715) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1301 ( .A0_t (n716), .B0_t (n715), .Z0_t (RoundOutput[39]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1302 ( .A0_t (MixColumnsOutput[3]), .B0_t (n577), .Z0_t (n718) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1303 ( .A0_t (n577), .B0_t (MixColumnsInput[3]), .Z0_t (n717) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1304 ( .A0_t (n718), .B0_t (n717), .Z0_t (RoundOutput[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1305 ( .A0_t (MixColumnsOutput[40]), .B0_t (n577), .Z0_t (n720) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1306 ( .A0_t (n577), .B0_t (MixColumnsInput[40]), .Z0_t (n719) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1307 ( .A0_t (n720), .B0_t (n719), .Z0_t (RoundOutput[40]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1308 ( .A0_t (MixColumnsOutput[41]), .B0_t (n577), .Z0_t (n722) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1309 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .Z0_t (n721) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1310 ( .A0_t (n722), .B0_t (n721), .Z0_t (RoundOutput[41]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1311 ( .A0_t (MixColumnsOutput[42]), .B0_t (n577), .Z0_t (n724) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1312 ( .A0_t (n577), .B0_t (MixColumnsInput[42]), .Z0_t (n723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1313 ( .A0_t (n724), .B0_t (n723), .Z0_t (RoundOutput[42]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1314 ( .A0_t (MixColumnsOutput[43]), .B0_t (n577), .Z0_t (n726) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1315 ( .A0_t (n577), .B0_t (MixColumnsInput[43]), .Z0_t (n725) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1316 ( .A0_t (n726), .B0_t (n725), .Z0_t (RoundOutput[43]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1317 ( .A0_t (MixColumnsOutput[44]), .B0_t (n577), .Z0_t (n728) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1318 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .Z0_t (n727) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1319 ( .A0_t (n728), .B0_t (n727), .Z0_t (RoundOutput[44]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1320 ( .A0_t (MixColumnsOutput[45]), .B0_t (n577), .Z0_t (n730) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1321 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .Z0_t (n729) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1322 ( .A0_t (n730), .B0_t (n729), .Z0_t (RoundOutput[45]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1323 ( .A0_t (MixColumnsOutput[46]), .B0_t (n577), .Z0_t (n732) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1324 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .Z0_t (n731) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1325 ( .A0_t (n732), .B0_t (n731), .Z0_t (RoundOutput[46]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1326 ( .A0_t (MixColumnsOutput[47]), .B0_t (n577), .Z0_t (n734) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1327 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .Z0_t (n733) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1328 ( .A0_t (n734), .B0_t (n733), .Z0_t (RoundOutput[47]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1329 ( .A0_t (MixColumnsOutput[48]), .B0_t (n577), .Z0_t (n736) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1330 ( .A0_t (n577), .B0_t (MixColumnsInput[48]), .Z0_t (n735) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1331 ( .A0_t (n736), .B0_t (n735), .Z0_t (RoundOutput[48]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1332 ( .A0_t (MixColumnsOutput[49]), .B0_t (n577), .Z0_t (n738) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1333 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .Z0_t (n737) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1334 ( .A0_t (n738), .B0_t (n737), .Z0_t (RoundOutput[49]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1335 ( .A0_t (MixColumnsOutput[4]), .B0_t (n577), .Z0_t (n740) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1336 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .Z0_t (n739) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1337 ( .A0_t (n740), .B0_t (n739), .Z0_t (RoundOutput[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1338 ( .A0_t (MixColumnsOutput[50]), .B0_t (n577), .Z0_t (n742) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1339 ( .A0_t (n577), .B0_t (MixColumnsInput[50]), .Z0_t (n741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1340 ( .A0_t (n742), .B0_t (n741), .Z0_t (RoundOutput[50]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1341 ( .A0_t (MixColumnsOutput[51]), .B0_t (n577), .Z0_t (n744) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1342 ( .A0_t (n577), .B0_t (MixColumnsInput[51]), .Z0_t (n743) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1343 ( .A0_t (n744), .B0_t (n743), .Z0_t (RoundOutput[51]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1344 ( .A0_t (MixColumnsOutput[52]), .B0_t (n577), .Z0_t (n746) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1345 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .Z0_t (n745) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1346 ( .A0_t (n746), .B0_t (n745), .Z0_t (RoundOutput[52]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1347 ( .A0_t (MixColumnsOutput[53]), .B0_t (n577), .Z0_t (n748) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1348 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .Z0_t (n747) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1349 ( .A0_t (n748), .B0_t (n747), .Z0_t (RoundOutput[53]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1350 ( .A0_t (MixColumnsOutput[54]), .B0_t (n577), .Z0_t (n750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1351 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .Z0_t (n749) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1352 ( .A0_t (n750), .B0_t (n749), .Z0_t (RoundOutput[54]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1353 ( .A0_t (MixColumnsOutput[55]), .B0_t (n577), .Z0_t (n752) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1354 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .Z0_t (n751) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1355 ( .A0_t (n752), .B0_t (n751), .Z0_t (RoundOutput[55]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1356 ( .A0_t (MixColumnsOutput[56]), .B0_t (n577), .Z0_t (n754) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1357 ( .A0_t (n577), .B0_t (MixColumnsInput[56]), .Z0_t (n753) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1358 ( .A0_t (n754), .B0_t (n753), .Z0_t (RoundOutput[56]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1359 ( .A0_t (MixColumnsOutput[57]), .B0_t (n577), .Z0_t (n756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1360 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .Z0_t (n755) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1361 ( .A0_t (n756), .B0_t (n755), .Z0_t (RoundOutput[57]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1362 ( .A0_t (MixColumnsOutput[58]), .B0_t (n577), .Z0_t (n758) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1363 ( .A0_t (n577), .B0_t (MixColumnsInput[58]), .Z0_t (n757) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1364 ( .A0_t (n758), .B0_t (n757), .Z0_t (RoundOutput[58]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1365 ( .A0_t (MixColumnsOutput[59]), .B0_t (n577), .Z0_t (n760) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1366 ( .A0_t (n577), .B0_t (MixColumnsInput[59]), .Z0_t (n759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1367 ( .A0_t (n760), .B0_t (n759), .Z0_t (RoundOutput[59]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1368 ( .A0_t (MixColumnsOutput[5]), .B0_t (n577), .Z0_t (n762) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1369 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .Z0_t (n761) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1370 ( .A0_t (n762), .B0_t (n761), .Z0_t (RoundOutput[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1371 ( .A0_t (MixColumnsOutput[60]), .B0_t (n577), .Z0_t (n764) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1372 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .Z0_t (n763) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1373 ( .A0_t (n764), .B0_t (n763), .Z0_t (RoundOutput[60]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1374 ( .A0_t (MixColumnsOutput[61]), .B0_t (n577), .Z0_t (n766) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1375 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .Z0_t (n765) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1376 ( .A0_t (n766), .B0_t (n765), .Z0_t (RoundOutput[61]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1377 ( .A0_t (MixColumnsOutput[62]), .B0_t (n577), .Z0_t (n768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1378 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .Z0_t (n767) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1379 ( .A0_t (n768), .B0_t (n767), .Z0_t (RoundOutput[62]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1380 ( .A0_t (MixColumnsOutput[63]), .B0_t (n577), .Z0_t (n770) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1381 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .Z0_t (n769) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1382 ( .A0_t (n770), .B0_t (n769), .Z0_t (RoundOutput[63]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1383 ( .A0_t (MixColumnsOutput[64]), .B0_t (n577), .Z0_t (n772) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1384 ( .A0_t (n577), .B0_t (MixColumnsInput[64]), .Z0_t (n771) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1385 ( .A0_t (n772), .B0_t (n771), .Z0_t (RoundOutput[64]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1386 ( .A0_t (MixColumnsOutput[65]), .B0_t (n577), .Z0_t (n774) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1387 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .Z0_t (n773) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1388 ( .A0_t (n774), .B0_t (n773), .Z0_t (RoundOutput[65]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1389 ( .A0_t (MixColumnsOutput[66]), .B0_t (n577), .Z0_t (n776) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1390 ( .A0_t (n577), .B0_t (MixColumnsInput[66]), .Z0_t (n775) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1391 ( .A0_t (n776), .B0_t (n775), .Z0_t (RoundOutput[66]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1392 ( .A0_t (MixColumnsOutput[67]), .B0_t (n577), .Z0_t (n778) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1393 ( .A0_t (n577), .B0_t (MixColumnsInput[67]), .Z0_t (n777) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1394 ( .A0_t (n778), .B0_t (n777), .Z0_t (RoundOutput[67]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1395 ( .A0_t (MixColumnsOutput[68]), .B0_t (n577), .Z0_t (n780) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1396 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .Z0_t (n779) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1397 ( .A0_t (n780), .B0_t (n779), .Z0_t (RoundOutput[68]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1398 ( .A0_t (MixColumnsOutput[69]), .B0_t (n577), .Z0_t (n782) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1399 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .Z0_t (n781) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1400 ( .A0_t (n782), .B0_t (n781), .Z0_t (RoundOutput[69]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1401 ( .A0_t (MixColumnsOutput[6]), .B0_t (n577), .Z0_t (n784) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1402 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .Z0_t (n783) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1403 ( .A0_t (n784), .B0_t (n783), .Z0_t (RoundOutput[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1404 ( .A0_t (MixColumnsOutput[70]), .B0_t (n577), .Z0_t (n786) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1405 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .Z0_t (n785) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1406 ( .A0_t (n786), .B0_t (n785), .Z0_t (RoundOutput[70]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1407 ( .A0_t (MixColumnsOutput[71]), .B0_t (n577), .Z0_t (n788) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1408 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .Z0_t (n787) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1409 ( .A0_t (n788), .B0_t (n787), .Z0_t (RoundOutput[71]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1410 ( .A0_t (MixColumnsOutput[72]), .B0_t (n577), .Z0_t (n790) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1411 ( .A0_t (n577), .B0_t (MixColumnsInput[72]), .Z0_t (n789) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1412 ( .A0_t (n790), .B0_t (n789), .Z0_t (RoundOutput[72]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1413 ( .A0_t (MixColumnsOutput[73]), .B0_t (n577), .Z0_t (n792) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1414 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .Z0_t (n791) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1415 ( .A0_t (n792), .B0_t (n791), .Z0_t (RoundOutput[73]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1416 ( .A0_t (MixColumnsOutput[74]), .B0_t (n577), .Z0_t (n794) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1417 ( .A0_t (n577), .B0_t (MixColumnsInput[74]), .Z0_t (n793) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1418 ( .A0_t (n794), .B0_t (n793), .Z0_t (RoundOutput[74]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1419 ( .A0_t (MixColumnsOutput[75]), .B0_t (n577), .Z0_t (n796) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1420 ( .A0_t (n577), .B0_t (MixColumnsInput[75]), .Z0_t (n795) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1421 ( .A0_t (n796), .B0_t (n795), .Z0_t (RoundOutput[75]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1422 ( .A0_t (MixColumnsOutput[76]), .B0_t (n577), .Z0_t (n798) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1423 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .Z0_t (n797) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1424 ( .A0_t (n798), .B0_t (n797), .Z0_t (RoundOutput[76]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1425 ( .A0_t (MixColumnsOutput[77]), .B0_t (n577), .Z0_t (n800) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1426 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .Z0_t (n799) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1427 ( .A0_t (n800), .B0_t (n799), .Z0_t (RoundOutput[77]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1428 ( .A0_t (MixColumnsOutput[78]), .B0_t (n577), .Z0_t (n802) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1429 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .Z0_t (n801) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1430 ( .A0_t (n802), .B0_t (n801), .Z0_t (RoundOutput[78]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1431 ( .A0_t (MixColumnsOutput[79]), .B0_t (n577), .Z0_t (n804) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1432 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .Z0_t (n803) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1433 ( .A0_t (n804), .B0_t (n803), .Z0_t (RoundOutput[79]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1434 ( .A0_t (MixColumnsOutput[7]), .B0_t (n577), .Z0_t (n806) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1435 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .Z0_t (n805) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1436 ( .A0_t (n806), .B0_t (n805), .Z0_t (RoundOutput[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1437 ( .A0_t (MixColumnsOutput[80]), .B0_t (n577), .Z0_t (n808) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1438 ( .A0_t (n577), .B0_t (MixColumnsInput[80]), .Z0_t (n807) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1439 ( .A0_t (n808), .B0_t (n807), .Z0_t (RoundOutput[80]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1440 ( .A0_t (MixColumnsOutput[81]), .B0_t (n577), .Z0_t (n810) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1441 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .Z0_t (n809) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1442 ( .A0_t (n810), .B0_t (n809), .Z0_t (RoundOutput[81]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1443 ( .A0_t (MixColumnsOutput[82]), .B0_t (n577), .Z0_t (n812) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1444 ( .A0_t (n577), .B0_t (MixColumnsInput[82]), .Z0_t (n811) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1445 ( .A0_t (n812), .B0_t (n811), .Z0_t (RoundOutput[82]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1446 ( .A0_t (MixColumnsOutput[83]), .B0_t (n577), .Z0_t (n814) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1447 ( .A0_t (n577), .B0_t (MixColumnsInput[83]), .Z0_t (n813) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1448 ( .A0_t (n814), .B0_t (n813), .Z0_t (RoundOutput[83]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1449 ( .A0_t (MixColumnsOutput[84]), .B0_t (n577), .Z0_t (n816) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1450 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .Z0_t (n815) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1451 ( .A0_t (n816), .B0_t (n815), .Z0_t (RoundOutput[84]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1452 ( .A0_t (MixColumnsOutput[85]), .B0_t (n577), .Z0_t (n818) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1453 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .Z0_t (n817) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1454 ( .A0_t (n818), .B0_t (n817), .Z0_t (RoundOutput[85]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1455 ( .A0_t (MixColumnsOutput[86]), .B0_t (n577), .Z0_t (n820) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1456 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .Z0_t (n819) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1457 ( .A0_t (n820), .B0_t (n819), .Z0_t (RoundOutput[86]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1458 ( .A0_t (MixColumnsOutput[87]), .B0_t (n577), .Z0_t (n822) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1459 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .Z0_t (n821) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1460 ( .A0_t (n822), .B0_t (n821), .Z0_t (RoundOutput[87]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1461 ( .A0_t (MixColumnsOutput[88]), .B0_t (n577), .Z0_t (n824) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1462 ( .A0_t (n577), .B0_t (MixColumnsInput[88]), .Z0_t (n823) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1463 ( .A0_t (n824), .B0_t (n823), .Z0_t (RoundOutput[88]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1464 ( .A0_t (MixColumnsOutput[89]), .B0_t (n577), .Z0_t (n826) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1465 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .Z0_t (n825) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1466 ( .A0_t (n826), .B0_t (n825), .Z0_t (RoundOutput[89]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1467 ( .A0_t (MixColumnsOutput[8]), .B0_t (n577), .Z0_t (n828) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1468 ( .A0_t (n577), .B0_t (MixColumnsInput[8]), .Z0_t (n827) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1469 ( .A0_t (n828), .B0_t (n827), .Z0_t (RoundOutput[8]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1470 ( .A0_t (MixColumnsOutput[90]), .B0_t (n577), .Z0_t (n830) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1471 ( .A0_t (n577), .B0_t (MixColumnsInput[90]), .Z0_t (n829) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1472 ( .A0_t (n830), .B0_t (n829), .Z0_t (RoundOutput[90]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1473 ( .A0_t (MixColumnsOutput[91]), .B0_t (n577), .Z0_t (n832) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1474 ( .A0_t (n577), .B0_t (MixColumnsInput[91]), .Z0_t (n831) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1475 ( .A0_t (n832), .B0_t (n831), .Z0_t (RoundOutput[91]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1476 ( .A0_t (MixColumnsOutput[92]), .B0_t (n577), .Z0_t (n834) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1477 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .Z0_t (n833) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1478 ( .A0_t (n834), .B0_t (n833), .Z0_t (RoundOutput[92]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1479 ( .A0_t (MixColumnsOutput[93]), .B0_t (n577), .Z0_t (n836) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1480 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .Z0_t (n835) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1481 ( .A0_t (n836), .B0_t (n835), .Z0_t (RoundOutput[93]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1482 ( .A0_t (MixColumnsOutput[94]), .B0_t (n577), .Z0_t (n838) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1483 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .Z0_t (n837) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1484 ( .A0_t (n838), .B0_t (n837), .Z0_t (RoundOutput[94]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1485 ( .A0_t (MixColumnsOutput[95]), .B0_t (n577), .Z0_t (n840) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1486 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .Z0_t (n839) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1487 ( .A0_t (n840), .B0_t (n839), .Z0_t (RoundOutput[95]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1488 ( .A0_t (MixColumnsOutput[96]), .B0_t (n577), .Z0_t (n842) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1489 ( .A0_t (n577), .B0_t (MixColumnsInput[96]), .Z0_t (n841) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1490 ( .A0_t (n842), .B0_t (n841), .Z0_t (RoundOutput[96]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1491 ( .A0_t (MixColumnsOutput[97]), .B0_t (n577), .Z0_t (n844) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1492 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .Z0_t (n843) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1493 ( .A0_t (n844), .B0_t (n843), .Z0_t (RoundOutput[97]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1494 ( .A0_t (MixColumnsOutput[98]), .B0_t (n577), .Z0_t (n846) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1495 ( .A0_t (n577), .B0_t (MixColumnsInput[98]), .Z0_t (n845) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1496 ( .A0_t (n846), .B0_t (n845), .Z0_t (RoundOutput[98]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1497 ( .A0_t (MixColumnsOutput[99]), .B0_t (n577), .Z0_t (n848) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1498 ( .A0_t (n577), .B0_t (MixColumnsInput[99]), .Z0_t (n847) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1499 ( .A0_t (n848), .B0_t (n847), .Z0_t (RoundOutput[99]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1500 ( .A0_t (MixColumnsOutput[9]), .B0_t (n577), .Z0_t (n850) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1501 ( .A0_t (n577), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .Z0_t (n849) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) U1502 ( .A0_t (n850), .B0_t (n849), .Z0_t (RoundOutput[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1503 ( .A0_t (RoundInput[0]), .B0_t (RoundKey[0]), .Z0_t (ciphertext[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1504 ( .A0_t (RoundInput[100]), .B0_t (RoundKey[100]), .Z0_t (ciphertext[100]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1505 ( .A0_t (RoundInput[101]), .B0_t (RoundKey[101]), .Z0_t (ciphertext[101]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1506 ( .A0_t (RoundInput[102]), .B0_t (RoundKey[102]), .Z0_t (ciphertext[102]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1507 ( .A0_t (RoundInput[103]), .B0_t (RoundKey[103]), .Z0_t (ciphertext[103]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1508 ( .A0_t (RoundInput[104]), .B0_t (RoundKey[104]), .Z0_t (ciphertext[104]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1509 ( .A0_t (RoundInput[105]), .B0_t (RoundKey[105]), .Z0_t (ciphertext[105]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1510 ( .A0_t (RoundInput[106]), .B0_t (RoundKey[106]), .Z0_t (ciphertext[106]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1511 ( .A0_t (RoundInput[107]), .B0_t (RoundKey[107]), .Z0_t (ciphertext[107]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1512 ( .A0_t (RoundInput[108]), .B0_t (RoundKey[108]), .Z0_t (ciphertext[108]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1513 ( .A0_t (RoundInput[109]), .B0_t (RoundKey[109]), .Z0_t (ciphertext[109]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1514 ( .A0_t (RoundInput[10]), .B0_t (RoundKey[10]), .Z0_t (ciphertext[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1515 ( .A0_t (RoundInput[110]), .B0_t (RoundKey[110]), .Z0_t (ciphertext[110]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1516 ( .A0_t (RoundInput[111]), .B0_t (RoundKey[111]), .Z0_t (ciphertext[111]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1517 ( .A0_t (RoundInput[112]), .B0_t (RoundKey[112]), .Z0_t (ciphertext[112]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1518 ( .A0_t (RoundInput[113]), .B0_t (RoundKey[113]), .Z0_t (ciphertext[113]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1519 ( .A0_t (RoundInput[114]), .B0_t (RoundKey[114]), .Z0_t (ciphertext[114]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1520 ( .A0_t (RoundInput[115]), .B0_t (RoundKey[115]), .Z0_t (ciphertext[115]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1521 ( .A0_t (RoundInput[116]), .B0_t (RoundKey[116]), .Z0_t (ciphertext[116]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1522 ( .A0_t (RoundInput[117]), .B0_t (RoundKey[117]), .Z0_t (ciphertext[117]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1523 ( .A0_t (RoundInput[118]), .B0_t (RoundKey[118]), .Z0_t (ciphertext[118]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1524 ( .A0_t (RoundInput[119]), .B0_t (RoundKey[119]), .Z0_t (ciphertext[119]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1525 ( .A0_t (RoundInput[11]), .B0_t (RoundKey[11]), .Z0_t (ciphertext[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1526 ( .A0_t (RoundInput[120]), .B0_t (RoundKey[120]), .Z0_t (ciphertext[120]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1527 ( .A0_t (RoundInput[121]), .B0_t (RoundKey[121]), .Z0_t (ciphertext[121]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1528 ( .A0_t (RoundInput[122]), .B0_t (RoundKey[122]), .Z0_t (ciphertext[122]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1529 ( .A0_t (RoundInput[123]), .B0_t (RoundKey[123]), .Z0_t (ciphertext[123]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1530 ( .A0_t (RoundInput[124]), .B0_t (RoundKey[124]), .Z0_t (ciphertext[124]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1531 ( .A0_t (RoundInput[125]), .B0_t (RoundKey[125]), .Z0_t (ciphertext[125]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1532 ( .A0_t (RoundInput[126]), .B0_t (RoundKey[126]), .Z0_t (ciphertext[126]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1533 ( .A0_t (RoundInput[127]), .B0_t (RoundKey[127]), .Z0_t (ciphertext[127]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1534 ( .A0_t (RoundInput[12]), .B0_t (RoundKey[12]), .Z0_t (ciphertext[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1535 ( .A0_t (RoundInput[13]), .B0_t (RoundKey[13]), .Z0_t (ciphertext[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1536 ( .A0_t (RoundInput[14]), .B0_t (RoundKey[14]), .Z0_t (ciphertext[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1537 ( .A0_t (RoundInput[15]), .B0_t (RoundKey[15]), .Z0_t (ciphertext[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1538 ( .A0_t (RoundInput[16]), .B0_t (RoundKey[16]), .Z0_t (ciphertext[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1539 ( .A0_t (RoundInput[17]), .B0_t (RoundKey[17]), .Z0_t (ciphertext[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1540 ( .A0_t (RoundInput[18]), .B0_t (RoundKey[18]), .Z0_t (ciphertext[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1541 ( .A0_t (RoundInput[19]), .B0_t (RoundKey[19]), .Z0_t (ciphertext[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1542 ( .A0_t (RoundInput[1]), .B0_t (RoundKey[1]), .Z0_t (ciphertext[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1543 ( .A0_t (RoundInput[20]), .B0_t (RoundKey[20]), .Z0_t (ciphertext[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1544 ( .A0_t (RoundInput[21]), .B0_t (RoundKey[21]), .Z0_t (ciphertext[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1545 ( .A0_t (RoundInput[22]), .B0_t (RoundKey[22]), .Z0_t (ciphertext[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1546 ( .A0_t (RoundInput[23]), .B0_t (RoundKey[23]), .Z0_t (ciphertext[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1547 ( .A0_t (RoundInput[24]), .B0_t (RoundKey[24]), .Z0_t (ciphertext[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1548 ( .A0_t (RoundInput[25]), .B0_t (RoundKey[25]), .Z0_t (ciphertext[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1549 ( .A0_t (RoundInput[26]), .B0_t (RoundKey[26]), .Z0_t (ciphertext[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1550 ( .A0_t (RoundInput[27]), .B0_t (RoundKey[27]), .Z0_t (ciphertext[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1551 ( .A0_t (RoundInput[28]), .B0_t (RoundKey[28]), .Z0_t (ciphertext[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1552 ( .A0_t (RoundInput[29]), .B0_t (RoundKey[29]), .Z0_t (ciphertext[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1553 ( .A0_t (RoundInput[2]), .B0_t (RoundKey[2]), .Z0_t (ciphertext[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1554 ( .A0_t (RoundInput[30]), .B0_t (RoundKey[30]), .Z0_t (ciphertext[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1555 ( .A0_t (RoundInput[31]), .B0_t (RoundKey[31]), .Z0_t (ciphertext[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1556 ( .A0_t (RoundInput[32]), .B0_t (RoundKey[32]), .Z0_t (ciphertext[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1557 ( .A0_t (RoundInput[33]), .B0_t (RoundKey[33]), .Z0_t (ciphertext[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1558 ( .A0_t (RoundInput[34]), .B0_t (RoundKey[34]), .Z0_t (ciphertext[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1559 ( .A0_t (RoundInput[35]), .B0_t (RoundKey[35]), .Z0_t (ciphertext[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1560 ( .A0_t (RoundInput[36]), .B0_t (RoundKey[36]), .Z0_t (ciphertext[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1561 ( .A0_t (RoundInput[37]), .B0_t (RoundKey[37]), .Z0_t (ciphertext[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1562 ( .A0_t (RoundInput[38]), .B0_t (RoundKey[38]), .Z0_t (ciphertext[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1563 ( .A0_t (RoundInput[39]), .B0_t (RoundKey[39]), .Z0_t (ciphertext[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1564 ( .A0_t (RoundInput[3]), .B0_t (RoundKey[3]), .Z0_t (ciphertext[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1565 ( .A0_t (RoundInput[40]), .B0_t (RoundKey[40]), .Z0_t (ciphertext[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1566 ( .A0_t (RoundInput[41]), .B0_t (RoundKey[41]), .Z0_t (ciphertext[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1567 ( .A0_t (RoundInput[42]), .B0_t (RoundKey[42]), .Z0_t (ciphertext[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1568 ( .A0_t (RoundInput[43]), .B0_t (RoundKey[43]), .Z0_t (ciphertext[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1569 ( .A0_t (RoundInput[44]), .B0_t (RoundKey[44]), .Z0_t (ciphertext[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1570 ( .A0_t (RoundInput[45]), .B0_t (RoundKey[45]), .Z0_t (ciphertext[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1571 ( .A0_t (RoundInput[46]), .B0_t (RoundKey[46]), .Z0_t (ciphertext[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1572 ( .A0_t (RoundInput[47]), .B0_t (RoundKey[47]), .Z0_t (ciphertext[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1573 ( .A0_t (RoundInput[48]), .B0_t (RoundKey[48]), .Z0_t (ciphertext[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1574 ( .A0_t (RoundInput[49]), .B0_t (RoundKey[49]), .Z0_t (ciphertext[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1575 ( .A0_t (RoundInput[4]), .B0_t (RoundKey[4]), .Z0_t (ciphertext[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1576 ( .A0_t (RoundInput[50]), .B0_t (RoundKey[50]), .Z0_t (ciphertext[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1577 ( .A0_t (RoundInput[51]), .B0_t (RoundKey[51]), .Z0_t (ciphertext[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1578 ( .A0_t (RoundInput[52]), .B0_t (RoundKey[52]), .Z0_t (ciphertext[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1579 ( .A0_t (RoundInput[53]), .B0_t (RoundKey[53]), .Z0_t (ciphertext[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1580 ( .A0_t (RoundInput[54]), .B0_t (RoundKey[54]), .Z0_t (ciphertext[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1581 ( .A0_t (RoundInput[55]), .B0_t (RoundKey[55]), .Z0_t (ciphertext[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1582 ( .A0_t (RoundInput[56]), .B0_t (RoundKey[56]), .Z0_t (ciphertext[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1583 ( .A0_t (RoundInput[57]), .B0_t (RoundKey[57]), .Z0_t (ciphertext[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1584 ( .A0_t (RoundInput[58]), .B0_t (RoundKey[58]), .Z0_t (ciphertext[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1585 ( .A0_t (RoundInput[59]), .B0_t (RoundKey[59]), .Z0_t (ciphertext[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1586 ( .A0_t (RoundInput[5]), .B0_t (RoundKey[5]), .Z0_t (ciphertext[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1587 ( .A0_t (RoundInput[60]), .B0_t (RoundKey[60]), .Z0_t (ciphertext[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1588 ( .A0_t (RoundInput[61]), .B0_t (RoundKey[61]), .Z0_t (ciphertext[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1589 ( .A0_t (RoundInput[62]), .B0_t (RoundKey[62]), .Z0_t (ciphertext[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1590 ( .A0_t (RoundInput[63]), .B0_t (RoundKey[63]), .Z0_t (ciphertext[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1591 ( .A0_t (RoundInput[64]), .B0_t (RoundKey[64]), .Z0_t (ciphertext[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1592 ( .A0_t (RoundInput[65]), .B0_t (RoundKey[65]), .Z0_t (ciphertext[65]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1593 ( .A0_t (RoundInput[66]), .B0_t (RoundKey[66]), .Z0_t (ciphertext[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1594 ( .A0_t (RoundInput[67]), .B0_t (RoundKey[67]), .Z0_t (ciphertext[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1595 ( .A0_t (RoundInput[68]), .B0_t (RoundKey[68]), .Z0_t (ciphertext[68]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1596 ( .A0_t (RoundInput[69]), .B0_t (RoundKey[69]), .Z0_t (ciphertext[69]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1597 ( .A0_t (RoundInput[6]), .B0_t (RoundKey[6]), .Z0_t (ciphertext[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1598 ( .A0_t (RoundInput[70]), .B0_t (RoundKey[70]), .Z0_t (ciphertext[70]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1599 ( .A0_t (RoundInput[71]), .B0_t (RoundKey[71]), .Z0_t (ciphertext[71]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1600 ( .A0_t (RoundInput[72]), .B0_t (RoundKey[72]), .Z0_t (ciphertext[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1601 ( .A0_t (RoundInput[73]), .B0_t (RoundKey[73]), .Z0_t (ciphertext[73]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1602 ( .A0_t (RoundInput[74]), .B0_t (RoundKey[74]), .Z0_t (ciphertext[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1603 ( .A0_t (RoundInput[75]), .B0_t (RoundKey[75]), .Z0_t (ciphertext[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1604 ( .A0_t (RoundInput[76]), .B0_t (RoundKey[76]), .Z0_t (ciphertext[76]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1605 ( .A0_t (RoundInput[77]), .B0_t (RoundKey[77]), .Z0_t (ciphertext[77]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1606 ( .A0_t (RoundInput[78]), .B0_t (RoundKey[78]), .Z0_t (ciphertext[78]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1607 ( .A0_t (RoundInput[79]), .B0_t (RoundKey[79]), .Z0_t (ciphertext[79]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1608 ( .A0_t (RoundInput[7]), .B0_t (RoundKey[7]), .Z0_t (ciphertext[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1609 ( .A0_t (RoundInput[80]), .B0_t (RoundKey[80]), .Z0_t (ciphertext[80]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1610 ( .A0_t (RoundInput[81]), .B0_t (RoundKey[81]), .Z0_t (ciphertext[81]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1611 ( .A0_t (RoundInput[82]), .B0_t (RoundKey[82]), .Z0_t (ciphertext[82]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1612 ( .A0_t (RoundInput[83]), .B0_t (RoundKey[83]), .Z0_t (ciphertext[83]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1613 ( .A0_t (RoundInput[84]), .B0_t (RoundKey[84]), .Z0_t (ciphertext[84]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1614 ( .A0_t (RoundInput[85]), .B0_t (RoundKey[85]), .Z0_t (ciphertext[85]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1615 ( .A0_t (RoundInput[86]), .B0_t (RoundKey[86]), .Z0_t (ciphertext[86]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1616 ( .A0_t (RoundInput[87]), .B0_t (RoundKey[87]), .Z0_t (ciphertext[87]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1617 ( .A0_t (RoundInput[88]), .B0_t (RoundKey[88]), .Z0_t (ciphertext[88]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1618 ( .A0_t (RoundInput[89]), .B0_t (RoundKey[89]), .Z0_t (ciphertext[89]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1619 ( .A0_t (RoundInput[8]), .B0_t (RoundKey[8]), .Z0_t (ciphertext[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1620 ( .A0_t (RoundInput[90]), .B0_t (RoundKey[90]), .Z0_t (ciphertext[90]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1621 ( .A0_t (RoundInput[91]), .B0_t (RoundKey[91]), .Z0_t (ciphertext[91]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1622 ( .A0_t (RoundInput[92]), .B0_t (RoundKey[92]), .Z0_t (ciphertext[92]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1623 ( .A0_t (RoundInput[93]), .B0_t (RoundKey[93]), .Z0_t (ciphertext[93]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1624 ( .A0_t (RoundInput[94]), .B0_t (RoundKey[94]), .Z0_t (ciphertext[94]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1625 ( .A0_t (RoundInput[95]), .B0_t (RoundKey[95]), .Z0_t (ciphertext[95]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1626 ( .A0_t (RoundInput[96]), .B0_t (RoundKey[96]), .Z0_t (ciphertext[96]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1627 ( .A0_t (RoundInput[97]), .B0_t (RoundKey[97]), .Z0_t (ciphertext[97]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1628 ( .A0_t (RoundInput[98]), .B0_t (RoundKey[98]), .Z0_t (ciphertext[98]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1629 ( .A0_t (RoundInput[99]), .B0_t (RoundKey[99]), .Z0_t (ciphertext[99]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1630 ( .A0_t (RoundInput[9]), .B0_t (RoundKey[9]), .Z0_t (ciphertext[9]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1631 ( .A0_t (RoundCounter[3]), .B0_t (n851), .Z0_t (n852) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1632 ( .A0_t (RoundCounter[0]), .B0_t (n852), .Z0_t (done) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U1634 ( .A0_t (RoundCounter[1]), .B0_t (RoundCounter[2]), .Z0_t (n856) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1635 ( .A0_t (n853), .B0_t (n856), .Z0_t (n283) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U1637 ( .A0_t (n855), .B0_t (n856), .Z0_t (n285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_0_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[0]), .B0_t (plaintext[0]), .Z0_t (RoundReg_Inst_ff_SDE_0_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_0_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_0_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_0_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_0_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_0_MUX_inst_Y), .B0_t (RoundOutput[0]), .Z0_t (RoundInput[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_1_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[1]), .B0_t (plaintext[1]), .Z0_t (RoundReg_Inst_ff_SDE_1_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_1_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_1_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_1_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_1_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_1_MUX_inst_Y), .B0_t (RoundOutput[1]), .Z0_t (RoundInput[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_2_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[2]), .B0_t (plaintext[2]), .Z0_t (RoundReg_Inst_ff_SDE_2_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_2_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_2_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_2_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_2_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_2_MUX_inst_Y), .B0_t (RoundOutput[2]), .Z0_t (RoundInput[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_3_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[3]), .B0_t (plaintext[3]), .Z0_t (RoundReg_Inst_ff_SDE_3_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_3_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_3_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_3_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_3_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_3_MUX_inst_Y), .B0_t (RoundOutput[3]), .Z0_t (RoundInput[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_4_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[4]), .B0_t (plaintext[4]), .Z0_t (RoundReg_Inst_ff_SDE_4_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_4_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_4_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_4_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_4_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_4_MUX_inst_Y), .B0_t (RoundOutput[4]), .Z0_t (RoundInput[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_5_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[5]), .B0_t (plaintext[5]), .Z0_t (RoundReg_Inst_ff_SDE_5_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_5_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_5_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_5_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_5_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_5_MUX_inst_Y), .B0_t (RoundOutput[5]), .Z0_t (RoundInput[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_6_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[6]), .B0_t (plaintext[6]), .Z0_t (RoundReg_Inst_ff_SDE_6_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_6_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_6_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_6_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_6_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_6_MUX_inst_Y), .B0_t (RoundOutput[6]), .Z0_t (RoundInput[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_7_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[7]), .B0_t (plaintext[7]), .Z0_t (RoundReg_Inst_ff_SDE_7_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_7_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_7_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_7_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_7_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_7_MUX_inst_Y), .B0_t (RoundOutput[7]), .Z0_t (RoundInput[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_8_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[8]), .B0_t (plaintext[8]), .Z0_t (RoundReg_Inst_ff_SDE_8_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_8_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_8_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_8_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_8_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_8_MUX_inst_Y), .B0_t (RoundOutput[8]), .Z0_t (RoundInput[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_9_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[9]), .B0_t (plaintext[9]), .Z0_t (RoundReg_Inst_ff_SDE_9_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_9_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_9_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_9_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_9_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_9_MUX_inst_Y), .B0_t (RoundOutput[9]), .Z0_t (RoundInput[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_10_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[10]), .B0_t (plaintext[10]), .Z0_t (RoundReg_Inst_ff_SDE_10_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_10_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_10_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_10_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_10_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_10_MUX_inst_Y), .B0_t (RoundOutput[10]), .Z0_t (RoundInput[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_11_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[11]), .B0_t (plaintext[11]), .Z0_t (RoundReg_Inst_ff_SDE_11_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_11_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_11_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_11_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_11_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_11_MUX_inst_Y), .B0_t (RoundOutput[11]), .Z0_t (RoundInput[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_12_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[12]), .B0_t (plaintext[12]), .Z0_t (RoundReg_Inst_ff_SDE_12_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_12_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_12_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_12_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_12_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_12_MUX_inst_Y), .B0_t (RoundOutput[12]), .Z0_t (RoundInput[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_13_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[13]), .B0_t (plaintext[13]), .Z0_t (RoundReg_Inst_ff_SDE_13_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_13_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_13_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_13_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_13_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_13_MUX_inst_Y), .B0_t (RoundOutput[13]), .Z0_t (RoundInput[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_14_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[14]), .B0_t (plaintext[14]), .Z0_t (RoundReg_Inst_ff_SDE_14_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_14_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_14_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_14_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_14_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_14_MUX_inst_Y), .B0_t (RoundOutput[14]), .Z0_t (RoundInput[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_15_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[15]), .B0_t (plaintext[15]), .Z0_t (RoundReg_Inst_ff_SDE_15_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_15_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_15_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_15_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_15_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_15_MUX_inst_Y), .B0_t (RoundOutput[15]), .Z0_t (RoundInput[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_16_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[16]), .B0_t (plaintext[16]), .Z0_t (RoundReg_Inst_ff_SDE_16_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_16_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_16_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_16_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_16_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_16_MUX_inst_Y), .B0_t (RoundOutput[16]), .Z0_t (RoundInput[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_17_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[17]), .B0_t (plaintext[17]), .Z0_t (RoundReg_Inst_ff_SDE_17_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_17_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_17_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_17_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_17_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_17_MUX_inst_Y), .B0_t (RoundOutput[17]), .Z0_t (RoundInput[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_18_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[18]), .B0_t (plaintext[18]), .Z0_t (RoundReg_Inst_ff_SDE_18_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_18_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_18_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_18_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_18_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_18_MUX_inst_Y), .B0_t (RoundOutput[18]), .Z0_t (RoundInput[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_19_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[19]), .B0_t (plaintext[19]), .Z0_t (RoundReg_Inst_ff_SDE_19_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_19_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_19_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_19_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_19_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_19_MUX_inst_Y), .B0_t (RoundOutput[19]), .Z0_t (RoundInput[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_20_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[20]), .B0_t (plaintext[20]), .Z0_t (RoundReg_Inst_ff_SDE_20_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_20_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_20_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_20_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_20_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_20_MUX_inst_Y), .B0_t (RoundOutput[20]), .Z0_t (RoundInput[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_21_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[21]), .B0_t (plaintext[21]), .Z0_t (RoundReg_Inst_ff_SDE_21_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_21_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_21_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_21_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_21_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_21_MUX_inst_Y), .B0_t (RoundOutput[21]), .Z0_t (RoundInput[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_22_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[22]), .B0_t (plaintext[22]), .Z0_t (RoundReg_Inst_ff_SDE_22_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_22_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_22_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_22_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_22_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_22_MUX_inst_Y), .B0_t (RoundOutput[22]), .Z0_t (RoundInput[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_23_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[23]), .B0_t (plaintext[23]), .Z0_t (RoundReg_Inst_ff_SDE_23_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_23_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_23_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_23_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_23_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_23_MUX_inst_Y), .B0_t (RoundOutput[23]), .Z0_t (RoundInput[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_24_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[24]), .B0_t (plaintext[24]), .Z0_t (RoundReg_Inst_ff_SDE_24_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_24_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_24_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_24_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_24_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_24_MUX_inst_Y), .B0_t (RoundOutput[24]), .Z0_t (RoundInput[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_25_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[25]), .B0_t (plaintext[25]), .Z0_t (RoundReg_Inst_ff_SDE_25_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_25_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_25_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_25_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_25_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_25_MUX_inst_Y), .B0_t (RoundOutput[25]), .Z0_t (RoundInput[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_26_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[26]), .B0_t (plaintext[26]), .Z0_t (RoundReg_Inst_ff_SDE_26_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_26_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_26_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_26_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_26_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_26_MUX_inst_Y), .B0_t (RoundOutput[26]), .Z0_t (RoundInput[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_27_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[27]), .B0_t (plaintext[27]), .Z0_t (RoundReg_Inst_ff_SDE_27_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_27_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_27_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_27_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_27_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_27_MUX_inst_Y), .B0_t (RoundOutput[27]), .Z0_t (RoundInput[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_28_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[28]), .B0_t (plaintext[28]), .Z0_t (RoundReg_Inst_ff_SDE_28_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_28_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_28_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_28_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_28_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_28_MUX_inst_Y), .B0_t (RoundOutput[28]), .Z0_t (RoundInput[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_29_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[29]), .B0_t (plaintext[29]), .Z0_t (RoundReg_Inst_ff_SDE_29_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_29_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_29_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_29_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_29_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_29_MUX_inst_Y), .B0_t (RoundOutput[29]), .Z0_t (RoundInput[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_30_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[30]), .B0_t (plaintext[30]), .Z0_t (RoundReg_Inst_ff_SDE_30_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_30_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_30_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_30_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_30_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_30_MUX_inst_Y), .B0_t (RoundOutput[30]), .Z0_t (RoundInput[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_31_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[31]), .B0_t (plaintext[31]), .Z0_t (RoundReg_Inst_ff_SDE_31_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_31_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_31_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_31_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_31_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_31_MUX_inst_Y), .B0_t (RoundOutput[31]), .Z0_t (RoundInput[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_32_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[32]), .B0_t (plaintext[32]), .Z0_t (RoundReg_Inst_ff_SDE_32_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_32_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_32_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_32_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_32_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_32_MUX_inst_Y), .B0_t (RoundOutput[32]), .Z0_t (RoundInput[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_33_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[33]), .B0_t (plaintext[33]), .Z0_t (RoundReg_Inst_ff_SDE_33_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_33_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_33_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_33_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_33_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_33_MUX_inst_Y), .B0_t (RoundOutput[33]), .Z0_t (RoundInput[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_34_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[34]), .B0_t (plaintext[34]), .Z0_t (RoundReg_Inst_ff_SDE_34_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_34_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_34_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_34_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_34_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_34_MUX_inst_Y), .B0_t (RoundOutput[34]), .Z0_t (RoundInput[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_35_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[35]), .B0_t (plaintext[35]), .Z0_t (RoundReg_Inst_ff_SDE_35_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_35_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_35_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_35_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_35_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_35_MUX_inst_Y), .B0_t (RoundOutput[35]), .Z0_t (RoundInput[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_36_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[36]), .B0_t (plaintext[36]), .Z0_t (RoundReg_Inst_ff_SDE_36_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_36_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_36_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_36_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_36_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_36_MUX_inst_Y), .B0_t (RoundOutput[36]), .Z0_t (RoundInput[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_37_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[37]), .B0_t (plaintext[37]), .Z0_t (RoundReg_Inst_ff_SDE_37_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_37_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_37_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_37_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_37_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_37_MUX_inst_Y), .B0_t (RoundOutput[37]), .Z0_t (RoundInput[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_38_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[38]), .B0_t (plaintext[38]), .Z0_t (RoundReg_Inst_ff_SDE_38_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_38_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_38_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_38_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_38_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_38_MUX_inst_Y), .B0_t (RoundOutput[38]), .Z0_t (RoundInput[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_39_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[39]), .B0_t (plaintext[39]), .Z0_t (RoundReg_Inst_ff_SDE_39_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_39_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_39_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_39_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_39_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_39_MUX_inst_Y), .B0_t (RoundOutput[39]), .Z0_t (RoundInput[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_40_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[40]), .B0_t (plaintext[40]), .Z0_t (RoundReg_Inst_ff_SDE_40_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_40_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_40_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_40_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_40_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_40_MUX_inst_Y), .B0_t (RoundOutput[40]), .Z0_t (RoundInput[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_41_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[41]), .B0_t (plaintext[41]), .Z0_t (RoundReg_Inst_ff_SDE_41_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_41_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_41_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_41_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_41_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_41_MUX_inst_Y), .B0_t (RoundOutput[41]), .Z0_t (RoundInput[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_42_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[42]), .B0_t (plaintext[42]), .Z0_t (RoundReg_Inst_ff_SDE_42_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_42_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_42_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_42_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_42_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_42_MUX_inst_Y), .B0_t (RoundOutput[42]), .Z0_t (RoundInput[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_43_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[43]), .B0_t (plaintext[43]), .Z0_t (RoundReg_Inst_ff_SDE_43_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_43_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_43_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_43_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_43_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_43_MUX_inst_Y), .B0_t (RoundOutput[43]), .Z0_t (RoundInput[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_44_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[44]), .B0_t (plaintext[44]), .Z0_t (RoundReg_Inst_ff_SDE_44_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_44_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_44_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_44_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_44_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_44_MUX_inst_Y), .B0_t (RoundOutput[44]), .Z0_t (RoundInput[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_45_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[45]), .B0_t (plaintext[45]), .Z0_t (RoundReg_Inst_ff_SDE_45_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_45_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_45_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_45_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_45_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_45_MUX_inst_Y), .B0_t (RoundOutput[45]), .Z0_t (RoundInput[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_46_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[46]), .B0_t (plaintext[46]), .Z0_t (RoundReg_Inst_ff_SDE_46_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_46_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_46_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_46_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_46_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_46_MUX_inst_Y), .B0_t (RoundOutput[46]), .Z0_t (RoundInput[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_47_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[47]), .B0_t (plaintext[47]), .Z0_t (RoundReg_Inst_ff_SDE_47_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_47_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_47_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_47_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_47_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_47_MUX_inst_Y), .B0_t (RoundOutput[47]), .Z0_t (RoundInput[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_48_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[48]), .B0_t (plaintext[48]), .Z0_t (RoundReg_Inst_ff_SDE_48_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_48_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_48_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_48_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_48_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_48_MUX_inst_Y), .B0_t (RoundOutput[48]), .Z0_t (RoundInput[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_49_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[49]), .B0_t (plaintext[49]), .Z0_t (RoundReg_Inst_ff_SDE_49_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_49_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_49_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_49_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_49_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_49_MUX_inst_Y), .B0_t (RoundOutput[49]), .Z0_t (RoundInput[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_50_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[50]), .B0_t (plaintext[50]), .Z0_t (RoundReg_Inst_ff_SDE_50_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_50_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_50_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_50_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_50_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_50_MUX_inst_Y), .B0_t (RoundOutput[50]), .Z0_t (RoundInput[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_51_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[51]), .B0_t (plaintext[51]), .Z0_t (RoundReg_Inst_ff_SDE_51_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_51_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_51_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_51_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_51_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_51_MUX_inst_Y), .B0_t (RoundOutput[51]), .Z0_t (RoundInput[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_52_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[52]), .B0_t (plaintext[52]), .Z0_t (RoundReg_Inst_ff_SDE_52_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_52_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_52_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_52_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_52_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_52_MUX_inst_Y), .B0_t (RoundOutput[52]), .Z0_t (RoundInput[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_53_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[53]), .B0_t (plaintext[53]), .Z0_t (RoundReg_Inst_ff_SDE_53_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_53_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_53_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_53_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_53_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_53_MUX_inst_Y), .B0_t (RoundOutput[53]), .Z0_t (RoundInput[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_54_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[54]), .B0_t (plaintext[54]), .Z0_t (RoundReg_Inst_ff_SDE_54_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_54_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_54_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_54_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_54_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_54_MUX_inst_Y), .B0_t (RoundOutput[54]), .Z0_t (RoundInput[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_55_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[55]), .B0_t (plaintext[55]), .Z0_t (RoundReg_Inst_ff_SDE_55_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_55_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_55_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_55_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_55_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_55_MUX_inst_Y), .B0_t (RoundOutput[55]), .Z0_t (RoundInput[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_56_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[56]), .B0_t (plaintext[56]), .Z0_t (RoundReg_Inst_ff_SDE_56_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_56_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_56_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_56_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_56_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_56_MUX_inst_Y), .B0_t (RoundOutput[56]), .Z0_t (RoundInput[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_57_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[57]), .B0_t (plaintext[57]), .Z0_t (RoundReg_Inst_ff_SDE_57_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_57_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_57_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_57_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_57_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_57_MUX_inst_Y), .B0_t (RoundOutput[57]), .Z0_t (RoundInput[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_58_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[58]), .B0_t (plaintext[58]), .Z0_t (RoundReg_Inst_ff_SDE_58_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_58_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_58_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_58_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_58_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_58_MUX_inst_Y), .B0_t (RoundOutput[58]), .Z0_t (RoundInput[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_59_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[59]), .B0_t (plaintext[59]), .Z0_t (RoundReg_Inst_ff_SDE_59_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_59_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_59_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_59_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_59_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_59_MUX_inst_Y), .B0_t (RoundOutput[59]), .Z0_t (RoundInput[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_60_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[60]), .B0_t (plaintext[60]), .Z0_t (RoundReg_Inst_ff_SDE_60_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_60_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_60_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_60_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_60_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_60_MUX_inst_Y), .B0_t (RoundOutput[60]), .Z0_t (RoundInput[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_61_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[61]), .B0_t (plaintext[61]), .Z0_t (RoundReg_Inst_ff_SDE_61_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_61_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_61_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_61_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_61_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_61_MUX_inst_Y), .B0_t (RoundOutput[61]), .Z0_t (RoundInput[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_62_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[62]), .B0_t (plaintext[62]), .Z0_t (RoundReg_Inst_ff_SDE_62_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_62_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_62_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_62_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_62_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_62_MUX_inst_Y), .B0_t (RoundOutput[62]), .Z0_t (RoundInput[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_63_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[63]), .B0_t (plaintext[63]), .Z0_t (RoundReg_Inst_ff_SDE_63_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_63_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_63_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_63_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_63_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_63_MUX_inst_Y), .B0_t (RoundOutput[63]), .Z0_t (RoundInput[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_64_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[64]), .B0_t (plaintext[64]), .Z0_t (RoundReg_Inst_ff_SDE_64_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_64_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_64_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_64_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_64_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_64_MUX_inst_Y), .B0_t (RoundOutput[64]), .Z0_t (RoundInput[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_65_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[65]), .B0_t (plaintext[65]), .Z0_t (RoundReg_Inst_ff_SDE_65_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_65_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_65_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_65_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_65_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_65_MUX_inst_Y), .B0_t (RoundOutput[65]), .Z0_t (RoundInput[65]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_66_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[66]), .B0_t (plaintext[66]), .Z0_t (RoundReg_Inst_ff_SDE_66_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_66_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_66_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_66_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_66_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_66_MUX_inst_Y), .B0_t (RoundOutput[66]), .Z0_t (RoundInput[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_67_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[67]), .B0_t (plaintext[67]), .Z0_t (RoundReg_Inst_ff_SDE_67_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_67_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_67_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_67_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_67_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_67_MUX_inst_Y), .B0_t (RoundOutput[67]), .Z0_t (RoundInput[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_68_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[68]), .B0_t (plaintext[68]), .Z0_t (RoundReg_Inst_ff_SDE_68_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_68_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_68_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_68_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_68_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_68_MUX_inst_Y), .B0_t (RoundOutput[68]), .Z0_t (RoundInput[68]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_69_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[69]), .B0_t (plaintext[69]), .Z0_t (RoundReg_Inst_ff_SDE_69_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_69_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_69_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_69_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_69_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_69_MUX_inst_Y), .B0_t (RoundOutput[69]), .Z0_t (RoundInput[69]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_70_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[70]), .B0_t (plaintext[70]), .Z0_t (RoundReg_Inst_ff_SDE_70_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_70_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_70_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_70_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_70_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_70_MUX_inst_Y), .B0_t (RoundOutput[70]), .Z0_t (RoundInput[70]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_71_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[71]), .B0_t (plaintext[71]), .Z0_t (RoundReg_Inst_ff_SDE_71_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_71_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_71_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_71_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_71_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_71_MUX_inst_Y), .B0_t (RoundOutput[71]), .Z0_t (RoundInput[71]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_72_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[72]), .B0_t (plaintext[72]), .Z0_t (RoundReg_Inst_ff_SDE_72_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_72_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_72_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_72_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_72_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_72_MUX_inst_Y), .B0_t (RoundOutput[72]), .Z0_t (RoundInput[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_73_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[73]), .B0_t (plaintext[73]), .Z0_t (RoundReg_Inst_ff_SDE_73_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_73_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_73_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_73_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_73_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_73_MUX_inst_Y), .B0_t (RoundOutput[73]), .Z0_t (RoundInput[73]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_74_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[74]), .B0_t (plaintext[74]), .Z0_t (RoundReg_Inst_ff_SDE_74_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_74_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_74_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_74_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_74_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_74_MUX_inst_Y), .B0_t (RoundOutput[74]), .Z0_t (RoundInput[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_75_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[75]), .B0_t (plaintext[75]), .Z0_t (RoundReg_Inst_ff_SDE_75_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_75_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_75_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_75_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_75_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_75_MUX_inst_Y), .B0_t (RoundOutput[75]), .Z0_t (RoundInput[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_76_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[76]), .B0_t (plaintext[76]), .Z0_t (RoundReg_Inst_ff_SDE_76_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_76_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_76_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_76_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_76_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_76_MUX_inst_Y), .B0_t (RoundOutput[76]), .Z0_t (RoundInput[76]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_77_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[77]), .B0_t (plaintext[77]), .Z0_t (RoundReg_Inst_ff_SDE_77_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_77_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_77_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_77_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_77_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_77_MUX_inst_Y), .B0_t (RoundOutput[77]), .Z0_t (RoundInput[77]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_78_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[78]), .B0_t (plaintext[78]), .Z0_t (RoundReg_Inst_ff_SDE_78_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_78_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_78_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_78_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_78_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_78_MUX_inst_Y), .B0_t (RoundOutput[78]), .Z0_t (RoundInput[78]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_79_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[79]), .B0_t (plaintext[79]), .Z0_t (RoundReg_Inst_ff_SDE_79_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_79_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_79_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_79_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_79_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_79_MUX_inst_Y), .B0_t (RoundOutput[79]), .Z0_t (RoundInput[79]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_80_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[80]), .B0_t (plaintext[80]), .Z0_t (RoundReg_Inst_ff_SDE_80_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_80_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_80_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_80_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_80_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_80_MUX_inst_Y), .B0_t (RoundOutput[80]), .Z0_t (RoundInput[80]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_81_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[81]), .B0_t (plaintext[81]), .Z0_t (RoundReg_Inst_ff_SDE_81_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_81_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_81_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_81_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_81_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_81_MUX_inst_Y), .B0_t (RoundOutput[81]), .Z0_t (RoundInput[81]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_82_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[82]), .B0_t (plaintext[82]), .Z0_t (RoundReg_Inst_ff_SDE_82_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_82_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_82_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_82_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_82_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_82_MUX_inst_Y), .B0_t (RoundOutput[82]), .Z0_t (RoundInput[82]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_83_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[83]), .B0_t (plaintext[83]), .Z0_t (RoundReg_Inst_ff_SDE_83_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_83_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_83_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_83_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_83_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_83_MUX_inst_Y), .B0_t (RoundOutput[83]), .Z0_t (RoundInput[83]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_84_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[84]), .B0_t (plaintext[84]), .Z0_t (RoundReg_Inst_ff_SDE_84_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_84_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_84_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_84_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_84_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_84_MUX_inst_Y), .B0_t (RoundOutput[84]), .Z0_t (RoundInput[84]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_85_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[85]), .B0_t (plaintext[85]), .Z0_t (RoundReg_Inst_ff_SDE_85_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_85_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_85_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_85_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_85_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_85_MUX_inst_Y), .B0_t (RoundOutput[85]), .Z0_t (RoundInput[85]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_86_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[86]), .B0_t (plaintext[86]), .Z0_t (RoundReg_Inst_ff_SDE_86_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_86_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_86_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_86_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_86_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_86_MUX_inst_Y), .B0_t (RoundOutput[86]), .Z0_t (RoundInput[86]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_87_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[87]), .B0_t (plaintext[87]), .Z0_t (RoundReg_Inst_ff_SDE_87_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_87_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_87_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_87_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_87_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_87_MUX_inst_Y), .B0_t (RoundOutput[87]), .Z0_t (RoundInput[87]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_88_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[88]), .B0_t (plaintext[88]), .Z0_t (RoundReg_Inst_ff_SDE_88_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_88_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_88_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_88_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_88_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_88_MUX_inst_Y), .B0_t (RoundOutput[88]), .Z0_t (RoundInput[88]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_89_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[89]), .B0_t (plaintext[89]), .Z0_t (RoundReg_Inst_ff_SDE_89_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_89_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_89_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_89_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_89_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_89_MUX_inst_Y), .B0_t (RoundOutput[89]), .Z0_t (RoundInput[89]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_90_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[90]), .B0_t (plaintext[90]), .Z0_t (RoundReg_Inst_ff_SDE_90_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_90_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_90_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_90_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_90_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_90_MUX_inst_Y), .B0_t (RoundOutput[90]), .Z0_t (RoundInput[90]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_91_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[91]), .B0_t (plaintext[91]), .Z0_t (RoundReg_Inst_ff_SDE_91_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_91_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_91_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_91_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_91_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_91_MUX_inst_Y), .B0_t (RoundOutput[91]), .Z0_t (RoundInput[91]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_92_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[92]), .B0_t (plaintext[92]), .Z0_t (RoundReg_Inst_ff_SDE_92_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_92_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_92_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_92_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_92_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_92_MUX_inst_Y), .B0_t (RoundOutput[92]), .Z0_t (RoundInput[92]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_93_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[93]), .B0_t (plaintext[93]), .Z0_t (RoundReg_Inst_ff_SDE_93_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_93_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_93_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_93_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_93_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_93_MUX_inst_Y), .B0_t (RoundOutput[93]), .Z0_t (RoundInput[93]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_94_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[94]), .B0_t (plaintext[94]), .Z0_t (RoundReg_Inst_ff_SDE_94_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_94_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_94_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_94_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_94_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_94_MUX_inst_Y), .B0_t (RoundOutput[94]), .Z0_t (RoundInput[94]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_95_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[95]), .B0_t (plaintext[95]), .Z0_t (RoundReg_Inst_ff_SDE_95_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_95_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_95_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_95_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_95_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_95_MUX_inst_Y), .B0_t (RoundOutput[95]), .Z0_t (RoundInput[95]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_96_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[96]), .B0_t (plaintext[96]), .Z0_t (RoundReg_Inst_ff_SDE_96_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_96_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_96_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_96_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_96_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_96_MUX_inst_Y), .B0_t (RoundOutput[96]), .Z0_t (RoundInput[96]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_97_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[97]), .B0_t (plaintext[97]), .Z0_t (RoundReg_Inst_ff_SDE_97_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_97_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_97_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_97_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_97_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_97_MUX_inst_Y), .B0_t (RoundOutput[97]), .Z0_t (RoundInput[97]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_98_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[98]), .B0_t (plaintext[98]), .Z0_t (RoundReg_Inst_ff_SDE_98_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_98_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_98_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_98_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_98_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_98_MUX_inst_Y), .B0_t (RoundOutput[98]), .Z0_t (RoundInput[98]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_99_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[99]), .B0_t (plaintext[99]), .Z0_t (RoundReg_Inst_ff_SDE_99_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_99_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_99_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_99_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_99_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_99_MUX_inst_Y), .B0_t (RoundOutput[99]), .Z0_t (RoundInput[99]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_100_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[100]), .B0_t (plaintext[100]), .Z0_t (RoundReg_Inst_ff_SDE_100_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_100_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_100_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_100_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_100_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_100_MUX_inst_Y), .B0_t (RoundOutput[100]), .Z0_t (RoundInput[100]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_101_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[101]), .B0_t (plaintext[101]), .Z0_t (RoundReg_Inst_ff_SDE_101_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_101_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_101_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_101_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_101_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_101_MUX_inst_Y), .B0_t (RoundOutput[101]), .Z0_t (RoundInput[101]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_102_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[102]), .B0_t (plaintext[102]), .Z0_t (RoundReg_Inst_ff_SDE_102_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_102_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_102_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_102_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_102_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_102_MUX_inst_Y), .B0_t (RoundOutput[102]), .Z0_t (RoundInput[102]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_103_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[103]), .B0_t (plaintext[103]), .Z0_t (RoundReg_Inst_ff_SDE_103_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_103_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_103_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_103_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_103_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_103_MUX_inst_Y), .B0_t (RoundOutput[103]), .Z0_t (RoundInput[103]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_104_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[104]), .B0_t (plaintext[104]), .Z0_t (RoundReg_Inst_ff_SDE_104_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_104_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_104_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_104_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_104_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_104_MUX_inst_Y), .B0_t (RoundOutput[104]), .Z0_t (RoundInput[104]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_105_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[105]), .B0_t (plaintext[105]), .Z0_t (RoundReg_Inst_ff_SDE_105_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_105_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_105_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_105_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_105_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_105_MUX_inst_Y), .B0_t (RoundOutput[105]), .Z0_t (RoundInput[105]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_106_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[106]), .B0_t (plaintext[106]), .Z0_t (RoundReg_Inst_ff_SDE_106_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_106_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_106_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_106_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_106_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_106_MUX_inst_Y), .B0_t (RoundOutput[106]), .Z0_t (RoundInput[106]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_107_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[107]), .B0_t (plaintext[107]), .Z0_t (RoundReg_Inst_ff_SDE_107_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_107_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_107_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_107_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_107_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_107_MUX_inst_Y), .B0_t (RoundOutput[107]), .Z0_t (RoundInput[107]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_108_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[108]), .B0_t (plaintext[108]), .Z0_t (RoundReg_Inst_ff_SDE_108_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_108_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_108_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_108_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_108_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_108_MUX_inst_Y), .B0_t (RoundOutput[108]), .Z0_t (RoundInput[108]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_109_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[109]), .B0_t (plaintext[109]), .Z0_t (RoundReg_Inst_ff_SDE_109_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_109_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_109_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_109_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_109_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_109_MUX_inst_Y), .B0_t (RoundOutput[109]), .Z0_t (RoundInput[109]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_110_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[110]), .B0_t (plaintext[110]), .Z0_t (RoundReg_Inst_ff_SDE_110_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_110_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_110_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_110_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_110_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_110_MUX_inst_Y), .B0_t (RoundOutput[110]), .Z0_t (RoundInput[110]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_111_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[111]), .B0_t (plaintext[111]), .Z0_t (RoundReg_Inst_ff_SDE_111_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_111_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_111_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_111_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_111_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_111_MUX_inst_Y), .B0_t (RoundOutput[111]), .Z0_t (RoundInput[111]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_112_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[112]), .B0_t (plaintext[112]), .Z0_t (RoundReg_Inst_ff_SDE_112_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_112_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_112_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_112_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_112_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_112_MUX_inst_Y), .B0_t (RoundOutput[112]), .Z0_t (RoundInput[112]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_113_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[113]), .B0_t (plaintext[113]), .Z0_t (RoundReg_Inst_ff_SDE_113_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_113_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_113_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_113_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_113_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_113_MUX_inst_Y), .B0_t (RoundOutput[113]), .Z0_t (RoundInput[113]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_114_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[114]), .B0_t (plaintext[114]), .Z0_t (RoundReg_Inst_ff_SDE_114_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_114_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_114_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_114_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_114_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_114_MUX_inst_Y), .B0_t (RoundOutput[114]), .Z0_t (RoundInput[114]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_115_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[115]), .B0_t (plaintext[115]), .Z0_t (RoundReg_Inst_ff_SDE_115_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_115_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_115_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_115_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_115_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_115_MUX_inst_Y), .B0_t (RoundOutput[115]), .Z0_t (RoundInput[115]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_116_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[116]), .B0_t (plaintext[116]), .Z0_t (RoundReg_Inst_ff_SDE_116_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_116_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_116_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_116_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_116_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_116_MUX_inst_Y), .B0_t (RoundOutput[116]), .Z0_t (RoundInput[116]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_117_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[117]), .B0_t (plaintext[117]), .Z0_t (RoundReg_Inst_ff_SDE_117_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_117_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_117_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_117_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_117_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_117_MUX_inst_Y), .B0_t (RoundOutput[117]), .Z0_t (RoundInput[117]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_118_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[118]), .B0_t (plaintext[118]), .Z0_t (RoundReg_Inst_ff_SDE_118_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_118_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_118_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_118_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_118_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_118_MUX_inst_Y), .B0_t (RoundOutput[118]), .Z0_t (RoundInput[118]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_119_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[119]), .B0_t (plaintext[119]), .Z0_t (RoundReg_Inst_ff_SDE_119_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_119_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_119_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_119_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_119_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_119_MUX_inst_Y), .B0_t (RoundOutput[119]), .Z0_t (RoundInput[119]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_120_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[120]), .B0_t (plaintext[120]), .Z0_t (RoundReg_Inst_ff_SDE_120_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_120_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_120_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_120_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_120_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_120_MUX_inst_Y), .B0_t (RoundOutput[120]), .Z0_t (RoundInput[120]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_121_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[121]), .B0_t (plaintext[121]), .Z0_t (RoundReg_Inst_ff_SDE_121_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_121_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_121_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_121_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_121_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_121_MUX_inst_Y), .B0_t (RoundOutput[121]), .Z0_t (RoundInput[121]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_122_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[122]), .B0_t (plaintext[122]), .Z0_t (RoundReg_Inst_ff_SDE_122_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_122_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_122_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_122_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_122_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_122_MUX_inst_Y), .B0_t (RoundOutput[122]), .Z0_t (RoundInput[122]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_123_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[123]), .B0_t (plaintext[123]), .Z0_t (RoundReg_Inst_ff_SDE_123_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_123_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_123_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_123_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_123_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_123_MUX_inst_Y), .B0_t (RoundOutput[123]), .Z0_t (RoundInput[123]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_124_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[124]), .B0_t (plaintext[124]), .Z0_t (RoundReg_Inst_ff_SDE_124_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_124_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_124_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_124_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_124_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_124_MUX_inst_Y), .B0_t (RoundOutput[124]), .Z0_t (RoundInput[124]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_125_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[125]), .B0_t (plaintext[125]), .Z0_t (RoundReg_Inst_ff_SDE_125_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_125_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_125_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_125_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_125_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_125_MUX_inst_Y), .B0_t (RoundOutput[125]), .Z0_t (RoundInput[125]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_126_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[126]), .B0_t (plaintext[126]), .Z0_t (RoundReg_Inst_ff_SDE_126_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_126_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_126_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_126_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_126_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_126_MUX_inst_Y), .B0_t (RoundOutput[126]), .Z0_t (RoundInput[126]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_127_MUX_inst_XOR1_U1 ( .A0_t (RoundOutput[127]), .B0_t (plaintext[127]), .Z0_t (RoundReg_Inst_ff_SDE_127_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) RoundReg_Inst_ff_SDE_127_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (RoundReg_Inst_ff_SDE_127_MUX_inst_X), .Z0_t (RoundReg_Inst_ff_SDE_127_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) RoundReg_Inst_ff_SDE_127_MUX_inst_XOR2_U1 ( .A0_t (RoundReg_Inst_ff_SDE_127_MUX_inst_Y), .B0_t (RoundOutput[127]), .Z0_t (RoundInput[127]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .A0_t (ciphertext[7]), .B0_t (ciphertext[4]), .Z0_t (SubBytesIns_Inst_Sbox_0_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .A0_t (ciphertext[7]), .B0_t (ciphertext[2]), .Z0_t (SubBytesIns_Inst_Sbox_0_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .A0_t (ciphertext[7]), .B0_t (ciphertext[1]), .Z0_t (SubBytesIns_Inst_Sbox_0_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .A0_t (ciphertext[4]), .B0_t (ciphertext[2]), .Z0_t (SubBytesIns_Inst_Sbox_0_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .A0_t (ciphertext[3]), .B0_t (ciphertext[1]), .Z0_t (SubBytesIns_Inst_Sbox_0_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T1), .B0_t (SubBytesIns_Inst_Sbox_0_T5), .Z0_t (SubBytesIns_Inst_Sbox_0_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .A0_t (ciphertext[6]), .B0_t (ciphertext[5]), .Z0_t (SubBytesIns_Inst_Sbox_0_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .A0_t (ciphertext[0]), .B0_t (SubBytesIns_Inst_Sbox_0_T6), .Z0_t (SubBytesIns_Inst_Sbox_0_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .A0_t (ciphertext[0]), .B0_t (SubBytesIns_Inst_Sbox_0_T7), .Z0_t (SubBytesIns_Inst_Sbox_0_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T6), .B0_t (SubBytesIns_Inst_Sbox_0_T7), .Z0_t (SubBytesIns_Inst_Sbox_0_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .A0_t (ciphertext[6]), .B0_t (ciphertext[2]), .Z0_t (SubBytesIns_Inst_Sbox_0_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .A0_t (ciphertext[5]), .B0_t (ciphertext[2]), .Z0_t (SubBytesIns_Inst_Sbox_0_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T3), .B0_t (SubBytesIns_Inst_Sbox_0_T4), .Z0_t (SubBytesIns_Inst_Sbox_0_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T6), .B0_t (SubBytesIns_Inst_Sbox_0_T11), .Z0_t (SubBytesIns_Inst_Sbox_0_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T5), .B0_t (SubBytesIns_Inst_Sbox_0_T11), .Z0_t (SubBytesIns_Inst_Sbox_0_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T5), .B0_t (SubBytesIns_Inst_Sbox_0_T12), .Z0_t (SubBytesIns_Inst_Sbox_0_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T9), .B0_t (SubBytesIns_Inst_Sbox_0_T16), .Z0_t (SubBytesIns_Inst_Sbox_0_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .A0_t (ciphertext[4]), .B0_t (ciphertext[0]), .Z0_t (SubBytesIns_Inst_Sbox_0_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T7), .B0_t (SubBytesIns_Inst_Sbox_0_T18), .Z0_t (SubBytesIns_Inst_Sbox_0_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T1), .B0_t (SubBytesIns_Inst_Sbox_0_T19), .Z0_t (SubBytesIns_Inst_Sbox_0_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .A0_t (ciphertext[1]), .B0_t (ciphertext[0]), .Z0_t (SubBytesIns_Inst_Sbox_0_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T7), .B0_t (SubBytesIns_Inst_Sbox_0_T21), .Z0_t (SubBytesIns_Inst_Sbox_0_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T2), .B0_t (SubBytesIns_Inst_Sbox_0_T22), .Z0_t (SubBytesIns_Inst_Sbox_0_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T2), .B0_t (SubBytesIns_Inst_Sbox_0_T10), .Z0_t (SubBytesIns_Inst_Sbox_0_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T20), .B0_t (SubBytesIns_Inst_Sbox_0_T17), .Z0_t (SubBytesIns_Inst_Sbox_0_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T3), .B0_t (SubBytesIns_Inst_Sbox_0_T16), .Z0_t (SubBytesIns_Inst_Sbox_0_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T1), .B0_t (SubBytesIns_Inst_Sbox_0_T12), .Z0_t (SubBytesIns_Inst_Sbox_0_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T13), .B0_t (SubBytesIns_Inst_Sbox_0_T6), .Z0_t (SubBytesIns_Inst_Sbox_0_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T23), .B0_t (SubBytesIns_Inst_Sbox_0_T8), .Z0_t (SubBytesIns_Inst_Sbox_0_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T14), .B0_t (SubBytesIns_Inst_Sbox_0_M1), .Z0_t (SubBytesIns_Inst_Sbox_0_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T19), .B0_t (ciphertext[0]), .Z0_t (SubBytesIns_Inst_Sbox_0_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M4), .B0_t (SubBytesIns_Inst_Sbox_0_M1), .Z0_t (SubBytesIns_Inst_Sbox_0_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T3), .B0_t (SubBytesIns_Inst_Sbox_0_T16), .Z0_t (SubBytesIns_Inst_Sbox_0_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T22), .B0_t (SubBytesIns_Inst_Sbox_0_T9), .Z0_t (SubBytesIns_Inst_Sbox_0_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T26), .B0_t (SubBytesIns_Inst_Sbox_0_M6), .Z0_t (SubBytesIns_Inst_Sbox_0_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T20), .B0_t (SubBytesIns_Inst_Sbox_0_T17), .Z0_t (SubBytesIns_Inst_Sbox_0_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M9), .B0_t (SubBytesIns_Inst_Sbox_0_M6), .Z0_t (SubBytesIns_Inst_Sbox_0_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T1), .B0_t (SubBytesIns_Inst_Sbox_0_T15), .Z0_t (SubBytesIns_Inst_Sbox_0_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T4), .B0_t (SubBytesIns_Inst_Sbox_0_T27), .Z0_t (SubBytesIns_Inst_Sbox_0_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M12), .B0_t (SubBytesIns_Inst_Sbox_0_M11), .Z0_t (SubBytesIns_Inst_Sbox_0_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_T2), .B0_t (SubBytesIns_Inst_Sbox_0_T10), .Z0_t (SubBytesIns_Inst_Sbox_0_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M14), .B0_t (SubBytesIns_Inst_Sbox_0_M11), .Z0_t (SubBytesIns_Inst_Sbox_0_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M3), .B0_t (SubBytesIns_Inst_Sbox_0_M2), .Z0_t (SubBytesIns_Inst_Sbox_0_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M5), .B0_t (SubBytesIns_Inst_Sbox_0_T24), .Z0_t (SubBytesIns_Inst_Sbox_0_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M8), .B0_t (SubBytesIns_Inst_Sbox_0_M7), .Z0_t (SubBytesIns_Inst_Sbox_0_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M10), .B0_t (SubBytesIns_Inst_Sbox_0_M15), .Z0_t (SubBytesIns_Inst_Sbox_0_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M16), .B0_t (SubBytesIns_Inst_Sbox_0_M13), .Z0_t (SubBytesIns_Inst_Sbox_0_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M17), .B0_t (SubBytesIns_Inst_Sbox_0_M15), .Z0_t (SubBytesIns_Inst_Sbox_0_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M18), .B0_t (SubBytesIns_Inst_Sbox_0_M13), .Z0_t (SubBytesIns_Inst_Sbox_0_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M19), .B0_t (SubBytesIns_Inst_Sbox_0_T25), .Z0_t (SubBytesIns_Inst_Sbox_0_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M22), .B0_t (SubBytesIns_Inst_Sbox_0_M23), .Z0_t (SubBytesIns_Inst_Sbox_0_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M22), .B0_t (SubBytesIns_Inst_Sbox_0_M20), .Z0_t (SubBytesIns_Inst_Sbox_0_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M21), .B0_t (SubBytesIns_Inst_Sbox_0_M25), .Z0_t (SubBytesIns_Inst_Sbox_0_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M20), .B0_t (SubBytesIns_Inst_Sbox_0_M21), .Z0_t (SubBytesIns_Inst_Sbox_0_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M23), .B0_t (SubBytesIns_Inst_Sbox_0_M25), .Z0_t (SubBytesIns_Inst_Sbox_0_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M28), .B0_t (SubBytesIns_Inst_Sbox_0_M27), .Z0_t (SubBytesIns_Inst_Sbox_0_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M26), .B0_t (SubBytesIns_Inst_Sbox_0_M24), .Z0_t (SubBytesIns_Inst_Sbox_0_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M20), .B0_t (SubBytesIns_Inst_Sbox_0_M23), .Z0_t (SubBytesIns_Inst_Sbox_0_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M27), .B0_t (SubBytesIns_Inst_Sbox_0_M31), .Z0_t (SubBytesIns_Inst_Sbox_0_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M27), .B0_t (SubBytesIns_Inst_Sbox_0_M25), .Z0_t (SubBytesIns_Inst_Sbox_0_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M21), .B0_t (SubBytesIns_Inst_Sbox_0_M22), .Z0_t (SubBytesIns_Inst_Sbox_0_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M24), .B0_t (SubBytesIns_Inst_Sbox_0_M34), .Z0_t (SubBytesIns_Inst_Sbox_0_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M24), .B0_t (SubBytesIns_Inst_Sbox_0_M25), .Z0_t (SubBytesIns_Inst_Sbox_0_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M21), .B0_t (SubBytesIns_Inst_Sbox_0_M29), .Z0_t (SubBytesIns_Inst_Sbox_0_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M32), .B0_t (SubBytesIns_Inst_Sbox_0_M33), .Z0_t (SubBytesIns_Inst_Sbox_0_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M23), .B0_t (SubBytesIns_Inst_Sbox_0_M30), .Z0_t (SubBytesIns_Inst_Sbox_0_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M35), .B0_t (SubBytesIns_Inst_Sbox_0_M36), .Z0_t (SubBytesIns_Inst_Sbox_0_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M38), .B0_t (SubBytesIns_Inst_Sbox_0_M40), .Z0_t (SubBytesIns_Inst_Sbox_0_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M37), .B0_t (SubBytesIns_Inst_Sbox_0_M39), .Z0_t (SubBytesIns_Inst_Sbox_0_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M37), .B0_t (SubBytesIns_Inst_Sbox_0_M38), .Z0_t (SubBytesIns_Inst_Sbox_0_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M39), .B0_t (SubBytesIns_Inst_Sbox_0_M40), .Z0_t (SubBytesIns_Inst_Sbox_0_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M42), .B0_t (SubBytesIns_Inst_Sbox_0_M41), .Z0_t (SubBytesIns_Inst_Sbox_0_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M44), .B0_t (SubBytesIns_Inst_Sbox_0_T6), .Z0_t (SubBytesIns_Inst_Sbox_0_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M40), .B0_t (SubBytesIns_Inst_Sbox_0_T8), .Z0_t (SubBytesIns_Inst_Sbox_0_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M39), .B0_t (ciphertext[0]), .Z0_t (SubBytesIns_Inst_Sbox_0_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M43), .B0_t (SubBytesIns_Inst_Sbox_0_T16), .Z0_t (SubBytesIns_Inst_Sbox_0_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M38), .B0_t (SubBytesIns_Inst_Sbox_0_T9), .Z0_t (SubBytesIns_Inst_Sbox_0_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M37), .B0_t (SubBytesIns_Inst_Sbox_0_T17), .Z0_t (SubBytesIns_Inst_Sbox_0_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M42), .B0_t (SubBytesIns_Inst_Sbox_0_T15), .Z0_t (SubBytesIns_Inst_Sbox_0_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M45), .B0_t (SubBytesIns_Inst_Sbox_0_T27), .Z0_t (SubBytesIns_Inst_Sbox_0_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M41), .B0_t (SubBytesIns_Inst_Sbox_0_T10), .Z0_t (SubBytesIns_Inst_Sbox_0_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M44), .B0_t (SubBytesIns_Inst_Sbox_0_T13), .Z0_t (SubBytesIns_Inst_Sbox_0_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M40), .B0_t (SubBytesIns_Inst_Sbox_0_T23), .Z0_t (SubBytesIns_Inst_Sbox_0_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M39), .B0_t (SubBytesIns_Inst_Sbox_0_T19), .Z0_t (SubBytesIns_Inst_Sbox_0_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M43), .B0_t (SubBytesIns_Inst_Sbox_0_T3), .Z0_t (SubBytesIns_Inst_Sbox_0_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M38), .B0_t (SubBytesIns_Inst_Sbox_0_T22), .Z0_t (SubBytesIns_Inst_Sbox_0_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M37), .B0_t (SubBytesIns_Inst_Sbox_0_T20), .Z0_t (SubBytesIns_Inst_Sbox_0_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M42), .B0_t (SubBytesIns_Inst_Sbox_0_T1), .Z0_t (SubBytesIns_Inst_Sbox_0_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M45), .B0_t (SubBytesIns_Inst_Sbox_0_T4), .Z0_t (SubBytesIns_Inst_Sbox_0_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M41), .B0_t (SubBytesIns_Inst_Sbox_0_T2), .Z0_t (SubBytesIns_Inst_Sbox_0_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M61), .B0_t (SubBytesIns_Inst_Sbox_0_M62), .Z0_t (SubBytesIns_Inst_Sbox_0_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M50), .B0_t (SubBytesIns_Inst_Sbox_0_M56), .Z0_t (SubBytesIns_Inst_Sbox_0_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M46), .B0_t (SubBytesIns_Inst_Sbox_0_M48), .Z0_t (SubBytesIns_Inst_Sbox_0_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M47), .B0_t (SubBytesIns_Inst_Sbox_0_M55), .Z0_t (SubBytesIns_Inst_Sbox_0_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M54), .B0_t (SubBytesIns_Inst_Sbox_0_M58), .Z0_t (SubBytesIns_Inst_Sbox_0_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M49), .B0_t (SubBytesIns_Inst_Sbox_0_M61), .Z0_t (SubBytesIns_Inst_Sbox_0_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M62), .B0_t (SubBytesIns_Inst_Sbox_0_L5), .Z0_t (SubBytesIns_Inst_Sbox_0_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M46), .B0_t (SubBytesIns_Inst_Sbox_0_L3), .Z0_t (SubBytesIns_Inst_Sbox_0_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M51), .B0_t (SubBytesIns_Inst_Sbox_0_M59), .Z0_t (SubBytesIns_Inst_Sbox_0_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M52), .B0_t (SubBytesIns_Inst_Sbox_0_M53), .Z0_t (SubBytesIns_Inst_Sbox_0_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M53), .B0_t (SubBytesIns_Inst_Sbox_0_L4), .Z0_t (SubBytesIns_Inst_Sbox_0_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M60), .B0_t (SubBytesIns_Inst_Sbox_0_L2), .Z0_t (SubBytesIns_Inst_Sbox_0_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M48), .B0_t (SubBytesIns_Inst_Sbox_0_M51), .Z0_t (SubBytesIns_Inst_Sbox_0_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M50), .B0_t (SubBytesIns_Inst_Sbox_0_L0), .Z0_t (SubBytesIns_Inst_Sbox_0_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M52), .B0_t (SubBytesIns_Inst_Sbox_0_M61), .Z0_t (SubBytesIns_Inst_Sbox_0_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M55), .B0_t (SubBytesIns_Inst_Sbox_0_L1), .Z0_t (SubBytesIns_Inst_Sbox_0_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M56), .B0_t (SubBytesIns_Inst_Sbox_0_L0), .Z0_t (SubBytesIns_Inst_Sbox_0_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M57), .B0_t (SubBytesIns_Inst_Sbox_0_L1), .Z0_t (SubBytesIns_Inst_Sbox_0_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M58), .B0_t (SubBytesIns_Inst_Sbox_0_L8), .Z0_t (SubBytesIns_Inst_Sbox_0_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_M63), .B0_t (SubBytesIns_Inst_Sbox_0_L4), .Z0_t (SubBytesIns_Inst_Sbox_0_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L0), .B0_t (SubBytesIns_Inst_Sbox_0_L1), .Z0_t (SubBytesIns_Inst_Sbox_0_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L1), .B0_t (SubBytesIns_Inst_Sbox_0_L7), .Z0_t (SubBytesIns_Inst_Sbox_0_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L3), .B0_t (SubBytesIns_Inst_Sbox_0_L12), .Z0_t (SubBytesIns_Inst_Sbox_0_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L18), .B0_t (SubBytesIns_Inst_Sbox_0_L2), .Z0_t (SubBytesIns_Inst_Sbox_0_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L15), .B0_t (SubBytesIns_Inst_Sbox_0_L9), .Z0_t (SubBytesIns_Inst_Sbox_0_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L6), .B0_t (SubBytesIns_Inst_Sbox_0_L10), .Z0_t (SubBytesIns_Inst_Sbox_0_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L7), .B0_t (SubBytesIns_Inst_Sbox_0_L9), .Z0_t (SubBytesIns_Inst_Sbox_0_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L8), .B0_t (SubBytesIns_Inst_Sbox_0_L10), .Z0_t (SubBytesIns_Inst_Sbox_0_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L11), .B0_t (SubBytesIns_Inst_Sbox_0_L14), .Z0_t (SubBytesIns_Inst_Sbox_0_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L11), .B0_t (SubBytesIns_Inst_Sbox_0_L17), .Z0_t (SubBytesIns_Inst_Sbox_0_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L6), .B0_t (SubBytesIns_Inst_Sbox_0_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L16), .B0_t (SubBytesIns_Inst_Sbox_0_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L19), .B0_t (SubBytesIns_Inst_Sbox_0_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L6), .B0_t (SubBytesIns_Inst_Sbox_0_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L20), .B0_t (SubBytesIns_Inst_Sbox_0_L22), .Z0_t (MixColumnsInput[99]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L25), .B0_t (SubBytesIns_Inst_Sbox_0_L29), .Z0_t (MixColumnsInput[98]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L13), .B0_t (SubBytesIns_Inst_Sbox_0_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_0_L6), .B0_t (SubBytesIns_Inst_Sbox_0_L23), .Z0_t (MixColumnsInput[96]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .A0_t (ciphertext[15]), .B0_t (ciphertext[12]), .Z0_t (SubBytesIns_Inst_Sbox_1_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .A0_t (ciphertext[15]), .B0_t (ciphertext[10]), .Z0_t (SubBytesIns_Inst_Sbox_1_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .A0_t (ciphertext[15]), .B0_t (ciphertext[9]), .Z0_t (SubBytesIns_Inst_Sbox_1_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .A0_t (ciphertext[12]), .B0_t (ciphertext[10]), .Z0_t (SubBytesIns_Inst_Sbox_1_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .A0_t (ciphertext[11]), .B0_t (ciphertext[9]), .Z0_t (SubBytesIns_Inst_Sbox_1_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T1), .B0_t (SubBytesIns_Inst_Sbox_1_T5), .Z0_t (SubBytesIns_Inst_Sbox_1_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .A0_t (ciphertext[14]), .B0_t (ciphertext[13]), .Z0_t (SubBytesIns_Inst_Sbox_1_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .A0_t (ciphertext[8]), .B0_t (SubBytesIns_Inst_Sbox_1_T6), .Z0_t (SubBytesIns_Inst_Sbox_1_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .A0_t (ciphertext[8]), .B0_t (SubBytesIns_Inst_Sbox_1_T7), .Z0_t (SubBytesIns_Inst_Sbox_1_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T6), .B0_t (SubBytesIns_Inst_Sbox_1_T7), .Z0_t (SubBytesIns_Inst_Sbox_1_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .A0_t (ciphertext[14]), .B0_t (ciphertext[10]), .Z0_t (SubBytesIns_Inst_Sbox_1_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .A0_t (ciphertext[13]), .B0_t (ciphertext[10]), .Z0_t (SubBytesIns_Inst_Sbox_1_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T3), .B0_t (SubBytesIns_Inst_Sbox_1_T4), .Z0_t (SubBytesIns_Inst_Sbox_1_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T6), .B0_t (SubBytesIns_Inst_Sbox_1_T11), .Z0_t (SubBytesIns_Inst_Sbox_1_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T5), .B0_t (SubBytesIns_Inst_Sbox_1_T11), .Z0_t (SubBytesIns_Inst_Sbox_1_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T5), .B0_t (SubBytesIns_Inst_Sbox_1_T12), .Z0_t (SubBytesIns_Inst_Sbox_1_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T9), .B0_t (SubBytesIns_Inst_Sbox_1_T16), .Z0_t (SubBytesIns_Inst_Sbox_1_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .A0_t (ciphertext[12]), .B0_t (ciphertext[8]), .Z0_t (SubBytesIns_Inst_Sbox_1_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T7), .B0_t (SubBytesIns_Inst_Sbox_1_T18), .Z0_t (SubBytesIns_Inst_Sbox_1_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T1), .B0_t (SubBytesIns_Inst_Sbox_1_T19), .Z0_t (SubBytesIns_Inst_Sbox_1_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .A0_t (ciphertext[9]), .B0_t (ciphertext[8]), .Z0_t (SubBytesIns_Inst_Sbox_1_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T7), .B0_t (SubBytesIns_Inst_Sbox_1_T21), .Z0_t (SubBytesIns_Inst_Sbox_1_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T2), .B0_t (SubBytesIns_Inst_Sbox_1_T22), .Z0_t (SubBytesIns_Inst_Sbox_1_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T2), .B0_t (SubBytesIns_Inst_Sbox_1_T10), .Z0_t (SubBytesIns_Inst_Sbox_1_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T20), .B0_t (SubBytesIns_Inst_Sbox_1_T17), .Z0_t (SubBytesIns_Inst_Sbox_1_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T3), .B0_t (SubBytesIns_Inst_Sbox_1_T16), .Z0_t (SubBytesIns_Inst_Sbox_1_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T1), .B0_t (SubBytesIns_Inst_Sbox_1_T12), .Z0_t (SubBytesIns_Inst_Sbox_1_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T13), .B0_t (SubBytesIns_Inst_Sbox_1_T6), .Z0_t (SubBytesIns_Inst_Sbox_1_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T23), .B0_t (SubBytesIns_Inst_Sbox_1_T8), .Z0_t (SubBytesIns_Inst_Sbox_1_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T14), .B0_t (SubBytesIns_Inst_Sbox_1_M1), .Z0_t (SubBytesIns_Inst_Sbox_1_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T19), .B0_t (ciphertext[8]), .Z0_t (SubBytesIns_Inst_Sbox_1_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M4), .B0_t (SubBytesIns_Inst_Sbox_1_M1), .Z0_t (SubBytesIns_Inst_Sbox_1_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T3), .B0_t (SubBytesIns_Inst_Sbox_1_T16), .Z0_t (SubBytesIns_Inst_Sbox_1_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T22), .B0_t (SubBytesIns_Inst_Sbox_1_T9), .Z0_t (SubBytesIns_Inst_Sbox_1_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T26), .B0_t (SubBytesIns_Inst_Sbox_1_M6), .Z0_t (SubBytesIns_Inst_Sbox_1_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T20), .B0_t (SubBytesIns_Inst_Sbox_1_T17), .Z0_t (SubBytesIns_Inst_Sbox_1_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M9), .B0_t (SubBytesIns_Inst_Sbox_1_M6), .Z0_t (SubBytesIns_Inst_Sbox_1_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T1), .B0_t (SubBytesIns_Inst_Sbox_1_T15), .Z0_t (SubBytesIns_Inst_Sbox_1_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T4), .B0_t (SubBytesIns_Inst_Sbox_1_T27), .Z0_t (SubBytesIns_Inst_Sbox_1_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M12), .B0_t (SubBytesIns_Inst_Sbox_1_M11), .Z0_t (SubBytesIns_Inst_Sbox_1_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_T2), .B0_t (SubBytesIns_Inst_Sbox_1_T10), .Z0_t (SubBytesIns_Inst_Sbox_1_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M14), .B0_t (SubBytesIns_Inst_Sbox_1_M11), .Z0_t (SubBytesIns_Inst_Sbox_1_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M3), .B0_t (SubBytesIns_Inst_Sbox_1_M2), .Z0_t (SubBytesIns_Inst_Sbox_1_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M5), .B0_t (SubBytesIns_Inst_Sbox_1_T24), .Z0_t (SubBytesIns_Inst_Sbox_1_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M8), .B0_t (SubBytesIns_Inst_Sbox_1_M7), .Z0_t (SubBytesIns_Inst_Sbox_1_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M10), .B0_t (SubBytesIns_Inst_Sbox_1_M15), .Z0_t (SubBytesIns_Inst_Sbox_1_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M16), .B0_t (SubBytesIns_Inst_Sbox_1_M13), .Z0_t (SubBytesIns_Inst_Sbox_1_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M17), .B0_t (SubBytesIns_Inst_Sbox_1_M15), .Z0_t (SubBytesIns_Inst_Sbox_1_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M18), .B0_t (SubBytesIns_Inst_Sbox_1_M13), .Z0_t (SubBytesIns_Inst_Sbox_1_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M19), .B0_t (SubBytesIns_Inst_Sbox_1_T25), .Z0_t (SubBytesIns_Inst_Sbox_1_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M22), .B0_t (SubBytesIns_Inst_Sbox_1_M23), .Z0_t (SubBytesIns_Inst_Sbox_1_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M22), .B0_t (SubBytesIns_Inst_Sbox_1_M20), .Z0_t (SubBytesIns_Inst_Sbox_1_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M21), .B0_t (SubBytesIns_Inst_Sbox_1_M25), .Z0_t (SubBytesIns_Inst_Sbox_1_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M20), .B0_t (SubBytesIns_Inst_Sbox_1_M21), .Z0_t (SubBytesIns_Inst_Sbox_1_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M23), .B0_t (SubBytesIns_Inst_Sbox_1_M25), .Z0_t (SubBytesIns_Inst_Sbox_1_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M28), .B0_t (SubBytesIns_Inst_Sbox_1_M27), .Z0_t (SubBytesIns_Inst_Sbox_1_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M26), .B0_t (SubBytesIns_Inst_Sbox_1_M24), .Z0_t (SubBytesIns_Inst_Sbox_1_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M20), .B0_t (SubBytesIns_Inst_Sbox_1_M23), .Z0_t (SubBytesIns_Inst_Sbox_1_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M27), .B0_t (SubBytesIns_Inst_Sbox_1_M31), .Z0_t (SubBytesIns_Inst_Sbox_1_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M27), .B0_t (SubBytesIns_Inst_Sbox_1_M25), .Z0_t (SubBytesIns_Inst_Sbox_1_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M21), .B0_t (SubBytesIns_Inst_Sbox_1_M22), .Z0_t (SubBytesIns_Inst_Sbox_1_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M24), .B0_t (SubBytesIns_Inst_Sbox_1_M34), .Z0_t (SubBytesIns_Inst_Sbox_1_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M24), .B0_t (SubBytesIns_Inst_Sbox_1_M25), .Z0_t (SubBytesIns_Inst_Sbox_1_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M21), .B0_t (SubBytesIns_Inst_Sbox_1_M29), .Z0_t (SubBytesIns_Inst_Sbox_1_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M32), .B0_t (SubBytesIns_Inst_Sbox_1_M33), .Z0_t (SubBytesIns_Inst_Sbox_1_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M23), .B0_t (SubBytesIns_Inst_Sbox_1_M30), .Z0_t (SubBytesIns_Inst_Sbox_1_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M35), .B0_t (SubBytesIns_Inst_Sbox_1_M36), .Z0_t (SubBytesIns_Inst_Sbox_1_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M38), .B0_t (SubBytesIns_Inst_Sbox_1_M40), .Z0_t (SubBytesIns_Inst_Sbox_1_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M37), .B0_t (SubBytesIns_Inst_Sbox_1_M39), .Z0_t (SubBytesIns_Inst_Sbox_1_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M37), .B0_t (SubBytesIns_Inst_Sbox_1_M38), .Z0_t (SubBytesIns_Inst_Sbox_1_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M39), .B0_t (SubBytesIns_Inst_Sbox_1_M40), .Z0_t (SubBytesIns_Inst_Sbox_1_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M42), .B0_t (SubBytesIns_Inst_Sbox_1_M41), .Z0_t (SubBytesIns_Inst_Sbox_1_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M44), .B0_t (SubBytesIns_Inst_Sbox_1_T6), .Z0_t (SubBytesIns_Inst_Sbox_1_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M40), .B0_t (SubBytesIns_Inst_Sbox_1_T8), .Z0_t (SubBytesIns_Inst_Sbox_1_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M39), .B0_t (ciphertext[8]), .Z0_t (SubBytesIns_Inst_Sbox_1_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M43), .B0_t (SubBytesIns_Inst_Sbox_1_T16), .Z0_t (SubBytesIns_Inst_Sbox_1_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M38), .B0_t (SubBytesIns_Inst_Sbox_1_T9), .Z0_t (SubBytesIns_Inst_Sbox_1_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M37), .B0_t (SubBytesIns_Inst_Sbox_1_T17), .Z0_t (SubBytesIns_Inst_Sbox_1_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M42), .B0_t (SubBytesIns_Inst_Sbox_1_T15), .Z0_t (SubBytesIns_Inst_Sbox_1_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M45), .B0_t (SubBytesIns_Inst_Sbox_1_T27), .Z0_t (SubBytesIns_Inst_Sbox_1_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M41), .B0_t (SubBytesIns_Inst_Sbox_1_T10), .Z0_t (SubBytesIns_Inst_Sbox_1_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M44), .B0_t (SubBytesIns_Inst_Sbox_1_T13), .Z0_t (SubBytesIns_Inst_Sbox_1_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M40), .B0_t (SubBytesIns_Inst_Sbox_1_T23), .Z0_t (SubBytesIns_Inst_Sbox_1_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M39), .B0_t (SubBytesIns_Inst_Sbox_1_T19), .Z0_t (SubBytesIns_Inst_Sbox_1_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M43), .B0_t (SubBytesIns_Inst_Sbox_1_T3), .Z0_t (SubBytesIns_Inst_Sbox_1_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M38), .B0_t (SubBytesIns_Inst_Sbox_1_T22), .Z0_t (SubBytesIns_Inst_Sbox_1_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M37), .B0_t (SubBytesIns_Inst_Sbox_1_T20), .Z0_t (SubBytesIns_Inst_Sbox_1_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M42), .B0_t (SubBytesIns_Inst_Sbox_1_T1), .Z0_t (SubBytesIns_Inst_Sbox_1_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M45), .B0_t (SubBytesIns_Inst_Sbox_1_T4), .Z0_t (SubBytesIns_Inst_Sbox_1_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M41), .B0_t (SubBytesIns_Inst_Sbox_1_T2), .Z0_t (SubBytesIns_Inst_Sbox_1_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M61), .B0_t (SubBytesIns_Inst_Sbox_1_M62), .Z0_t (SubBytesIns_Inst_Sbox_1_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M50), .B0_t (SubBytesIns_Inst_Sbox_1_M56), .Z0_t (SubBytesIns_Inst_Sbox_1_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M46), .B0_t (SubBytesIns_Inst_Sbox_1_M48), .Z0_t (SubBytesIns_Inst_Sbox_1_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M47), .B0_t (SubBytesIns_Inst_Sbox_1_M55), .Z0_t (SubBytesIns_Inst_Sbox_1_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M54), .B0_t (SubBytesIns_Inst_Sbox_1_M58), .Z0_t (SubBytesIns_Inst_Sbox_1_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M49), .B0_t (SubBytesIns_Inst_Sbox_1_M61), .Z0_t (SubBytesIns_Inst_Sbox_1_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M62), .B0_t (SubBytesIns_Inst_Sbox_1_L5), .Z0_t (SubBytesIns_Inst_Sbox_1_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M46), .B0_t (SubBytesIns_Inst_Sbox_1_L3), .Z0_t (SubBytesIns_Inst_Sbox_1_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M51), .B0_t (SubBytesIns_Inst_Sbox_1_M59), .Z0_t (SubBytesIns_Inst_Sbox_1_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M52), .B0_t (SubBytesIns_Inst_Sbox_1_M53), .Z0_t (SubBytesIns_Inst_Sbox_1_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M53), .B0_t (SubBytesIns_Inst_Sbox_1_L4), .Z0_t (SubBytesIns_Inst_Sbox_1_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M60), .B0_t (SubBytesIns_Inst_Sbox_1_L2), .Z0_t (SubBytesIns_Inst_Sbox_1_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M48), .B0_t (SubBytesIns_Inst_Sbox_1_M51), .Z0_t (SubBytesIns_Inst_Sbox_1_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M50), .B0_t (SubBytesIns_Inst_Sbox_1_L0), .Z0_t (SubBytesIns_Inst_Sbox_1_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M52), .B0_t (SubBytesIns_Inst_Sbox_1_M61), .Z0_t (SubBytesIns_Inst_Sbox_1_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M55), .B0_t (SubBytesIns_Inst_Sbox_1_L1), .Z0_t (SubBytesIns_Inst_Sbox_1_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M56), .B0_t (SubBytesIns_Inst_Sbox_1_L0), .Z0_t (SubBytesIns_Inst_Sbox_1_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M57), .B0_t (SubBytesIns_Inst_Sbox_1_L1), .Z0_t (SubBytesIns_Inst_Sbox_1_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M58), .B0_t (SubBytesIns_Inst_Sbox_1_L8), .Z0_t (SubBytesIns_Inst_Sbox_1_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_M63), .B0_t (SubBytesIns_Inst_Sbox_1_L4), .Z0_t (SubBytesIns_Inst_Sbox_1_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L0), .B0_t (SubBytesIns_Inst_Sbox_1_L1), .Z0_t (SubBytesIns_Inst_Sbox_1_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L1), .B0_t (SubBytesIns_Inst_Sbox_1_L7), .Z0_t (SubBytesIns_Inst_Sbox_1_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L3), .B0_t (SubBytesIns_Inst_Sbox_1_L12), .Z0_t (SubBytesIns_Inst_Sbox_1_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L18), .B0_t (SubBytesIns_Inst_Sbox_1_L2), .Z0_t (SubBytesIns_Inst_Sbox_1_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L15), .B0_t (SubBytesIns_Inst_Sbox_1_L9), .Z0_t (SubBytesIns_Inst_Sbox_1_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L6), .B0_t (SubBytesIns_Inst_Sbox_1_L10), .Z0_t (SubBytesIns_Inst_Sbox_1_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L7), .B0_t (SubBytesIns_Inst_Sbox_1_L9), .Z0_t (SubBytesIns_Inst_Sbox_1_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L8), .B0_t (SubBytesIns_Inst_Sbox_1_L10), .Z0_t (SubBytesIns_Inst_Sbox_1_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L11), .B0_t (SubBytesIns_Inst_Sbox_1_L14), .Z0_t (SubBytesIns_Inst_Sbox_1_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L11), .B0_t (SubBytesIns_Inst_Sbox_1_L17), .Z0_t (SubBytesIns_Inst_Sbox_1_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L6), .B0_t (SubBytesIns_Inst_Sbox_1_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L16), .B0_t (SubBytesIns_Inst_Sbox_1_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L19), .B0_t (SubBytesIns_Inst_Sbox_1_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L6), .B0_t (SubBytesIns_Inst_Sbox_1_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L20), .B0_t (SubBytesIns_Inst_Sbox_1_L22), .Z0_t (MixColumnsInput[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L25), .B0_t (SubBytesIns_Inst_Sbox_1_L29), .Z0_t (MixColumnsInput[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L13), .B0_t (SubBytesIns_Inst_Sbox_1_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_1_L6), .B0_t (SubBytesIns_Inst_Sbox_1_L23), .Z0_t (MixColumnsInput[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .A0_t (ciphertext[23]), .B0_t (ciphertext[20]), .Z0_t (SubBytesIns_Inst_Sbox_2_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .A0_t (ciphertext[23]), .B0_t (ciphertext[18]), .Z0_t (SubBytesIns_Inst_Sbox_2_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .A0_t (ciphertext[23]), .B0_t (ciphertext[17]), .Z0_t (SubBytesIns_Inst_Sbox_2_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .A0_t (ciphertext[20]), .B0_t (ciphertext[18]), .Z0_t (SubBytesIns_Inst_Sbox_2_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .A0_t (ciphertext[19]), .B0_t (ciphertext[17]), .Z0_t (SubBytesIns_Inst_Sbox_2_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T1), .B0_t (SubBytesIns_Inst_Sbox_2_T5), .Z0_t (SubBytesIns_Inst_Sbox_2_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .A0_t (ciphertext[22]), .B0_t (ciphertext[21]), .Z0_t (SubBytesIns_Inst_Sbox_2_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .A0_t (ciphertext[16]), .B0_t (SubBytesIns_Inst_Sbox_2_T6), .Z0_t (SubBytesIns_Inst_Sbox_2_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .A0_t (ciphertext[16]), .B0_t (SubBytesIns_Inst_Sbox_2_T7), .Z0_t (SubBytesIns_Inst_Sbox_2_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T6), .B0_t (SubBytesIns_Inst_Sbox_2_T7), .Z0_t (SubBytesIns_Inst_Sbox_2_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .A0_t (ciphertext[22]), .B0_t (ciphertext[18]), .Z0_t (SubBytesIns_Inst_Sbox_2_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .A0_t (ciphertext[21]), .B0_t (ciphertext[18]), .Z0_t (SubBytesIns_Inst_Sbox_2_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T3), .B0_t (SubBytesIns_Inst_Sbox_2_T4), .Z0_t (SubBytesIns_Inst_Sbox_2_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T6), .B0_t (SubBytesIns_Inst_Sbox_2_T11), .Z0_t (SubBytesIns_Inst_Sbox_2_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T5), .B0_t (SubBytesIns_Inst_Sbox_2_T11), .Z0_t (SubBytesIns_Inst_Sbox_2_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T5), .B0_t (SubBytesIns_Inst_Sbox_2_T12), .Z0_t (SubBytesIns_Inst_Sbox_2_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T9), .B0_t (SubBytesIns_Inst_Sbox_2_T16), .Z0_t (SubBytesIns_Inst_Sbox_2_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .A0_t (ciphertext[20]), .B0_t (ciphertext[16]), .Z0_t (SubBytesIns_Inst_Sbox_2_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T7), .B0_t (SubBytesIns_Inst_Sbox_2_T18), .Z0_t (SubBytesIns_Inst_Sbox_2_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T1), .B0_t (SubBytesIns_Inst_Sbox_2_T19), .Z0_t (SubBytesIns_Inst_Sbox_2_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .A0_t (ciphertext[17]), .B0_t (ciphertext[16]), .Z0_t (SubBytesIns_Inst_Sbox_2_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T7), .B0_t (SubBytesIns_Inst_Sbox_2_T21), .Z0_t (SubBytesIns_Inst_Sbox_2_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T2), .B0_t (SubBytesIns_Inst_Sbox_2_T22), .Z0_t (SubBytesIns_Inst_Sbox_2_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T2), .B0_t (SubBytesIns_Inst_Sbox_2_T10), .Z0_t (SubBytesIns_Inst_Sbox_2_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T20), .B0_t (SubBytesIns_Inst_Sbox_2_T17), .Z0_t (SubBytesIns_Inst_Sbox_2_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T3), .B0_t (SubBytesIns_Inst_Sbox_2_T16), .Z0_t (SubBytesIns_Inst_Sbox_2_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T1), .B0_t (SubBytesIns_Inst_Sbox_2_T12), .Z0_t (SubBytesIns_Inst_Sbox_2_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T13), .B0_t (SubBytesIns_Inst_Sbox_2_T6), .Z0_t (SubBytesIns_Inst_Sbox_2_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T23), .B0_t (SubBytesIns_Inst_Sbox_2_T8), .Z0_t (SubBytesIns_Inst_Sbox_2_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T14), .B0_t (SubBytesIns_Inst_Sbox_2_M1), .Z0_t (SubBytesIns_Inst_Sbox_2_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T19), .B0_t (ciphertext[16]), .Z0_t (SubBytesIns_Inst_Sbox_2_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M4), .B0_t (SubBytesIns_Inst_Sbox_2_M1), .Z0_t (SubBytesIns_Inst_Sbox_2_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T3), .B0_t (SubBytesIns_Inst_Sbox_2_T16), .Z0_t (SubBytesIns_Inst_Sbox_2_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T22), .B0_t (SubBytesIns_Inst_Sbox_2_T9), .Z0_t (SubBytesIns_Inst_Sbox_2_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T26), .B0_t (SubBytesIns_Inst_Sbox_2_M6), .Z0_t (SubBytesIns_Inst_Sbox_2_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T20), .B0_t (SubBytesIns_Inst_Sbox_2_T17), .Z0_t (SubBytesIns_Inst_Sbox_2_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M9), .B0_t (SubBytesIns_Inst_Sbox_2_M6), .Z0_t (SubBytesIns_Inst_Sbox_2_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T1), .B0_t (SubBytesIns_Inst_Sbox_2_T15), .Z0_t (SubBytesIns_Inst_Sbox_2_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T4), .B0_t (SubBytesIns_Inst_Sbox_2_T27), .Z0_t (SubBytesIns_Inst_Sbox_2_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M12), .B0_t (SubBytesIns_Inst_Sbox_2_M11), .Z0_t (SubBytesIns_Inst_Sbox_2_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_T2), .B0_t (SubBytesIns_Inst_Sbox_2_T10), .Z0_t (SubBytesIns_Inst_Sbox_2_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M14), .B0_t (SubBytesIns_Inst_Sbox_2_M11), .Z0_t (SubBytesIns_Inst_Sbox_2_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M3), .B0_t (SubBytesIns_Inst_Sbox_2_M2), .Z0_t (SubBytesIns_Inst_Sbox_2_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M5), .B0_t (SubBytesIns_Inst_Sbox_2_T24), .Z0_t (SubBytesIns_Inst_Sbox_2_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M8), .B0_t (SubBytesIns_Inst_Sbox_2_M7), .Z0_t (SubBytesIns_Inst_Sbox_2_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M10), .B0_t (SubBytesIns_Inst_Sbox_2_M15), .Z0_t (SubBytesIns_Inst_Sbox_2_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M16), .B0_t (SubBytesIns_Inst_Sbox_2_M13), .Z0_t (SubBytesIns_Inst_Sbox_2_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M17), .B0_t (SubBytesIns_Inst_Sbox_2_M15), .Z0_t (SubBytesIns_Inst_Sbox_2_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M18), .B0_t (SubBytesIns_Inst_Sbox_2_M13), .Z0_t (SubBytesIns_Inst_Sbox_2_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M19), .B0_t (SubBytesIns_Inst_Sbox_2_T25), .Z0_t (SubBytesIns_Inst_Sbox_2_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M22), .B0_t (SubBytesIns_Inst_Sbox_2_M23), .Z0_t (SubBytesIns_Inst_Sbox_2_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M22), .B0_t (SubBytesIns_Inst_Sbox_2_M20), .Z0_t (SubBytesIns_Inst_Sbox_2_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M21), .B0_t (SubBytesIns_Inst_Sbox_2_M25), .Z0_t (SubBytesIns_Inst_Sbox_2_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M20), .B0_t (SubBytesIns_Inst_Sbox_2_M21), .Z0_t (SubBytesIns_Inst_Sbox_2_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M23), .B0_t (SubBytesIns_Inst_Sbox_2_M25), .Z0_t (SubBytesIns_Inst_Sbox_2_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M28), .B0_t (SubBytesIns_Inst_Sbox_2_M27), .Z0_t (SubBytesIns_Inst_Sbox_2_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M26), .B0_t (SubBytesIns_Inst_Sbox_2_M24), .Z0_t (SubBytesIns_Inst_Sbox_2_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M20), .B0_t (SubBytesIns_Inst_Sbox_2_M23), .Z0_t (SubBytesIns_Inst_Sbox_2_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M27), .B0_t (SubBytesIns_Inst_Sbox_2_M31), .Z0_t (SubBytesIns_Inst_Sbox_2_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M27), .B0_t (SubBytesIns_Inst_Sbox_2_M25), .Z0_t (SubBytesIns_Inst_Sbox_2_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M21), .B0_t (SubBytesIns_Inst_Sbox_2_M22), .Z0_t (SubBytesIns_Inst_Sbox_2_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M24), .B0_t (SubBytesIns_Inst_Sbox_2_M34), .Z0_t (SubBytesIns_Inst_Sbox_2_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M24), .B0_t (SubBytesIns_Inst_Sbox_2_M25), .Z0_t (SubBytesIns_Inst_Sbox_2_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M21), .B0_t (SubBytesIns_Inst_Sbox_2_M29), .Z0_t (SubBytesIns_Inst_Sbox_2_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M32), .B0_t (SubBytesIns_Inst_Sbox_2_M33), .Z0_t (SubBytesIns_Inst_Sbox_2_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M23), .B0_t (SubBytesIns_Inst_Sbox_2_M30), .Z0_t (SubBytesIns_Inst_Sbox_2_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M35), .B0_t (SubBytesIns_Inst_Sbox_2_M36), .Z0_t (SubBytesIns_Inst_Sbox_2_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M38), .B0_t (SubBytesIns_Inst_Sbox_2_M40), .Z0_t (SubBytesIns_Inst_Sbox_2_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M37), .B0_t (SubBytesIns_Inst_Sbox_2_M39), .Z0_t (SubBytesIns_Inst_Sbox_2_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M37), .B0_t (SubBytesIns_Inst_Sbox_2_M38), .Z0_t (SubBytesIns_Inst_Sbox_2_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M39), .B0_t (SubBytesIns_Inst_Sbox_2_M40), .Z0_t (SubBytesIns_Inst_Sbox_2_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M42), .B0_t (SubBytesIns_Inst_Sbox_2_M41), .Z0_t (SubBytesIns_Inst_Sbox_2_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M44), .B0_t (SubBytesIns_Inst_Sbox_2_T6), .Z0_t (SubBytesIns_Inst_Sbox_2_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M40), .B0_t (SubBytesIns_Inst_Sbox_2_T8), .Z0_t (SubBytesIns_Inst_Sbox_2_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M39), .B0_t (ciphertext[16]), .Z0_t (SubBytesIns_Inst_Sbox_2_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M43), .B0_t (SubBytesIns_Inst_Sbox_2_T16), .Z0_t (SubBytesIns_Inst_Sbox_2_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M38), .B0_t (SubBytesIns_Inst_Sbox_2_T9), .Z0_t (SubBytesIns_Inst_Sbox_2_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M37), .B0_t (SubBytesIns_Inst_Sbox_2_T17), .Z0_t (SubBytesIns_Inst_Sbox_2_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M42), .B0_t (SubBytesIns_Inst_Sbox_2_T15), .Z0_t (SubBytesIns_Inst_Sbox_2_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M45), .B0_t (SubBytesIns_Inst_Sbox_2_T27), .Z0_t (SubBytesIns_Inst_Sbox_2_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M41), .B0_t (SubBytesIns_Inst_Sbox_2_T10), .Z0_t (SubBytesIns_Inst_Sbox_2_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M44), .B0_t (SubBytesIns_Inst_Sbox_2_T13), .Z0_t (SubBytesIns_Inst_Sbox_2_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M40), .B0_t (SubBytesIns_Inst_Sbox_2_T23), .Z0_t (SubBytesIns_Inst_Sbox_2_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M39), .B0_t (SubBytesIns_Inst_Sbox_2_T19), .Z0_t (SubBytesIns_Inst_Sbox_2_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M43), .B0_t (SubBytesIns_Inst_Sbox_2_T3), .Z0_t (SubBytesIns_Inst_Sbox_2_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M38), .B0_t (SubBytesIns_Inst_Sbox_2_T22), .Z0_t (SubBytesIns_Inst_Sbox_2_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M37), .B0_t (SubBytesIns_Inst_Sbox_2_T20), .Z0_t (SubBytesIns_Inst_Sbox_2_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M42), .B0_t (SubBytesIns_Inst_Sbox_2_T1), .Z0_t (SubBytesIns_Inst_Sbox_2_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M45), .B0_t (SubBytesIns_Inst_Sbox_2_T4), .Z0_t (SubBytesIns_Inst_Sbox_2_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M41), .B0_t (SubBytesIns_Inst_Sbox_2_T2), .Z0_t (SubBytesIns_Inst_Sbox_2_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M61), .B0_t (SubBytesIns_Inst_Sbox_2_M62), .Z0_t (SubBytesIns_Inst_Sbox_2_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M50), .B0_t (SubBytesIns_Inst_Sbox_2_M56), .Z0_t (SubBytesIns_Inst_Sbox_2_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M46), .B0_t (SubBytesIns_Inst_Sbox_2_M48), .Z0_t (SubBytesIns_Inst_Sbox_2_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M47), .B0_t (SubBytesIns_Inst_Sbox_2_M55), .Z0_t (SubBytesIns_Inst_Sbox_2_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M54), .B0_t (SubBytesIns_Inst_Sbox_2_M58), .Z0_t (SubBytesIns_Inst_Sbox_2_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M49), .B0_t (SubBytesIns_Inst_Sbox_2_M61), .Z0_t (SubBytesIns_Inst_Sbox_2_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M62), .B0_t (SubBytesIns_Inst_Sbox_2_L5), .Z0_t (SubBytesIns_Inst_Sbox_2_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M46), .B0_t (SubBytesIns_Inst_Sbox_2_L3), .Z0_t (SubBytesIns_Inst_Sbox_2_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M51), .B0_t (SubBytesIns_Inst_Sbox_2_M59), .Z0_t (SubBytesIns_Inst_Sbox_2_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M52), .B0_t (SubBytesIns_Inst_Sbox_2_M53), .Z0_t (SubBytesIns_Inst_Sbox_2_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M53), .B0_t (SubBytesIns_Inst_Sbox_2_L4), .Z0_t (SubBytesIns_Inst_Sbox_2_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M60), .B0_t (SubBytesIns_Inst_Sbox_2_L2), .Z0_t (SubBytesIns_Inst_Sbox_2_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M48), .B0_t (SubBytesIns_Inst_Sbox_2_M51), .Z0_t (SubBytesIns_Inst_Sbox_2_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M50), .B0_t (SubBytesIns_Inst_Sbox_2_L0), .Z0_t (SubBytesIns_Inst_Sbox_2_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M52), .B0_t (SubBytesIns_Inst_Sbox_2_M61), .Z0_t (SubBytesIns_Inst_Sbox_2_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M55), .B0_t (SubBytesIns_Inst_Sbox_2_L1), .Z0_t (SubBytesIns_Inst_Sbox_2_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M56), .B0_t (SubBytesIns_Inst_Sbox_2_L0), .Z0_t (SubBytesIns_Inst_Sbox_2_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M57), .B0_t (SubBytesIns_Inst_Sbox_2_L1), .Z0_t (SubBytesIns_Inst_Sbox_2_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M58), .B0_t (SubBytesIns_Inst_Sbox_2_L8), .Z0_t (SubBytesIns_Inst_Sbox_2_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_M63), .B0_t (SubBytesIns_Inst_Sbox_2_L4), .Z0_t (SubBytesIns_Inst_Sbox_2_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L0), .B0_t (SubBytesIns_Inst_Sbox_2_L1), .Z0_t (SubBytesIns_Inst_Sbox_2_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L1), .B0_t (SubBytesIns_Inst_Sbox_2_L7), .Z0_t (SubBytesIns_Inst_Sbox_2_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L3), .B0_t (SubBytesIns_Inst_Sbox_2_L12), .Z0_t (SubBytesIns_Inst_Sbox_2_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L18), .B0_t (SubBytesIns_Inst_Sbox_2_L2), .Z0_t (SubBytesIns_Inst_Sbox_2_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L15), .B0_t (SubBytesIns_Inst_Sbox_2_L9), .Z0_t (SubBytesIns_Inst_Sbox_2_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L6), .B0_t (SubBytesIns_Inst_Sbox_2_L10), .Z0_t (SubBytesIns_Inst_Sbox_2_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L7), .B0_t (SubBytesIns_Inst_Sbox_2_L9), .Z0_t (SubBytesIns_Inst_Sbox_2_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L8), .B0_t (SubBytesIns_Inst_Sbox_2_L10), .Z0_t (SubBytesIns_Inst_Sbox_2_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L11), .B0_t (SubBytesIns_Inst_Sbox_2_L14), .Z0_t (SubBytesIns_Inst_Sbox_2_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L11), .B0_t (SubBytesIns_Inst_Sbox_2_L17), .Z0_t (SubBytesIns_Inst_Sbox_2_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L6), .B0_t (SubBytesIns_Inst_Sbox_2_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L16), .B0_t (SubBytesIns_Inst_Sbox_2_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L19), .B0_t (SubBytesIns_Inst_Sbox_2_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L6), .B0_t (SubBytesIns_Inst_Sbox_2_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L20), .B0_t (SubBytesIns_Inst_Sbox_2_L22), .Z0_t (MixColumnsInput[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L25), .B0_t (SubBytesIns_Inst_Sbox_2_L29), .Z0_t (MixColumnsInput[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L13), .B0_t (SubBytesIns_Inst_Sbox_2_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_2_L6), .B0_t (SubBytesIns_Inst_Sbox_2_L23), .Z0_t (MixColumnsInput[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .A0_t (ciphertext[31]), .B0_t (ciphertext[28]), .Z0_t (SubBytesIns_Inst_Sbox_3_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .A0_t (ciphertext[31]), .B0_t (ciphertext[26]), .Z0_t (SubBytesIns_Inst_Sbox_3_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .A0_t (ciphertext[31]), .B0_t (ciphertext[25]), .Z0_t (SubBytesIns_Inst_Sbox_3_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .A0_t (ciphertext[28]), .B0_t (ciphertext[26]), .Z0_t (SubBytesIns_Inst_Sbox_3_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .A0_t (ciphertext[27]), .B0_t (ciphertext[25]), .Z0_t (SubBytesIns_Inst_Sbox_3_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T1), .B0_t (SubBytesIns_Inst_Sbox_3_T5), .Z0_t (SubBytesIns_Inst_Sbox_3_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .A0_t (ciphertext[30]), .B0_t (ciphertext[29]), .Z0_t (SubBytesIns_Inst_Sbox_3_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .A0_t (ciphertext[24]), .B0_t (SubBytesIns_Inst_Sbox_3_T6), .Z0_t (SubBytesIns_Inst_Sbox_3_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .A0_t (ciphertext[24]), .B0_t (SubBytesIns_Inst_Sbox_3_T7), .Z0_t (SubBytesIns_Inst_Sbox_3_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T6), .B0_t (SubBytesIns_Inst_Sbox_3_T7), .Z0_t (SubBytesIns_Inst_Sbox_3_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .A0_t (ciphertext[30]), .B0_t (ciphertext[26]), .Z0_t (SubBytesIns_Inst_Sbox_3_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .A0_t (ciphertext[29]), .B0_t (ciphertext[26]), .Z0_t (SubBytesIns_Inst_Sbox_3_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T3), .B0_t (SubBytesIns_Inst_Sbox_3_T4), .Z0_t (SubBytesIns_Inst_Sbox_3_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T6), .B0_t (SubBytesIns_Inst_Sbox_3_T11), .Z0_t (SubBytesIns_Inst_Sbox_3_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T5), .B0_t (SubBytesIns_Inst_Sbox_3_T11), .Z0_t (SubBytesIns_Inst_Sbox_3_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T5), .B0_t (SubBytesIns_Inst_Sbox_3_T12), .Z0_t (SubBytesIns_Inst_Sbox_3_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T9), .B0_t (SubBytesIns_Inst_Sbox_3_T16), .Z0_t (SubBytesIns_Inst_Sbox_3_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .A0_t (ciphertext[28]), .B0_t (ciphertext[24]), .Z0_t (SubBytesIns_Inst_Sbox_3_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T7), .B0_t (SubBytesIns_Inst_Sbox_3_T18), .Z0_t (SubBytesIns_Inst_Sbox_3_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T1), .B0_t (SubBytesIns_Inst_Sbox_3_T19), .Z0_t (SubBytesIns_Inst_Sbox_3_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .A0_t (ciphertext[25]), .B0_t (ciphertext[24]), .Z0_t (SubBytesIns_Inst_Sbox_3_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T7), .B0_t (SubBytesIns_Inst_Sbox_3_T21), .Z0_t (SubBytesIns_Inst_Sbox_3_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T2), .B0_t (SubBytesIns_Inst_Sbox_3_T22), .Z0_t (SubBytesIns_Inst_Sbox_3_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T2), .B0_t (SubBytesIns_Inst_Sbox_3_T10), .Z0_t (SubBytesIns_Inst_Sbox_3_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T20), .B0_t (SubBytesIns_Inst_Sbox_3_T17), .Z0_t (SubBytesIns_Inst_Sbox_3_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T3), .B0_t (SubBytesIns_Inst_Sbox_3_T16), .Z0_t (SubBytesIns_Inst_Sbox_3_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T1), .B0_t (SubBytesIns_Inst_Sbox_3_T12), .Z0_t (SubBytesIns_Inst_Sbox_3_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T13), .B0_t (SubBytesIns_Inst_Sbox_3_T6), .Z0_t (SubBytesIns_Inst_Sbox_3_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T23), .B0_t (SubBytesIns_Inst_Sbox_3_T8), .Z0_t (SubBytesIns_Inst_Sbox_3_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T14), .B0_t (SubBytesIns_Inst_Sbox_3_M1), .Z0_t (SubBytesIns_Inst_Sbox_3_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T19), .B0_t (ciphertext[24]), .Z0_t (SubBytesIns_Inst_Sbox_3_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M4), .B0_t (SubBytesIns_Inst_Sbox_3_M1), .Z0_t (SubBytesIns_Inst_Sbox_3_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T3), .B0_t (SubBytesIns_Inst_Sbox_3_T16), .Z0_t (SubBytesIns_Inst_Sbox_3_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T22), .B0_t (SubBytesIns_Inst_Sbox_3_T9), .Z0_t (SubBytesIns_Inst_Sbox_3_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T26), .B0_t (SubBytesIns_Inst_Sbox_3_M6), .Z0_t (SubBytesIns_Inst_Sbox_3_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T20), .B0_t (SubBytesIns_Inst_Sbox_3_T17), .Z0_t (SubBytesIns_Inst_Sbox_3_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M9), .B0_t (SubBytesIns_Inst_Sbox_3_M6), .Z0_t (SubBytesIns_Inst_Sbox_3_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T1), .B0_t (SubBytesIns_Inst_Sbox_3_T15), .Z0_t (SubBytesIns_Inst_Sbox_3_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T4), .B0_t (SubBytesIns_Inst_Sbox_3_T27), .Z0_t (SubBytesIns_Inst_Sbox_3_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M12), .B0_t (SubBytesIns_Inst_Sbox_3_M11), .Z0_t (SubBytesIns_Inst_Sbox_3_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_T2), .B0_t (SubBytesIns_Inst_Sbox_3_T10), .Z0_t (SubBytesIns_Inst_Sbox_3_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M14), .B0_t (SubBytesIns_Inst_Sbox_3_M11), .Z0_t (SubBytesIns_Inst_Sbox_3_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M3), .B0_t (SubBytesIns_Inst_Sbox_3_M2), .Z0_t (SubBytesIns_Inst_Sbox_3_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M5), .B0_t (SubBytesIns_Inst_Sbox_3_T24), .Z0_t (SubBytesIns_Inst_Sbox_3_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M8), .B0_t (SubBytesIns_Inst_Sbox_3_M7), .Z0_t (SubBytesIns_Inst_Sbox_3_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M10), .B0_t (SubBytesIns_Inst_Sbox_3_M15), .Z0_t (SubBytesIns_Inst_Sbox_3_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M16), .B0_t (SubBytesIns_Inst_Sbox_3_M13), .Z0_t (SubBytesIns_Inst_Sbox_3_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M17), .B0_t (SubBytesIns_Inst_Sbox_3_M15), .Z0_t (SubBytesIns_Inst_Sbox_3_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M18), .B0_t (SubBytesIns_Inst_Sbox_3_M13), .Z0_t (SubBytesIns_Inst_Sbox_3_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M19), .B0_t (SubBytesIns_Inst_Sbox_3_T25), .Z0_t (SubBytesIns_Inst_Sbox_3_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M22), .B0_t (SubBytesIns_Inst_Sbox_3_M23), .Z0_t (SubBytesIns_Inst_Sbox_3_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M22), .B0_t (SubBytesIns_Inst_Sbox_3_M20), .Z0_t (SubBytesIns_Inst_Sbox_3_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M21), .B0_t (SubBytesIns_Inst_Sbox_3_M25), .Z0_t (SubBytesIns_Inst_Sbox_3_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M20), .B0_t (SubBytesIns_Inst_Sbox_3_M21), .Z0_t (SubBytesIns_Inst_Sbox_3_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M23), .B0_t (SubBytesIns_Inst_Sbox_3_M25), .Z0_t (SubBytesIns_Inst_Sbox_3_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M28), .B0_t (SubBytesIns_Inst_Sbox_3_M27), .Z0_t (SubBytesIns_Inst_Sbox_3_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M26), .B0_t (SubBytesIns_Inst_Sbox_3_M24), .Z0_t (SubBytesIns_Inst_Sbox_3_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M20), .B0_t (SubBytesIns_Inst_Sbox_3_M23), .Z0_t (SubBytesIns_Inst_Sbox_3_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M27), .B0_t (SubBytesIns_Inst_Sbox_3_M31), .Z0_t (SubBytesIns_Inst_Sbox_3_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M27), .B0_t (SubBytesIns_Inst_Sbox_3_M25), .Z0_t (SubBytesIns_Inst_Sbox_3_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M21), .B0_t (SubBytesIns_Inst_Sbox_3_M22), .Z0_t (SubBytesIns_Inst_Sbox_3_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M24), .B0_t (SubBytesIns_Inst_Sbox_3_M34), .Z0_t (SubBytesIns_Inst_Sbox_3_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M24), .B0_t (SubBytesIns_Inst_Sbox_3_M25), .Z0_t (SubBytesIns_Inst_Sbox_3_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M21), .B0_t (SubBytesIns_Inst_Sbox_3_M29), .Z0_t (SubBytesIns_Inst_Sbox_3_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M32), .B0_t (SubBytesIns_Inst_Sbox_3_M33), .Z0_t (SubBytesIns_Inst_Sbox_3_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M23), .B0_t (SubBytesIns_Inst_Sbox_3_M30), .Z0_t (SubBytesIns_Inst_Sbox_3_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M35), .B0_t (SubBytesIns_Inst_Sbox_3_M36), .Z0_t (SubBytesIns_Inst_Sbox_3_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M38), .B0_t (SubBytesIns_Inst_Sbox_3_M40), .Z0_t (SubBytesIns_Inst_Sbox_3_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M37), .B0_t (SubBytesIns_Inst_Sbox_3_M39), .Z0_t (SubBytesIns_Inst_Sbox_3_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M37), .B0_t (SubBytesIns_Inst_Sbox_3_M38), .Z0_t (SubBytesIns_Inst_Sbox_3_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M39), .B0_t (SubBytesIns_Inst_Sbox_3_M40), .Z0_t (SubBytesIns_Inst_Sbox_3_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M42), .B0_t (SubBytesIns_Inst_Sbox_3_M41), .Z0_t (SubBytesIns_Inst_Sbox_3_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M44), .B0_t (SubBytesIns_Inst_Sbox_3_T6), .Z0_t (SubBytesIns_Inst_Sbox_3_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M40), .B0_t (SubBytesIns_Inst_Sbox_3_T8), .Z0_t (SubBytesIns_Inst_Sbox_3_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M39), .B0_t (ciphertext[24]), .Z0_t (SubBytesIns_Inst_Sbox_3_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M43), .B0_t (SubBytesIns_Inst_Sbox_3_T16), .Z0_t (SubBytesIns_Inst_Sbox_3_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M38), .B0_t (SubBytesIns_Inst_Sbox_3_T9), .Z0_t (SubBytesIns_Inst_Sbox_3_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M37), .B0_t (SubBytesIns_Inst_Sbox_3_T17), .Z0_t (SubBytesIns_Inst_Sbox_3_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M42), .B0_t (SubBytesIns_Inst_Sbox_3_T15), .Z0_t (SubBytesIns_Inst_Sbox_3_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M45), .B0_t (SubBytesIns_Inst_Sbox_3_T27), .Z0_t (SubBytesIns_Inst_Sbox_3_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M41), .B0_t (SubBytesIns_Inst_Sbox_3_T10), .Z0_t (SubBytesIns_Inst_Sbox_3_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M44), .B0_t (SubBytesIns_Inst_Sbox_3_T13), .Z0_t (SubBytesIns_Inst_Sbox_3_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M40), .B0_t (SubBytesIns_Inst_Sbox_3_T23), .Z0_t (SubBytesIns_Inst_Sbox_3_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M39), .B0_t (SubBytesIns_Inst_Sbox_3_T19), .Z0_t (SubBytesIns_Inst_Sbox_3_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M43), .B0_t (SubBytesIns_Inst_Sbox_3_T3), .Z0_t (SubBytesIns_Inst_Sbox_3_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M38), .B0_t (SubBytesIns_Inst_Sbox_3_T22), .Z0_t (SubBytesIns_Inst_Sbox_3_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M37), .B0_t (SubBytesIns_Inst_Sbox_3_T20), .Z0_t (SubBytesIns_Inst_Sbox_3_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M42), .B0_t (SubBytesIns_Inst_Sbox_3_T1), .Z0_t (SubBytesIns_Inst_Sbox_3_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M45), .B0_t (SubBytesIns_Inst_Sbox_3_T4), .Z0_t (SubBytesIns_Inst_Sbox_3_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M41), .B0_t (SubBytesIns_Inst_Sbox_3_T2), .Z0_t (SubBytesIns_Inst_Sbox_3_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M61), .B0_t (SubBytesIns_Inst_Sbox_3_M62), .Z0_t (SubBytesIns_Inst_Sbox_3_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M50), .B0_t (SubBytesIns_Inst_Sbox_3_M56), .Z0_t (SubBytesIns_Inst_Sbox_3_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M46), .B0_t (SubBytesIns_Inst_Sbox_3_M48), .Z0_t (SubBytesIns_Inst_Sbox_3_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M47), .B0_t (SubBytesIns_Inst_Sbox_3_M55), .Z0_t (SubBytesIns_Inst_Sbox_3_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M54), .B0_t (SubBytesIns_Inst_Sbox_3_M58), .Z0_t (SubBytesIns_Inst_Sbox_3_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M49), .B0_t (SubBytesIns_Inst_Sbox_3_M61), .Z0_t (SubBytesIns_Inst_Sbox_3_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M62), .B0_t (SubBytesIns_Inst_Sbox_3_L5), .Z0_t (SubBytesIns_Inst_Sbox_3_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M46), .B0_t (SubBytesIns_Inst_Sbox_3_L3), .Z0_t (SubBytesIns_Inst_Sbox_3_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M51), .B0_t (SubBytesIns_Inst_Sbox_3_M59), .Z0_t (SubBytesIns_Inst_Sbox_3_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M52), .B0_t (SubBytesIns_Inst_Sbox_3_M53), .Z0_t (SubBytesIns_Inst_Sbox_3_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M53), .B0_t (SubBytesIns_Inst_Sbox_3_L4), .Z0_t (SubBytesIns_Inst_Sbox_3_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M60), .B0_t (SubBytesIns_Inst_Sbox_3_L2), .Z0_t (SubBytesIns_Inst_Sbox_3_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M48), .B0_t (SubBytesIns_Inst_Sbox_3_M51), .Z0_t (SubBytesIns_Inst_Sbox_3_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M50), .B0_t (SubBytesIns_Inst_Sbox_3_L0), .Z0_t (SubBytesIns_Inst_Sbox_3_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M52), .B0_t (SubBytesIns_Inst_Sbox_3_M61), .Z0_t (SubBytesIns_Inst_Sbox_3_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M55), .B0_t (SubBytesIns_Inst_Sbox_3_L1), .Z0_t (SubBytesIns_Inst_Sbox_3_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M56), .B0_t (SubBytesIns_Inst_Sbox_3_L0), .Z0_t (SubBytesIns_Inst_Sbox_3_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M57), .B0_t (SubBytesIns_Inst_Sbox_3_L1), .Z0_t (SubBytesIns_Inst_Sbox_3_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M58), .B0_t (SubBytesIns_Inst_Sbox_3_L8), .Z0_t (SubBytesIns_Inst_Sbox_3_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_M63), .B0_t (SubBytesIns_Inst_Sbox_3_L4), .Z0_t (SubBytesIns_Inst_Sbox_3_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L0), .B0_t (SubBytesIns_Inst_Sbox_3_L1), .Z0_t (SubBytesIns_Inst_Sbox_3_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L1), .B0_t (SubBytesIns_Inst_Sbox_3_L7), .Z0_t (SubBytesIns_Inst_Sbox_3_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L3), .B0_t (SubBytesIns_Inst_Sbox_3_L12), .Z0_t (SubBytesIns_Inst_Sbox_3_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L18), .B0_t (SubBytesIns_Inst_Sbox_3_L2), .Z0_t (SubBytesIns_Inst_Sbox_3_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L15), .B0_t (SubBytesIns_Inst_Sbox_3_L9), .Z0_t (SubBytesIns_Inst_Sbox_3_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L6), .B0_t (SubBytesIns_Inst_Sbox_3_L10), .Z0_t (SubBytesIns_Inst_Sbox_3_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L7), .B0_t (SubBytesIns_Inst_Sbox_3_L9), .Z0_t (SubBytesIns_Inst_Sbox_3_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L8), .B0_t (SubBytesIns_Inst_Sbox_3_L10), .Z0_t (SubBytesIns_Inst_Sbox_3_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L11), .B0_t (SubBytesIns_Inst_Sbox_3_L14), .Z0_t (SubBytesIns_Inst_Sbox_3_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L11), .B0_t (SubBytesIns_Inst_Sbox_3_L17), .Z0_t (SubBytesIns_Inst_Sbox_3_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L6), .B0_t (SubBytesIns_Inst_Sbox_3_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L16), .B0_t (SubBytesIns_Inst_Sbox_3_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L19), .B0_t (SubBytesIns_Inst_Sbox_3_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L6), .B0_t (SubBytesIns_Inst_Sbox_3_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L20), .B0_t (SubBytesIns_Inst_Sbox_3_L22), .Z0_t (MixColumnsInput[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L25), .B0_t (SubBytesIns_Inst_Sbox_3_L29), .Z0_t (MixColumnsInput[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L13), .B0_t (SubBytesIns_Inst_Sbox_3_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_3_L6), .B0_t (SubBytesIns_Inst_Sbox_3_L23), .Z0_t (MixColumnsInput[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T1_U1 ( .A0_t (ciphertext[39]), .B0_t (ciphertext[36]), .Z0_t (SubBytesIns_Inst_Sbox_4_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T2_U1 ( .A0_t (ciphertext[39]), .B0_t (ciphertext[34]), .Z0_t (SubBytesIns_Inst_Sbox_4_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T3_U1 ( .A0_t (ciphertext[39]), .B0_t (ciphertext[33]), .Z0_t (SubBytesIns_Inst_Sbox_4_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T4_U1 ( .A0_t (ciphertext[36]), .B0_t (ciphertext[34]), .Z0_t (SubBytesIns_Inst_Sbox_4_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T5_U1 ( .A0_t (ciphertext[35]), .B0_t (ciphertext[33]), .Z0_t (SubBytesIns_Inst_Sbox_4_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T1), .B0_t (SubBytesIns_Inst_Sbox_4_T5), .Z0_t (SubBytesIns_Inst_Sbox_4_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T7_U1 ( .A0_t (ciphertext[38]), .B0_t (ciphertext[37]), .Z0_t (SubBytesIns_Inst_Sbox_4_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T8_U1 ( .A0_t (ciphertext[32]), .B0_t (SubBytesIns_Inst_Sbox_4_T6), .Z0_t (SubBytesIns_Inst_Sbox_4_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T9_U1 ( .A0_t (ciphertext[32]), .B0_t (SubBytesIns_Inst_Sbox_4_T7), .Z0_t (SubBytesIns_Inst_Sbox_4_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T6), .B0_t (SubBytesIns_Inst_Sbox_4_T7), .Z0_t (SubBytesIns_Inst_Sbox_4_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T11_U1 ( .A0_t (ciphertext[38]), .B0_t (ciphertext[34]), .Z0_t (SubBytesIns_Inst_Sbox_4_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T12_U1 ( .A0_t (ciphertext[37]), .B0_t (ciphertext[34]), .Z0_t (SubBytesIns_Inst_Sbox_4_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T3), .B0_t (SubBytesIns_Inst_Sbox_4_T4), .Z0_t (SubBytesIns_Inst_Sbox_4_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T6), .B0_t (SubBytesIns_Inst_Sbox_4_T11), .Z0_t (SubBytesIns_Inst_Sbox_4_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T5), .B0_t (SubBytesIns_Inst_Sbox_4_T11), .Z0_t (SubBytesIns_Inst_Sbox_4_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T5), .B0_t (SubBytesIns_Inst_Sbox_4_T12), .Z0_t (SubBytesIns_Inst_Sbox_4_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T9), .B0_t (SubBytesIns_Inst_Sbox_4_T16), .Z0_t (SubBytesIns_Inst_Sbox_4_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T18_U1 ( .A0_t (ciphertext[36]), .B0_t (ciphertext[32]), .Z0_t (SubBytesIns_Inst_Sbox_4_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T7), .B0_t (SubBytesIns_Inst_Sbox_4_T18), .Z0_t (SubBytesIns_Inst_Sbox_4_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T1), .B0_t (SubBytesIns_Inst_Sbox_4_T19), .Z0_t (SubBytesIns_Inst_Sbox_4_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T21_U1 ( .A0_t (ciphertext[33]), .B0_t (ciphertext[32]), .Z0_t (SubBytesIns_Inst_Sbox_4_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T7), .B0_t (SubBytesIns_Inst_Sbox_4_T21), .Z0_t (SubBytesIns_Inst_Sbox_4_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T2), .B0_t (SubBytesIns_Inst_Sbox_4_T22), .Z0_t (SubBytesIns_Inst_Sbox_4_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T2), .B0_t (SubBytesIns_Inst_Sbox_4_T10), .Z0_t (SubBytesIns_Inst_Sbox_4_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T20), .B0_t (SubBytesIns_Inst_Sbox_4_T17), .Z0_t (SubBytesIns_Inst_Sbox_4_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T3), .B0_t (SubBytesIns_Inst_Sbox_4_T16), .Z0_t (SubBytesIns_Inst_Sbox_4_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T1), .B0_t (SubBytesIns_Inst_Sbox_4_T12), .Z0_t (SubBytesIns_Inst_Sbox_4_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T13), .B0_t (SubBytesIns_Inst_Sbox_4_T6), .Z0_t (SubBytesIns_Inst_Sbox_4_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T23), .B0_t (SubBytesIns_Inst_Sbox_4_T8), .Z0_t (SubBytesIns_Inst_Sbox_4_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T14), .B0_t (SubBytesIns_Inst_Sbox_4_M1), .Z0_t (SubBytesIns_Inst_Sbox_4_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T19), .B0_t (ciphertext[32]), .Z0_t (SubBytesIns_Inst_Sbox_4_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M4), .B0_t (SubBytesIns_Inst_Sbox_4_M1), .Z0_t (SubBytesIns_Inst_Sbox_4_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T3), .B0_t (SubBytesIns_Inst_Sbox_4_T16), .Z0_t (SubBytesIns_Inst_Sbox_4_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T22), .B0_t (SubBytesIns_Inst_Sbox_4_T9), .Z0_t (SubBytesIns_Inst_Sbox_4_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T26), .B0_t (SubBytesIns_Inst_Sbox_4_M6), .Z0_t (SubBytesIns_Inst_Sbox_4_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T20), .B0_t (SubBytesIns_Inst_Sbox_4_T17), .Z0_t (SubBytesIns_Inst_Sbox_4_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M9), .B0_t (SubBytesIns_Inst_Sbox_4_M6), .Z0_t (SubBytesIns_Inst_Sbox_4_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T1), .B0_t (SubBytesIns_Inst_Sbox_4_T15), .Z0_t (SubBytesIns_Inst_Sbox_4_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T4), .B0_t (SubBytesIns_Inst_Sbox_4_T27), .Z0_t (SubBytesIns_Inst_Sbox_4_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M12), .B0_t (SubBytesIns_Inst_Sbox_4_M11), .Z0_t (SubBytesIns_Inst_Sbox_4_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_T2), .B0_t (SubBytesIns_Inst_Sbox_4_T10), .Z0_t (SubBytesIns_Inst_Sbox_4_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M14), .B0_t (SubBytesIns_Inst_Sbox_4_M11), .Z0_t (SubBytesIns_Inst_Sbox_4_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M3), .B0_t (SubBytesIns_Inst_Sbox_4_M2), .Z0_t (SubBytesIns_Inst_Sbox_4_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M5), .B0_t (SubBytesIns_Inst_Sbox_4_T24), .Z0_t (SubBytesIns_Inst_Sbox_4_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M8), .B0_t (SubBytesIns_Inst_Sbox_4_M7), .Z0_t (SubBytesIns_Inst_Sbox_4_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M10), .B0_t (SubBytesIns_Inst_Sbox_4_M15), .Z0_t (SubBytesIns_Inst_Sbox_4_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M16), .B0_t (SubBytesIns_Inst_Sbox_4_M13), .Z0_t (SubBytesIns_Inst_Sbox_4_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M17), .B0_t (SubBytesIns_Inst_Sbox_4_M15), .Z0_t (SubBytesIns_Inst_Sbox_4_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M18), .B0_t (SubBytesIns_Inst_Sbox_4_M13), .Z0_t (SubBytesIns_Inst_Sbox_4_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M19), .B0_t (SubBytesIns_Inst_Sbox_4_T25), .Z0_t (SubBytesIns_Inst_Sbox_4_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M22), .B0_t (SubBytesIns_Inst_Sbox_4_M23), .Z0_t (SubBytesIns_Inst_Sbox_4_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M22), .B0_t (SubBytesIns_Inst_Sbox_4_M20), .Z0_t (SubBytesIns_Inst_Sbox_4_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M21), .B0_t (SubBytesIns_Inst_Sbox_4_M25), .Z0_t (SubBytesIns_Inst_Sbox_4_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M20), .B0_t (SubBytesIns_Inst_Sbox_4_M21), .Z0_t (SubBytesIns_Inst_Sbox_4_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M23), .B0_t (SubBytesIns_Inst_Sbox_4_M25), .Z0_t (SubBytesIns_Inst_Sbox_4_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M28), .B0_t (SubBytesIns_Inst_Sbox_4_M27), .Z0_t (SubBytesIns_Inst_Sbox_4_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M26), .B0_t (SubBytesIns_Inst_Sbox_4_M24), .Z0_t (SubBytesIns_Inst_Sbox_4_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M20), .B0_t (SubBytesIns_Inst_Sbox_4_M23), .Z0_t (SubBytesIns_Inst_Sbox_4_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M27), .B0_t (SubBytesIns_Inst_Sbox_4_M31), .Z0_t (SubBytesIns_Inst_Sbox_4_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M27), .B0_t (SubBytesIns_Inst_Sbox_4_M25), .Z0_t (SubBytesIns_Inst_Sbox_4_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M21), .B0_t (SubBytesIns_Inst_Sbox_4_M22), .Z0_t (SubBytesIns_Inst_Sbox_4_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M24), .B0_t (SubBytesIns_Inst_Sbox_4_M34), .Z0_t (SubBytesIns_Inst_Sbox_4_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M24), .B0_t (SubBytesIns_Inst_Sbox_4_M25), .Z0_t (SubBytesIns_Inst_Sbox_4_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M21), .B0_t (SubBytesIns_Inst_Sbox_4_M29), .Z0_t (SubBytesIns_Inst_Sbox_4_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M32), .B0_t (SubBytesIns_Inst_Sbox_4_M33), .Z0_t (SubBytesIns_Inst_Sbox_4_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M23), .B0_t (SubBytesIns_Inst_Sbox_4_M30), .Z0_t (SubBytesIns_Inst_Sbox_4_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M35), .B0_t (SubBytesIns_Inst_Sbox_4_M36), .Z0_t (SubBytesIns_Inst_Sbox_4_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M38), .B0_t (SubBytesIns_Inst_Sbox_4_M40), .Z0_t (SubBytesIns_Inst_Sbox_4_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M37), .B0_t (SubBytesIns_Inst_Sbox_4_M39), .Z0_t (SubBytesIns_Inst_Sbox_4_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M37), .B0_t (SubBytesIns_Inst_Sbox_4_M38), .Z0_t (SubBytesIns_Inst_Sbox_4_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M39), .B0_t (SubBytesIns_Inst_Sbox_4_M40), .Z0_t (SubBytesIns_Inst_Sbox_4_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M42), .B0_t (SubBytesIns_Inst_Sbox_4_M41), .Z0_t (SubBytesIns_Inst_Sbox_4_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M44), .B0_t (SubBytesIns_Inst_Sbox_4_T6), .Z0_t (SubBytesIns_Inst_Sbox_4_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M40), .B0_t (SubBytesIns_Inst_Sbox_4_T8), .Z0_t (SubBytesIns_Inst_Sbox_4_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M39), .B0_t (ciphertext[32]), .Z0_t (SubBytesIns_Inst_Sbox_4_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M43), .B0_t (SubBytesIns_Inst_Sbox_4_T16), .Z0_t (SubBytesIns_Inst_Sbox_4_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M38), .B0_t (SubBytesIns_Inst_Sbox_4_T9), .Z0_t (SubBytesIns_Inst_Sbox_4_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M37), .B0_t (SubBytesIns_Inst_Sbox_4_T17), .Z0_t (SubBytesIns_Inst_Sbox_4_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M42), .B0_t (SubBytesIns_Inst_Sbox_4_T15), .Z0_t (SubBytesIns_Inst_Sbox_4_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M45), .B0_t (SubBytesIns_Inst_Sbox_4_T27), .Z0_t (SubBytesIns_Inst_Sbox_4_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M41), .B0_t (SubBytesIns_Inst_Sbox_4_T10), .Z0_t (SubBytesIns_Inst_Sbox_4_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M44), .B0_t (SubBytesIns_Inst_Sbox_4_T13), .Z0_t (SubBytesIns_Inst_Sbox_4_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M40), .B0_t (SubBytesIns_Inst_Sbox_4_T23), .Z0_t (SubBytesIns_Inst_Sbox_4_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M39), .B0_t (SubBytesIns_Inst_Sbox_4_T19), .Z0_t (SubBytesIns_Inst_Sbox_4_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M43), .B0_t (SubBytesIns_Inst_Sbox_4_T3), .Z0_t (SubBytesIns_Inst_Sbox_4_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M38), .B0_t (SubBytesIns_Inst_Sbox_4_T22), .Z0_t (SubBytesIns_Inst_Sbox_4_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M37), .B0_t (SubBytesIns_Inst_Sbox_4_T20), .Z0_t (SubBytesIns_Inst_Sbox_4_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M42), .B0_t (SubBytesIns_Inst_Sbox_4_T1), .Z0_t (SubBytesIns_Inst_Sbox_4_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M45), .B0_t (SubBytesIns_Inst_Sbox_4_T4), .Z0_t (SubBytesIns_Inst_Sbox_4_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M41), .B0_t (SubBytesIns_Inst_Sbox_4_T2), .Z0_t (SubBytesIns_Inst_Sbox_4_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M61), .B0_t (SubBytesIns_Inst_Sbox_4_M62), .Z0_t (SubBytesIns_Inst_Sbox_4_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M50), .B0_t (SubBytesIns_Inst_Sbox_4_M56), .Z0_t (SubBytesIns_Inst_Sbox_4_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M46), .B0_t (SubBytesIns_Inst_Sbox_4_M48), .Z0_t (SubBytesIns_Inst_Sbox_4_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M47), .B0_t (SubBytesIns_Inst_Sbox_4_M55), .Z0_t (SubBytesIns_Inst_Sbox_4_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M54), .B0_t (SubBytesIns_Inst_Sbox_4_M58), .Z0_t (SubBytesIns_Inst_Sbox_4_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M49), .B0_t (SubBytesIns_Inst_Sbox_4_M61), .Z0_t (SubBytesIns_Inst_Sbox_4_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M62), .B0_t (SubBytesIns_Inst_Sbox_4_L5), .Z0_t (SubBytesIns_Inst_Sbox_4_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M46), .B0_t (SubBytesIns_Inst_Sbox_4_L3), .Z0_t (SubBytesIns_Inst_Sbox_4_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M51), .B0_t (SubBytesIns_Inst_Sbox_4_M59), .Z0_t (SubBytesIns_Inst_Sbox_4_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M52), .B0_t (SubBytesIns_Inst_Sbox_4_M53), .Z0_t (SubBytesIns_Inst_Sbox_4_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M53), .B0_t (SubBytesIns_Inst_Sbox_4_L4), .Z0_t (SubBytesIns_Inst_Sbox_4_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M60), .B0_t (SubBytesIns_Inst_Sbox_4_L2), .Z0_t (SubBytesIns_Inst_Sbox_4_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M48), .B0_t (SubBytesIns_Inst_Sbox_4_M51), .Z0_t (SubBytesIns_Inst_Sbox_4_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M50), .B0_t (SubBytesIns_Inst_Sbox_4_L0), .Z0_t (SubBytesIns_Inst_Sbox_4_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M52), .B0_t (SubBytesIns_Inst_Sbox_4_M61), .Z0_t (SubBytesIns_Inst_Sbox_4_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M55), .B0_t (SubBytesIns_Inst_Sbox_4_L1), .Z0_t (SubBytesIns_Inst_Sbox_4_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M56), .B0_t (SubBytesIns_Inst_Sbox_4_L0), .Z0_t (SubBytesIns_Inst_Sbox_4_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M57), .B0_t (SubBytesIns_Inst_Sbox_4_L1), .Z0_t (SubBytesIns_Inst_Sbox_4_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M58), .B0_t (SubBytesIns_Inst_Sbox_4_L8), .Z0_t (SubBytesIns_Inst_Sbox_4_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_M63), .B0_t (SubBytesIns_Inst_Sbox_4_L4), .Z0_t (SubBytesIns_Inst_Sbox_4_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L0), .B0_t (SubBytesIns_Inst_Sbox_4_L1), .Z0_t (SubBytesIns_Inst_Sbox_4_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L1), .B0_t (SubBytesIns_Inst_Sbox_4_L7), .Z0_t (SubBytesIns_Inst_Sbox_4_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L3), .B0_t (SubBytesIns_Inst_Sbox_4_L12), .Z0_t (SubBytesIns_Inst_Sbox_4_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L18), .B0_t (SubBytesIns_Inst_Sbox_4_L2), .Z0_t (SubBytesIns_Inst_Sbox_4_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L15), .B0_t (SubBytesIns_Inst_Sbox_4_L9), .Z0_t (SubBytesIns_Inst_Sbox_4_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L6), .B0_t (SubBytesIns_Inst_Sbox_4_L10), .Z0_t (SubBytesIns_Inst_Sbox_4_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L7), .B0_t (SubBytesIns_Inst_Sbox_4_L9), .Z0_t (SubBytesIns_Inst_Sbox_4_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L8), .B0_t (SubBytesIns_Inst_Sbox_4_L10), .Z0_t (SubBytesIns_Inst_Sbox_4_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L11), .B0_t (SubBytesIns_Inst_Sbox_4_L14), .Z0_t (SubBytesIns_Inst_Sbox_4_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L11), .B0_t (SubBytesIns_Inst_Sbox_4_L17), .Z0_t (SubBytesIns_Inst_Sbox_4_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L6), .B0_t (SubBytesIns_Inst_Sbox_4_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L16), .B0_t (SubBytesIns_Inst_Sbox_4_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L19), .B0_t (SubBytesIns_Inst_Sbox_4_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L6), .B0_t (SubBytesIns_Inst_Sbox_4_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L20), .B0_t (SubBytesIns_Inst_Sbox_4_L22), .Z0_t (MixColumnsInput[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L25), .B0_t (SubBytesIns_Inst_Sbox_4_L29), .Z0_t (MixColumnsInput[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L13), .B0_t (SubBytesIns_Inst_Sbox_4_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_4_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_4_L6), .B0_t (SubBytesIns_Inst_Sbox_4_L23), .Z0_t (MixColumnsInput[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T1_U1 ( .A0_t (ciphertext[47]), .B0_t (ciphertext[44]), .Z0_t (SubBytesIns_Inst_Sbox_5_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T2_U1 ( .A0_t (ciphertext[47]), .B0_t (ciphertext[42]), .Z0_t (SubBytesIns_Inst_Sbox_5_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T3_U1 ( .A0_t (ciphertext[47]), .B0_t (ciphertext[41]), .Z0_t (SubBytesIns_Inst_Sbox_5_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T4_U1 ( .A0_t (ciphertext[44]), .B0_t (ciphertext[42]), .Z0_t (SubBytesIns_Inst_Sbox_5_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T5_U1 ( .A0_t (ciphertext[43]), .B0_t (ciphertext[41]), .Z0_t (SubBytesIns_Inst_Sbox_5_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T1), .B0_t (SubBytesIns_Inst_Sbox_5_T5), .Z0_t (SubBytesIns_Inst_Sbox_5_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T7_U1 ( .A0_t (ciphertext[46]), .B0_t (ciphertext[45]), .Z0_t (SubBytesIns_Inst_Sbox_5_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T8_U1 ( .A0_t (ciphertext[40]), .B0_t (SubBytesIns_Inst_Sbox_5_T6), .Z0_t (SubBytesIns_Inst_Sbox_5_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T9_U1 ( .A0_t (ciphertext[40]), .B0_t (SubBytesIns_Inst_Sbox_5_T7), .Z0_t (SubBytesIns_Inst_Sbox_5_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T6), .B0_t (SubBytesIns_Inst_Sbox_5_T7), .Z0_t (SubBytesIns_Inst_Sbox_5_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T11_U1 ( .A0_t (ciphertext[46]), .B0_t (ciphertext[42]), .Z0_t (SubBytesIns_Inst_Sbox_5_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T12_U1 ( .A0_t (ciphertext[45]), .B0_t (ciphertext[42]), .Z0_t (SubBytesIns_Inst_Sbox_5_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T3), .B0_t (SubBytesIns_Inst_Sbox_5_T4), .Z0_t (SubBytesIns_Inst_Sbox_5_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T6), .B0_t (SubBytesIns_Inst_Sbox_5_T11), .Z0_t (SubBytesIns_Inst_Sbox_5_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T5), .B0_t (SubBytesIns_Inst_Sbox_5_T11), .Z0_t (SubBytesIns_Inst_Sbox_5_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T5), .B0_t (SubBytesIns_Inst_Sbox_5_T12), .Z0_t (SubBytesIns_Inst_Sbox_5_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T9), .B0_t (SubBytesIns_Inst_Sbox_5_T16), .Z0_t (SubBytesIns_Inst_Sbox_5_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T18_U1 ( .A0_t (ciphertext[44]), .B0_t (ciphertext[40]), .Z0_t (SubBytesIns_Inst_Sbox_5_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T7), .B0_t (SubBytesIns_Inst_Sbox_5_T18), .Z0_t (SubBytesIns_Inst_Sbox_5_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T1), .B0_t (SubBytesIns_Inst_Sbox_5_T19), .Z0_t (SubBytesIns_Inst_Sbox_5_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T21_U1 ( .A0_t (ciphertext[41]), .B0_t (ciphertext[40]), .Z0_t (SubBytesIns_Inst_Sbox_5_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T7), .B0_t (SubBytesIns_Inst_Sbox_5_T21), .Z0_t (SubBytesIns_Inst_Sbox_5_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T2), .B0_t (SubBytesIns_Inst_Sbox_5_T22), .Z0_t (SubBytesIns_Inst_Sbox_5_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T2), .B0_t (SubBytesIns_Inst_Sbox_5_T10), .Z0_t (SubBytesIns_Inst_Sbox_5_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T20), .B0_t (SubBytesIns_Inst_Sbox_5_T17), .Z0_t (SubBytesIns_Inst_Sbox_5_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T3), .B0_t (SubBytesIns_Inst_Sbox_5_T16), .Z0_t (SubBytesIns_Inst_Sbox_5_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T1), .B0_t (SubBytesIns_Inst_Sbox_5_T12), .Z0_t (SubBytesIns_Inst_Sbox_5_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T13), .B0_t (SubBytesIns_Inst_Sbox_5_T6), .Z0_t (SubBytesIns_Inst_Sbox_5_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T23), .B0_t (SubBytesIns_Inst_Sbox_5_T8), .Z0_t (SubBytesIns_Inst_Sbox_5_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T14), .B0_t (SubBytesIns_Inst_Sbox_5_M1), .Z0_t (SubBytesIns_Inst_Sbox_5_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T19), .B0_t (ciphertext[40]), .Z0_t (SubBytesIns_Inst_Sbox_5_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M4), .B0_t (SubBytesIns_Inst_Sbox_5_M1), .Z0_t (SubBytesIns_Inst_Sbox_5_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T3), .B0_t (SubBytesIns_Inst_Sbox_5_T16), .Z0_t (SubBytesIns_Inst_Sbox_5_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T22), .B0_t (SubBytesIns_Inst_Sbox_5_T9), .Z0_t (SubBytesIns_Inst_Sbox_5_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T26), .B0_t (SubBytesIns_Inst_Sbox_5_M6), .Z0_t (SubBytesIns_Inst_Sbox_5_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T20), .B0_t (SubBytesIns_Inst_Sbox_5_T17), .Z0_t (SubBytesIns_Inst_Sbox_5_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M9), .B0_t (SubBytesIns_Inst_Sbox_5_M6), .Z0_t (SubBytesIns_Inst_Sbox_5_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T1), .B0_t (SubBytesIns_Inst_Sbox_5_T15), .Z0_t (SubBytesIns_Inst_Sbox_5_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T4), .B0_t (SubBytesIns_Inst_Sbox_5_T27), .Z0_t (SubBytesIns_Inst_Sbox_5_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M12), .B0_t (SubBytesIns_Inst_Sbox_5_M11), .Z0_t (SubBytesIns_Inst_Sbox_5_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_T2), .B0_t (SubBytesIns_Inst_Sbox_5_T10), .Z0_t (SubBytesIns_Inst_Sbox_5_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M14), .B0_t (SubBytesIns_Inst_Sbox_5_M11), .Z0_t (SubBytesIns_Inst_Sbox_5_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M3), .B0_t (SubBytesIns_Inst_Sbox_5_M2), .Z0_t (SubBytesIns_Inst_Sbox_5_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M5), .B0_t (SubBytesIns_Inst_Sbox_5_T24), .Z0_t (SubBytesIns_Inst_Sbox_5_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M8), .B0_t (SubBytesIns_Inst_Sbox_5_M7), .Z0_t (SubBytesIns_Inst_Sbox_5_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M10), .B0_t (SubBytesIns_Inst_Sbox_5_M15), .Z0_t (SubBytesIns_Inst_Sbox_5_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M16), .B0_t (SubBytesIns_Inst_Sbox_5_M13), .Z0_t (SubBytesIns_Inst_Sbox_5_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M17), .B0_t (SubBytesIns_Inst_Sbox_5_M15), .Z0_t (SubBytesIns_Inst_Sbox_5_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M18), .B0_t (SubBytesIns_Inst_Sbox_5_M13), .Z0_t (SubBytesIns_Inst_Sbox_5_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M19), .B0_t (SubBytesIns_Inst_Sbox_5_T25), .Z0_t (SubBytesIns_Inst_Sbox_5_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M22), .B0_t (SubBytesIns_Inst_Sbox_5_M23), .Z0_t (SubBytesIns_Inst_Sbox_5_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M22), .B0_t (SubBytesIns_Inst_Sbox_5_M20), .Z0_t (SubBytesIns_Inst_Sbox_5_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M21), .B0_t (SubBytesIns_Inst_Sbox_5_M25), .Z0_t (SubBytesIns_Inst_Sbox_5_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M20), .B0_t (SubBytesIns_Inst_Sbox_5_M21), .Z0_t (SubBytesIns_Inst_Sbox_5_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M23), .B0_t (SubBytesIns_Inst_Sbox_5_M25), .Z0_t (SubBytesIns_Inst_Sbox_5_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M28), .B0_t (SubBytesIns_Inst_Sbox_5_M27), .Z0_t (SubBytesIns_Inst_Sbox_5_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M26), .B0_t (SubBytesIns_Inst_Sbox_5_M24), .Z0_t (SubBytesIns_Inst_Sbox_5_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M20), .B0_t (SubBytesIns_Inst_Sbox_5_M23), .Z0_t (SubBytesIns_Inst_Sbox_5_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M27), .B0_t (SubBytesIns_Inst_Sbox_5_M31), .Z0_t (SubBytesIns_Inst_Sbox_5_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M27), .B0_t (SubBytesIns_Inst_Sbox_5_M25), .Z0_t (SubBytesIns_Inst_Sbox_5_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M21), .B0_t (SubBytesIns_Inst_Sbox_5_M22), .Z0_t (SubBytesIns_Inst_Sbox_5_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M24), .B0_t (SubBytesIns_Inst_Sbox_5_M34), .Z0_t (SubBytesIns_Inst_Sbox_5_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M24), .B0_t (SubBytesIns_Inst_Sbox_5_M25), .Z0_t (SubBytesIns_Inst_Sbox_5_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M21), .B0_t (SubBytesIns_Inst_Sbox_5_M29), .Z0_t (SubBytesIns_Inst_Sbox_5_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M32), .B0_t (SubBytesIns_Inst_Sbox_5_M33), .Z0_t (SubBytesIns_Inst_Sbox_5_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M23), .B0_t (SubBytesIns_Inst_Sbox_5_M30), .Z0_t (SubBytesIns_Inst_Sbox_5_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M35), .B0_t (SubBytesIns_Inst_Sbox_5_M36), .Z0_t (SubBytesIns_Inst_Sbox_5_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M38), .B0_t (SubBytesIns_Inst_Sbox_5_M40), .Z0_t (SubBytesIns_Inst_Sbox_5_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M37), .B0_t (SubBytesIns_Inst_Sbox_5_M39), .Z0_t (SubBytesIns_Inst_Sbox_5_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M37), .B0_t (SubBytesIns_Inst_Sbox_5_M38), .Z0_t (SubBytesIns_Inst_Sbox_5_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M39), .B0_t (SubBytesIns_Inst_Sbox_5_M40), .Z0_t (SubBytesIns_Inst_Sbox_5_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M42), .B0_t (SubBytesIns_Inst_Sbox_5_M41), .Z0_t (SubBytesIns_Inst_Sbox_5_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M44), .B0_t (SubBytesIns_Inst_Sbox_5_T6), .Z0_t (SubBytesIns_Inst_Sbox_5_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M40), .B0_t (SubBytesIns_Inst_Sbox_5_T8), .Z0_t (SubBytesIns_Inst_Sbox_5_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M39), .B0_t (ciphertext[40]), .Z0_t (SubBytesIns_Inst_Sbox_5_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M43), .B0_t (SubBytesIns_Inst_Sbox_5_T16), .Z0_t (SubBytesIns_Inst_Sbox_5_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M38), .B0_t (SubBytesIns_Inst_Sbox_5_T9), .Z0_t (SubBytesIns_Inst_Sbox_5_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M37), .B0_t (SubBytesIns_Inst_Sbox_5_T17), .Z0_t (SubBytesIns_Inst_Sbox_5_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M42), .B0_t (SubBytesIns_Inst_Sbox_5_T15), .Z0_t (SubBytesIns_Inst_Sbox_5_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M45), .B0_t (SubBytesIns_Inst_Sbox_5_T27), .Z0_t (SubBytesIns_Inst_Sbox_5_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M41), .B0_t (SubBytesIns_Inst_Sbox_5_T10), .Z0_t (SubBytesIns_Inst_Sbox_5_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M44), .B0_t (SubBytesIns_Inst_Sbox_5_T13), .Z0_t (SubBytesIns_Inst_Sbox_5_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M40), .B0_t (SubBytesIns_Inst_Sbox_5_T23), .Z0_t (SubBytesIns_Inst_Sbox_5_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M39), .B0_t (SubBytesIns_Inst_Sbox_5_T19), .Z0_t (SubBytesIns_Inst_Sbox_5_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M43), .B0_t (SubBytesIns_Inst_Sbox_5_T3), .Z0_t (SubBytesIns_Inst_Sbox_5_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M38), .B0_t (SubBytesIns_Inst_Sbox_5_T22), .Z0_t (SubBytesIns_Inst_Sbox_5_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M37), .B0_t (SubBytesIns_Inst_Sbox_5_T20), .Z0_t (SubBytesIns_Inst_Sbox_5_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M42), .B0_t (SubBytesIns_Inst_Sbox_5_T1), .Z0_t (SubBytesIns_Inst_Sbox_5_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M45), .B0_t (SubBytesIns_Inst_Sbox_5_T4), .Z0_t (SubBytesIns_Inst_Sbox_5_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M41), .B0_t (SubBytesIns_Inst_Sbox_5_T2), .Z0_t (SubBytesIns_Inst_Sbox_5_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M61), .B0_t (SubBytesIns_Inst_Sbox_5_M62), .Z0_t (SubBytesIns_Inst_Sbox_5_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M50), .B0_t (SubBytesIns_Inst_Sbox_5_M56), .Z0_t (SubBytesIns_Inst_Sbox_5_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M46), .B0_t (SubBytesIns_Inst_Sbox_5_M48), .Z0_t (SubBytesIns_Inst_Sbox_5_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M47), .B0_t (SubBytesIns_Inst_Sbox_5_M55), .Z0_t (SubBytesIns_Inst_Sbox_5_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M54), .B0_t (SubBytesIns_Inst_Sbox_5_M58), .Z0_t (SubBytesIns_Inst_Sbox_5_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M49), .B0_t (SubBytesIns_Inst_Sbox_5_M61), .Z0_t (SubBytesIns_Inst_Sbox_5_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M62), .B0_t (SubBytesIns_Inst_Sbox_5_L5), .Z0_t (SubBytesIns_Inst_Sbox_5_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M46), .B0_t (SubBytesIns_Inst_Sbox_5_L3), .Z0_t (SubBytesIns_Inst_Sbox_5_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M51), .B0_t (SubBytesIns_Inst_Sbox_5_M59), .Z0_t (SubBytesIns_Inst_Sbox_5_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M52), .B0_t (SubBytesIns_Inst_Sbox_5_M53), .Z0_t (SubBytesIns_Inst_Sbox_5_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M53), .B0_t (SubBytesIns_Inst_Sbox_5_L4), .Z0_t (SubBytesIns_Inst_Sbox_5_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M60), .B0_t (SubBytesIns_Inst_Sbox_5_L2), .Z0_t (SubBytesIns_Inst_Sbox_5_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M48), .B0_t (SubBytesIns_Inst_Sbox_5_M51), .Z0_t (SubBytesIns_Inst_Sbox_5_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M50), .B0_t (SubBytesIns_Inst_Sbox_5_L0), .Z0_t (SubBytesIns_Inst_Sbox_5_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M52), .B0_t (SubBytesIns_Inst_Sbox_5_M61), .Z0_t (SubBytesIns_Inst_Sbox_5_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M55), .B0_t (SubBytesIns_Inst_Sbox_5_L1), .Z0_t (SubBytesIns_Inst_Sbox_5_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M56), .B0_t (SubBytesIns_Inst_Sbox_5_L0), .Z0_t (SubBytesIns_Inst_Sbox_5_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M57), .B0_t (SubBytesIns_Inst_Sbox_5_L1), .Z0_t (SubBytesIns_Inst_Sbox_5_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M58), .B0_t (SubBytesIns_Inst_Sbox_5_L8), .Z0_t (SubBytesIns_Inst_Sbox_5_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_M63), .B0_t (SubBytesIns_Inst_Sbox_5_L4), .Z0_t (SubBytesIns_Inst_Sbox_5_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L0), .B0_t (SubBytesIns_Inst_Sbox_5_L1), .Z0_t (SubBytesIns_Inst_Sbox_5_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L1), .B0_t (SubBytesIns_Inst_Sbox_5_L7), .Z0_t (SubBytesIns_Inst_Sbox_5_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L3), .B0_t (SubBytesIns_Inst_Sbox_5_L12), .Z0_t (SubBytesIns_Inst_Sbox_5_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L18), .B0_t (SubBytesIns_Inst_Sbox_5_L2), .Z0_t (SubBytesIns_Inst_Sbox_5_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L15), .B0_t (SubBytesIns_Inst_Sbox_5_L9), .Z0_t (SubBytesIns_Inst_Sbox_5_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L6), .B0_t (SubBytesIns_Inst_Sbox_5_L10), .Z0_t (SubBytesIns_Inst_Sbox_5_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L7), .B0_t (SubBytesIns_Inst_Sbox_5_L9), .Z0_t (SubBytesIns_Inst_Sbox_5_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L8), .B0_t (SubBytesIns_Inst_Sbox_5_L10), .Z0_t (SubBytesIns_Inst_Sbox_5_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L11), .B0_t (SubBytesIns_Inst_Sbox_5_L14), .Z0_t (SubBytesIns_Inst_Sbox_5_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L11), .B0_t (SubBytesIns_Inst_Sbox_5_L17), .Z0_t (SubBytesIns_Inst_Sbox_5_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L6), .B0_t (SubBytesIns_Inst_Sbox_5_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L16), .B0_t (SubBytesIns_Inst_Sbox_5_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L19), .B0_t (SubBytesIns_Inst_Sbox_5_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L6), .B0_t (SubBytesIns_Inst_Sbox_5_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L20), .B0_t (SubBytesIns_Inst_Sbox_5_L22), .Z0_t (MixColumnsInput[107]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L25), .B0_t (SubBytesIns_Inst_Sbox_5_L29), .Z0_t (MixColumnsInput[106]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L13), .B0_t (SubBytesIns_Inst_Sbox_5_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_5_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_5_L6), .B0_t (SubBytesIns_Inst_Sbox_5_L23), .Z0_t (MixColumnsInput[104]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T1_U1 ( .A0_t (ciphertext[55]), .B0_t (ciphertext[52]), .Z0_t (SubBytesIns_Inst_Sbox_6_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T2_U1 ( .A0_t (ciphertext[55]), .B0_t (ciphertext[50]), .Z0_t (SubBytesIns_Inst_Sbox_6_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T3_U1 ( .A0_t (ciphertext[55]), .B0_t (ciphertext[49]), .Z0_t (SubBytesIns_Inst_Sbox_6_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T4_U1 ( .A0_t (ciphertext[52]), .B0_t (ciphertext[50]), .Z0_t (SubBytesIns_Inst_Sbox_6_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T5_U1 ( .A0_t (ciphertext[51]), .B0_t (ciphertext[49]), .Z0_t (SubBytesIns_Inst_Sbox_6_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T1), .B0_t (SubBytesIns_Inst_Sbox_6_T5), .Z0_t (SubBytesIns_Inst_Sbox_6_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T7_U1 ( .A0_t (ciphertext[54]), .B0_t (ciphertext[53]), .Z0_t (SubBytesIns_Inst_Sbox_6_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T8_U1 ( .A0_t (ciphertext[48]), .B0_t (SubBytesIns_Inst_Sbox_6_T6), .Z0_t (SubBytesIns_Inst_Sbox_6_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T9_U1 ( .A0_t (ciphertext[48]), .B0_t (SubBytesIns_Inst_Sbox_6_T7), .Z0_t (SubBytesIns_Inst_Sbox_6_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T6), .B0_t (SubBytesIns_Inst_Sbox_6_T7), .Z0_t (SubBytesIns_Inst_Sbox_6_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T11_U1 ( .A0_t (ciphertext[54]), .B0_t (ciphertext[50]), .Z0_t (SubBytesIns_Inst_Sbox_6_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T12_U1 ( .A0_t (ciphertext[53]), .B0_t (ciphertext[50]), .Z0_t (SubBytesIns_Inst_Sbox_6_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T3), .B0_t (SubBytesIns_Inst_Sbox_6_T4), .Z0_t (SubBytesIns_Inst_Sbox_6_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T6), .B0_t (SubBytesIns_Inst_Sbox_6_T11), .Z0_t (SubBytesIns_Inst_Sbox_6_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T5), .B0_t (SubBytesIns_Inst_Sbox_6_T11), .Z0_t (SubBytesIns_Inst_Sbox_6_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T5), .B0_t (SubBytesIns_Inst_Sbox_6_T12), .Z0_t (SubBytesIns_Inst_Sbox_6_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T9), .B0_t (SubBytesIns_Inst_Sbox_6_T16), .Z0_t (SubBytesIns_Inst_Sbox_6_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T18_U1 ( .A0_t (ciphertext[52]), .B0_t (ciphertext[48]), .Z0_t (SubBytesIns_Inst_Sbox_6_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T7), .B0_t (SubBytesIns_Inst_Sbox_6_T18), .Z0_t (SubBytesIns_Inst_Sbox_6_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T1), .B0_t (SubBytesIns_Inst_Sbox_6_T19), .Z0_t (SubBytesIns_Inst_Sbox_6_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T21_U1 ( .A0_t (ciphertext[49]), .B0_t (ciphertext[48]), .Z0_t (SubBytesIns_Inst_Sbox_6_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T7), .B0_t (SubBytesIns_Inst_Sbox_6_T21), .Z0_t (SubBytesIns_Inst_Sbox_6_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T2), .B0_t (SubBytesIns_Inst_Sbox_6_T22), .Z0_t (SubBytesIns_Inst_Sbox_6_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T2), .B0_t (SubBytesIns_Inst_Sbox_6_T10), .Z0_t (SubBytesIns_Inst_Sbox_6_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T20), .B0_t (SubBytesIns_Inst_Sbox_6_T17), .Z0_t (SubBytesIns_Inst_Sbox_6_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T3), .B0_t (SubBytesIns_Inst_Sbox_6_T16), .Z0_t (SubBytesIns_Inst_Sbox_6_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T1), .B0_t (SubBytesIns_Inst_Sbox_6_T12), .Z0_t (SubBytesIns_Inst_Sbox_6_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T13), .B0_t (SubBytesIns_Inst_Sbox_6_T6), .Z0_t (SubBytesIns_Inst_Sbox_6_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T23), .B0_t (SubBytesIns_Inst_Sbox_6_T8), .Z0_t (SubBytesIns_Inst_Sbox_6_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T14), .B0_t (SubBytesIns_Inst_Sbox_6_M1), .Z0_t (SubBytesIns_Inst_Sbox_6_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T19), .B0_t (ciphertext[48]), .Z0_t (SubBytesIns_Inst_Sbox_6_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M4), .B0_t (SubBytesIns_Inst_Sbox_6_M1), .Z0_t (SubBytesIns_Inst_Sbox_6_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T3), .B0_t (SubBytesIns_Inst_Sbox_6_T16), .Z0_t (SubBytesIns_Inst_Sbox_6_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T22), .B0_t (SubBytesIns_Inst_Sbox_6_T9), .Z0_t (SubBytesIns_Inst_Sbox_6_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T26), .B0_t (SubBytesIns_Inst_Sbox_6_M6), .Z0_t (SubBytesIns_Inst_Sbox_6_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T20), .B0_t (SubBytesIns_Inst_Sbox_6_T17), .Z0_t (SubBytesIns_Inst_Sbox_6_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M9), .B0_t (SubBytesIns_Inst_Sbox_6_M6), .Z0_t (SubBytesIns_Inst_Sbox_6_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T1), .B0_t (SubBytesIns_Inst_Sbox_6_T15), .Z0_t (SubBytesIns_Inst_Sbox_6_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T4), .B0_t (SubBytesIns_Inst_Sbox_6_T27), .Z0_t (SubBytesIns_Inst_Sbox_6_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M12), .B0_t (SubBytesIns_Inst_Sbox_6_M11), .Z0_t (SubBytesIns_Inst_Sbox_6_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_T2), .B0_t (SubBytesIns_Inst_Sbox_6_T10), .Z0_t (SubBytesIns_Inst_Sbox_6_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M14), .B0_t (SubBytesIns_Inst_Sbox_6_M11), .Z0_t (SubBytesIns_Inst_Sbox_6_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M3), .B0_t (SubBytesIns_Inst_Sbox_6_M2), .Z0_t (SubBytesIns_Inst_Sbox_6_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M5), .B0_t (SubBytesIns_Inst_Sbox_6_T24), .Z0_t (SubBytesIns_Inst_Sbox_6_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M8), .B0_t (SubBytesIns_Inst_Sbox_6_M7), .Z0_t (SubBytesIns_Inst_Sbox_6_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M10), .B0_t (SubBytesIns_Inst_Sbox_6_M15), .Z0_t (SubBytesIns_Inst_Sbox_6_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M16), .B0_t (SubBytesIns_Inst_Sbox_6_M13), .Z0_t (SubBytesIns_Inst_Sbox_6_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M17), .B0_t (SubBytesIns_Inst_Sbox_6_M15), .Z0_t (SubBytesIns_Inst_Sbox_6_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M18), .B0_t (SubBytesIns_Inst_Sbox_6_M13), .Z0_t (SubBytesIns_Inst_Sbox_6_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M19), .B0_t (SubBytesIns_Inst_Sbox_6_T25), .Z0_t (SubBytesIns_Inst_Sbox_6_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M22), .B0_t (SubBytesIns_Inst_Sbox_6_M23), .Z0_t (SubBytesIns_Inst_Sbox_6_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M22), .B0_t (SubBytesIns_Inst_Sbox_6_M20), .Z0_t (SubBytesIns_Inst_Sbox_6_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M21), .B0_t (SubBytesIns_Inst_Sbox_6_M25), .Z0_t (SubBytesIns_Inst_Sbox_6_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M20), .B0_t (SubBytesIns_Inst_Sbox_6_M21), .Z0_t (SubBytesIns_Inst_Sbox_6_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M23), .B0_t (SubBytesIns_Inst_Sbox_6_M25), .Z0_t (SubBytesIns_Inst_Sbox_6_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M28), .B0_t (SubBytesIns_Inst_Sbox_6_M27), .Z0_t (SubBytesIns_Inst_Sbox_6_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M26), .B0_t (SubBytesIns_Inst_Sbox_6_M24), .Z0_t (SubBytesIns_Inst_Sbox_6_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M20), .B0_t (SubBytesIns_Inst_Sbox_6_M23), .Z0_t (SubBytesIns_Inst_Sbox_6_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M27), .B0_t (SubBytesIns_Inst_Sbox_6_M31), .Z0_t (SubBytesIns_Inst_Sbox_6_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M27), .B0_t (SubBytesIns_Inst_Sbox_6_M25), .Z0_t (SubBytesIns_Inst_Sbox_6_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M21), .B0_t (SubBytesIns_Inst_Sbox_6_M22), .Z0_t (SubBytesIns_Inst_Sbox_6_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M24), .B0_t (SubBytesIns_Inst_Sbox_6_M34), .Z0_t (SubBytesIns_Inst_Sbox_6_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M24), .B0_t (SubBytesIns_Inst_Sbox_6_M25), .Z0_t (SubBytesIns_Inst_Sbox_6_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M21), .B0_t (SubBytesIns_Inst_Sbox_6_M29), .Z0_t (SubBytesIns_Inst_Sbox_6_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M32), .B0_t (SubBytesIns_Inst_Sbox_6_M33), .Z0_t (SubBytesIns_Inst_Sbox_6_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M23), .B0_t (SubBytesIns_Inst_Sbox_6_M30), .Z0_t (SubBytesIns_Inst_Sbox_6_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M35), .B0_t (SubBytesIns_Inst_Sbox_6_M36), .Z0_t (SubBytesIns_Inst_Sbox_6_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M38), .B0_t (SubBytesIns_Inst_Sbox_6_M40), .Z0_t (SubBytesIns_Inst_Sbox_6_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M37), .B0_t (SubBytesIns_Inst_Sbox_6_M39), .Z0_t (SubBytesIns_Inst_Sbox_6_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M37), .B0_t (SubBytesIns_Inst_Sbox_6_M38), .Z0_t (SubBytesIns_Inst_Sbox_6_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M39), .B0_t (SubBytesIns_Inst_Sbox_6_M40), .Z0_t (SubBytesIns_Inst_Sbox_6_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M42), .B0_t (SubBytesIns_Inst_Sbox_6_M41), .Z0_t (SubBytesIns_Inst_Sbox_6_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M44), .B0_t (SubBytesIns_Inst_Sbox_6_T6), .Z0_t (SubBytesIns_Inst_Sbox_6_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M40), .B0_t (SubBytesIns_Inst_Sbox_6_T8), .Z0_t (SubBytesIns_Inst_Sbox_6_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M39), .B0_t (ciphertext[48]), .Z0_t (SubBytesIns_Inst_Sbox_6_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M43), .B0_t (SubBytesIns_Inst_Sbox_6_T16), .Z0_t (SubBytesIns_Inst_Sbox_6_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M38), .B0_t (SubBytesIns_Inst_Sbox_6_T9), .Z0_t (SubBytesIns_Inst_Sbox_6_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M37), .B0_t (SubBytesIns_Inst_Sbox_6_T17), .Z0_t (SubBytesIns_Inst_Sbox_6_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M42), .B0_t (SubBytesIns_Inst_Sbox_6_T15), .Z0_t (SubBytesIns_Inst_Sbox_6_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M45), .B0_t (SubBytesIns_Inst_Sbox_6_T27), .Z0_t (SubBytesIns_Inst_Sbox_6_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M41), .B0_t (SubBytesIns_Inst_Sbox_6_T10), .Z0_t (SubBytesIns_Inst_Sbox_6_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M44), .B0_t (SubBytesIns_Inst_Sbox_6_T13), .Z0_t (SubBytesIns_Inst_Sbox_6_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M40), .B0_t (SubBytesIns_Inst_Sbox_6_T23), .Z0_t (SubBytesIns_Inst_Sbox_6_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M39), .B0_t (SubBytesIns_Inst_Sbox_6_T19), .Z0_t (SubBytesIns_Inst_Sbox_6_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M43), .B0_t (SubBytesIns_Inst_Sbox_6_T3), .Z0_t (SubBytesIns_Inst_Sbox_6_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M38), .B0_t (SubBytesIns_Inst_Sbox_6_T22), .Z0_t (SubBytesIns_Inst_Sbox_6_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M37), .B0_t (SubBytesIns_Inst_Sbox_6_T20), .Z0_t (SubBytesIns_Inst_Sbox_6_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M42), .B0_t (SubBytesIns_Inst_Sbox_6_T1), .Z0_t (SubBytesIns_Inst_Sbox_6_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M45), .B0_t (SubBytesIns_Inst_Sbox_6_T4), .Z0_t (SubBytesIns_Inst_Sbox_6_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M41), .B0_t (SubBytesIns_Inst_Sbox_6_T2), .Z0_t (SubBytesIns_Inst_Sbox_6_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M61), .B0_t (SubBytesIns_Inst_Sbox_6_M62), .Z0_t (SubBytesIns_Inst_Sbox_6_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M50), .B0_t (SubBytesIns_Inst_Sbox_6_M56), .Z0_t (SubBytesIns_Inst_Sbox_6_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M46), .B0_t (SubBytesIns_Inst_Sbox_6_M48), .Z0_t (SubBytesIns_Inst_Sbox_6_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M47), .B0_t (SubBytesIns_Inst_Sbox_6_M55), .Z0_t (SubBytesIns_Inst_Sbox_6_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M54), .B0_t (SubBytesIns_Inst_Sbox_6_M58), .Z0_t (SubBytesIns_Inst_Sbox_6_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M49), .B0_t (SubBytesIns_Inst_Sbox_6_M61), .Z0_t (SubBytesIns_Inst_Sbox_6_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M62), .B0_t (SubBytesIns_Inst_Sbox_6_L5), .Z0_t (SubBytesIns_Inst_Sbox_6_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M46), .B0_t (SubBytesIns_Inst_Sbox_6_L3), .Z0_t (SubBytesIns_Inst_Sbox_6_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M51), .B0_t (SubBytesIns_Inst_Sbox_6_M59), .Z0_t (SubBytesIns_Inst_Sbox_6_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M52), .B0_t (SubBytesIns_Inst_Sbox_6_M53), .Z0_t (SubBytesIns_Inst_Sbox_6_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M53), .B0_t (SubBytesIns_Inst_Sbox_6_L4), .Z0_t (SubBytesIns_Inst_Sbox_6_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M60), .B0_t (SubBytesIns_Inst_Sbox_6_L2), .Z0_t (SubBytesIns_Inst_Sbox_6_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M48), .B0_t (SubBytesIns_Inst_Sbox_6_M51), .Z0_t (SubBytesIns_Inst_Sbox_6_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M50), .B0_t (SubBytesIns_Inst_Sbox_6_L0), .Z0_t (SubBytesIns_Inst_Sbox_6_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M52), .B0_t (SubBytesIns_Inst_Sbox_6_M61), .Z0_t (SubBytesIns_Inst_Sbox_6_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M55), .B0_t (SubBytesIns_Inst_Sbox_6_L1), .Z0_t (SubBytesIns_Inst_Sbox_6_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M56), .B0_t (SubBytesIns_Inst_Sbox_6_L0), .Z0_t (SubBytesIns_Inst_Sbox_6_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M57), .B0_t (SubBytesIns_Inst_Sbox_6_L1), .Z0_t (SubBytesIns_Inst_Sbox_6_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M58), .B0_t (SubBytesIns_Inst_Sbox_6_L8), .Z0_t (SubBytesIns_Inst_Sbox_6_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_M63), .B0_t (SubBytesIns_Inst_Sbox_6_L4), .Z0_t (SubBytesIns_Inst_Sbox_6_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L0), .B0_t (SubBytesIns_Inst_Sbox_6_L1), .Z0_t (SubBytesIns_Inst_Sbox_6_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L1), .B0_t (SubBytesIns_Inst_Sbox_6_L7), .Z0_t (SubBytesIns_Inst_Sbox_6_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L3), .B0_t (SubBytesIns_Inst_Sbox_6_L12), .Z0_t (SubBytesIns_Inst_Sbox_6_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L18), .B0_t (SubBytesIns_Inst_Sbox_6_L2), .Z0_t (SubBytesIns_Inst_Sbox_6_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L15), .B0_t (SubBytesIns_Inst_Sbox_6_L9), .Z0_t (SubBytesIns_Inst_Sbox_6_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L6), .B0_t (SubBytesIns_Inst_Sbox_6_L10), .Z0_t (SubBytesIns_Inst_Sbox_6_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L7), .B0_t (SubBytesIns_Inst_Sbox_6_L9), .Z0_t (SubBytesIns_Inst_Sbox_6_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L8), .B0_t (SubBytesIns_Inst_Sbox_6_L10), .Z0_t (SubBytesIns_Inst_Sbox_6_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L11), .B0_t (SubBytesIns_Inst_Sbox_6_L14), .Z0_t (SubBytesIns_Inst_Sbox_6_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L11), .B0_t (SubBytesIns_Inst_Sbox_6_L17), .Z0_t (SubBytesIns_Inst_Sbox_6_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L6), .B0_t (SubBytesIns_Inst_Sbox_6_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L16), .B0_t (SubBytesIns_Inst_Sbox_6_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L19), .B0_t (SubBytesIns_Inst_Sbox_6_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L6), .B0_t (SubBytesIns_Inst_Sbox_6_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L20), .B0_t (SubBytesIns_Inst_Sbox_6_L22), .Z0_t (MixColumnsInput[83]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L25), .B0_t (SubBytesIns_Inst_Sbox_6_L29), .Z0_t (MixColumnsInput[82]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L13), .B0_t (SubBytesIns_Inst_Sbox_6_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_6_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_6_L6), .B0_t (SubBytesIns_Inst_Sbox_6_L23), .Z0_t (MixColumnsInput[80]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T1_U1 ( .A0_t (ciphertext[63]), .B0_t (ciphertext[60]), .Z0_t (SubBytesIns_Inst_Sbox_7_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T2_U1 ( .A0_t (ciphertext[63]), .B0_t (ciphertext[58]), .Z0_t (SubBytesIns_Inst_Sbox_7_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T3_U1 ( .A0_t (ciphertext[63]), .B0_t (ciphertext[57]), .Z0_t (SubBytesIns_Inst_Sbox_7_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T4_U1 ( .A0_t (ciphertext[60]), .B0_t (ciphertext[58]), .Z0_t (SubBytesIns_Inst_Sbox_7_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T5_U1 ( .A0_t (ciphertext[59]), .B0_t (ciphertext[57]), .Z0_t (SubBytesIns_Inst_Sbox_7_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T1), .B0_t (SubBytesIns_Inst_Sbox_7_T5), .Z0_t (SubBytesIns_Inst_Sbox_7_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T7_U1 ( .A0_t (ciphertext[62]), .B0_t (ciphertext[61]), .Z0_t (SubBytesIns_Inst_Sbox_7_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T8_U1 ( .A0_t (ciphertext[56]), .B0_t (SubBytesIns_Inst_Sbox_7_T6), .Z0_t (SubBytesIns_Inst_Sbox_7_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T9_U1 ( .A0_t (ciphertext[56]), .B0_t (SubBytesIns_Inst_Sbox_7_T7), .Z0_t (SubBytesIns_Inst_Sbox_7_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T6), .B0_t (SubBytesIns_Inst_Sbox_7_T7), .Z0_t (SubBytesIns_Inst_Sbox_7_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T11_U1 ( .A0_t (ciphertext[62]), .B0_t (ciphertext[58]), .Z0_t (SubBytesIns_Inst_Sbox_7_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T12_U1 ( .A0_t (ciphertext[61]), .B0_t (ciphertext[58]), .Z0_t (SubBytesIns_Inst_Sbox_7_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T3), .B0_t (SubBytesIns_Inst_Sbox_7_T4), .Z0_t (SubBytesIns_Inst_Sbox_7_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T6), .B0_t (SubBytesIns_Inst_Sbox_7_T11), .Z0_t (SubBytesIns_Inst_Sbox_7_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T5), .B0_t (SubBytesIns_Inst_Sbox_7_T11), .Z0_t (SubBytesIns_Inst_Sbox_7_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T5), .B0_t (SubBytesIns_Inst_Sbox_7_T12), .Z0_t (SubBytesIns_Inst_Sbox_7_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T9), .B0_t (SubBytesIns_Inst_Sbox_7_T16), .Z0_t (SubBytesIns_Inst_Sbox_7_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T18_U1 ( .A0_t (ciphertext[60]), .B0_t (ciphertext[56]), .Z0_t (SubBytesIns_Inst_Sbox_7_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T7), .B0_t (SubBytesIns_Inst_Sbox_7_T18), .Z0_t (SubBytesIns_Inst_Sbox_7_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T1), .B0_t (SubBytesIns_Inst_Sbox_7_T19), .Z0_t (SubBytesIns_Inst_Sbox_7_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T21_U1 ( .A0_t (ciphertext[57]), .B0_t (ciphertext[56]), .Z0_t (SubBytesIns_Inst_Sbox_7_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T7), .B0_t (SubBytesIns_Inst_Sbox_7_T21), .Z0_t (SubBytesIns_Inst_Sbox_7_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T2), .B0_t (SubBytesIns_Inst_Sbox_7_T22), .Z0_t (SubBytesIns_Inst_Sbox_7_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T2), .B0_t (SubBytesIns_Inst_Sbox_7_T10), .Z0_t (SubBytesIns_Inst_Sbox_7_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T20), .B0_t (SubBytesIns_Inst_Sbox_7_T17), .Z0_t (SubBytesIns_Inst_Sbox_7_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T3), .B0_t (SubBytesIns_Inst_Sbox_7_T16), .Z0_t (SubBytesIns_Inst_Sbox_7_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T1), .B0_t (SubBytesIns_Inst_Sbox_7_T12), .Z0_t (SubBytesIns_Inst_Sbox_7_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T13), .B0_t (SubBytesIns_Inst_Sbox_7_T6), .Z0_t (SubBytesIns_Inst_Sbox_7_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T23), .B0_t (SubBytesIns_Inst_Sbox_7_T8), .Z0_t (SubBytesIns_Inst_Sbox_7_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T14), .B0_t (SubBytesIns_Inst_Sbox_7_M1), .Z0_t (SubBytesIns_Inst_Sbox_7_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T19), .B0_t (ciphertext[56]), .Z0_t (SubBytesIns_Inst_Sbox_7_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M4), .B0_t (SubBytesIns_Inst_Sbox_7_M1), .Z0_t (SubBytesIns_Inst_Sbox_7_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T3), .B0_t (SubBytesIns_Inst_Sbox_7_T16), .Z0_t (SubBytesIns_Inst_Sbox_7_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T22), .B0_t (SubBytesIns_Inst_Sbox_7_T9), .Z0_t (SubBytesIns_Inst_Sbox_7_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T26), .B0_t (SubBytesIns_Inst_Sbox_7_M6), .Z0_t (SubBytesIns_Inst_Sbox_7_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T20), .B0_t (SubBytesIns_Inst_Sbox_7_T17), .Z0_t (SubBytesIns_Inst_Sbox_7_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M9), .B0_t (SubBytesIns_Inst_Sbox_7_M6), .Z0_t (SubBytesIns_Inst_Sbox_7_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T1), .B0_t (SubBytesIns_Inst_Sbox_7_T15), .Z0_t (SubBytesIns_Inst_Sbox_7_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T4), .B0_t (SubBytesIns_Inst_Sbox_7_T27), .Z0_t (SubBytesIns_Inst_Sbox_7_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M12), .B0_t (SubBytesIns_Inst_Sbox_7_M11), .Z0_t (SubBytesIns_Inst_Sbox_7_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_T2), .B0_t (SubBytesIns_Inst_Sbox_7_T10), .Z0_t (SubBytesIns_Inst_Sbox_7_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M14), .B0_t (SubBytesIns_Inst_Sbox_7_M11), .Z0_t (SubBytesIns_Inst_Sbox_7_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M3), .B0_t (SubBytesIns_Inst_Sbox_7_M2), .Z0_t (SubBytesIns_Inst_Sbox_7_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M5), .B0_t (SubBytesIns_Inst_Sbox_7_T24), .Z0_t (SubBytesIns_Inst_Sbox_7_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M8), .B0_t (SubBytesIns_Inst_Sbox_7_M7), .Z0_t (SubBytesIns_Inst_Sbox_7_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M10), .B0_t (SubBytesIns_Inst_Sbox_7_M15), .Z0_t (SubBytesIns_Inst_Sbox_7_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M16), .B0_t (SubBytesIns_Inst_Sbox_7_M13), .Z0_t (SubBytesIns_Inst_Sbox_7_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M17), .B0_t (SubBytesIns_Inst_Sbox_7_M15), .Z0_t (SubBytesIns_Inst_Sbox_7_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M18), .B0_t (SubBytesIns_Inst_Sbox_7_M13), .Z0_t (SubBytesIns_Inst_Sbox_7_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M19), .B0_t (SubBytesIns_Inst_Sbox_7_T25), .Z0_t (SubBytesIns_Inst_Sbox_7_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M22), .B0_t (SubBytesIns_Inst_Sbox_7_M23), .Z0_t (SubBytesIns_Inst_Sbox_7_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M22), .B0_t (SubBytesIns_Inst_Sbox_7_M20), .Z0_t (SubBytesIns_Inst_Sbox_7_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M21), .B0_t (SubBytesIns_Inst_Sbox_7_M25), .Z0_t (SubBytesIns_Inst_Sbox_7_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M20), .B0_t (SubBytesIns_Inst_Sbox_7_M21), .Z0_t (SubBytesIns_Inst_Sbox_7_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M23), .B0_t (SubBytesIns_Inst_Sbox_7_M25), .Z0_t (SubBytesIns_Inst_Sbox_7_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M28), .B0_t (SubBytesIns_Inst_Sbox_7_M27), .Z0_t (SubBytesIns_Inst_Sbox_7_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M26), .B0_t (SubBytesIns_Inst_Sbox_7_M24), .Z0_t (SubBytesIns_Inst_Sbox_7_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M20), .B0_t (SubBytesIns_Inst_Sbox_7_M23), .Z0_t (SubBytesIns_Inst_Sbox_7_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M27), .B0_t (SubBytesIns_Inst_Sbox_7_M31), .Z0_t (SubBytesIns_Inst_Sbox_7_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M27), .B0_t (SubBytesIns_Inst_Sbox_7_M25), .Z0_t (SubBytesIns_Inst_Sbox_7_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M21), .B0_t (SubBytesIns_Inst_Sbox_7_M22), .Z0_t (SubBytesIns_Inst_Sbox_7_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M24), .B0_t (SubBytesIns_Inst_Sbox_7_M34), .Z0_t (SubBytesIns_Inst_Sbox_7_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M24), .B0_t (SubBytesIns_Inst_Sbox_7_M25), .Z0_t (SubBytesIns_Inst_Sbox_7_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M21), .B0_t (SubBytesIns_Inst_Sbox_7_M29), .Z0_t (SubBytesIns_Inst_Sbox_7_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M32), .B0_t (SubBytesIns_Inst_Sbox_7_M33), .Z0_t (SubBytesIns_Inst_Sbox_7_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M23), .B0_t (SubBytesIns_Inst_Sbox_7_M30), .Z0_t (SubBytesIns_Inst_Sbox_7_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M35), .B0_t (SubBytesIns_Inst_Sbox_7_M36), .Z0_t (SubBytesIns_Inst_Sbox_7_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M38), .B0_t (SubBytesIns_Inst_Sbox_7_M40), .Z0_t (SubBytesIns_Inst_Sbox_7_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M37), .B0_t (SubBytesIns_Inst_Sbox_7_M39), .Z0_t (SubBytesIns_Inst_Sbox_7_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M37), .B0_t (SubBytesIns_Inst_Sbox_7_M38), .Z0_t (SubBytesIns_Inst_Sbox_7_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M39), .B0_t (SubBytesIns_Inst_Sbox_7_M40), .Z0_t (SubBytesIns_Inst_Sbox_7_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M42), .B0_t (SubBytesIns_Inst_Sbox_7_M41), .Z0_t (SubBytesIns_Inst_Sbox_7_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M44), .B0_t (SubBytesIns_Inst_Sbox_7_T6), .Z0_t (SubBytesIns_Inst_Sbox_7_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M40), .B0_t (SubBytesIns_Inst_Sbox_7_T8), .Z0_t (SubBytesIns_Inst_Sbox_7_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M39), .B0_t (ciphertext[56]), .Z0_t (SubBytesIns_Inst_Sbox_7_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M43), .B0_t (SubBytesIns_Inst_Sbox_7_T16), .Z0_t (SubBytesIns_Inst_Sbox_7_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M38), .B0_t (SubBytesIns_Inst_Sbox_7_T9), .Z0_t (SubBytesIns_Inst_Sbox_7_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M37), .B0_t (SubBytesIns_Inst_Sbox_7_T17), .Z0_t (SubBytesIns_Inst_Sbox_7_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M42), .B0_t (SubBytesIns_Inst_Sbox_7_T15), .Z0_t (SubBytesIns_Inst_Sbox_7_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M45), .B0_t (SubBytesIns_Inst_Sbox_7_T27), .Z0_t (SubBytesIns_Inst_Sbox_7_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M41), .B0_t (SubBytesIns_Inst_Sbox_7_T10), .Z0_t (SubBytesIns_Inst_Sbox_7_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M44), .B0_t (SubBytesIns_Inst_Sbox_7_T13), .Z0_t (SubBytesIns_Inst_Sbox_7_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M40), .B0_t (SubBytesIns_Inst_Sbox_7_T23), .Z0_t (SubBytesIns_Inst_Sbox_7_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M39), .B0_t (SubBytesIns_Inst_Sbox_7_T19), .Z0_t (SubBytesIns_Inst_Sbox_7_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M43), .B0_t (SubBytesIns_Inst_Sbox_7_T3), .Z0_t (SubBytesIns_Inst_Sbox_7_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M38), .B0_t (SubBytesIns_Inst_Sbox_7_T22), .Z0_t (SubBytesIns_Inst_Sbox_7_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M37), .B0_t (SubBytesIns_Inst_Sbox_7_T20), .Z0_t (SubBytesIns_Inst_Sbox_7_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M42), .B0_t (SubBytesIns_Inst_Sbox_7_T1), .Z0_t (SubBytesIns_Inst_Sbox_7_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M45), .B0_t (SubBytesIns_Inst_Sbox_7_T4), .Z0_t (SubBytesIns_Inst_Sbox_7_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M41), .B0_t (SubBytesIns_Inst_Sbox_7_T2), .Z0_t (SubBytesIns_Inst_Sbox_7_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M61), .B0_t (SubBytesIns_Inst_Sbox_7_M62), .Z0_t (SubBytesIns_Inst_Sbox_7_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M50), .B0_t (SubBytesIns_Inst_Sbox_7_M56), .Z0_t (SubBytesIns_Inst_Sbox_7_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M46), .B0_t (SubBytesIns_Inst_Sbox_7_M48), .Z0_t (SubBytesIns_Inst_Sbox_7_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M47), .B0_t (SubBytesIns_Inst_Sbox_7_M55), .Z0_t (SubBytesIns_Inst_Sbox_7_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M54), .B0_t (SubBytesIns_Inst_Sbox_7_M58), .Z0_t (SubBytesIns_Inst_Sbox_7_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M49), .B0_t (SubBytesIns_Inst_Sbox_7_M61), .Z0_t (SubBytesIns_Inst_Sbox_7_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M62), .B0_t (SubBytesIns_Inst_Sbox_7_L5), .Z0_t (SubBytesIns_Inst_Sbox_7_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M46), .B0_t (SubBytesIns_Inst_Sbox_7_L3), .Z0_t (SubBytesIns_Inst_Sbox_7_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M51), .B0_t (SubBytesIns_Inst_Sbox_7_M59), .Z0_t (SubBytesIns_Inst_Sbox_7_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M52), .B0_t (SubBytesIns_Inst_Sbox_7_M53), .Z0_t (SubBytesIns_Inst_Sbox_7_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M53), .B0_t (SubBytesIns_Inst_Sbox_7_L4), .Z0_t (SubBytesIns_Inst_Sbox_7_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M60), .B0_t (SubBytesIns_Inst_Sbox_7_L2), .Z0_t (SubBytesIns_Inst_Sbox_7_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M48), .B0_t (SubBytesIns_Inst_Sbox_7_M51), .Z0_t (SubBytesIns_Inst_Sbox_7_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M50), .B0_t (SubBytesIns_Inst_Sbox_7_L0), .Z0_t (SubBytesIns_Inst_Sbox_7_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M52), .B0_t (SubBytesIns_Inst_Sbox_7_M61), .Z0_t (SubBytesIns_Inst_Sbox_7_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M55), .B0_t (SubBytesIns_Inst_Sbox_7_L1), .Z0_t (SubBytesIns_Inst_Sbox_7_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M56), .B0_t (SubBytesIns_Inst_Sbox_7_L0), .Z0_t (SubBytesIns_Inst_Sbox_7_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M57), .B0_t (SubBytesIns_Inst_Sbox_7_L1), .Z0_t (SubBytesIns_Inst_Sbox_7_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M58), .B0_t (SubBytesIns_Inst_Sbox_7_L8), .Z0_t (SubBytesIns_Inst_Sbox_7_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_M63), .B0_t (SubBytesIns_Inst_Sbox_7_L4), .Z0_t (SubBytesIns_Inst_Sbox_7_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L0), .B0_t (SubBytesIns_Inst_Sbox_7_L1), .Z0_t (SubBytesIns_Inst_Sbox_7_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L1), .B0_t (SubBytesIns_Inst_Sbox_7_L7), .Z0_t (SubBytesIns_Inst_Sbox_7_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L3), .B0_t (SubBytesIns_Inst_Sbox_7_L12), .Z0_t (SubBytesIns_Inst_Sbox_7_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L18), .B0_t (SubBytesIns_Inst_Sbox_7_L2), .Z0_t (SubBytesIns_Inst_Sbox_7_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L15), .B0_t (SubBytesIns_Inst_Sbox_7_L9), .Z0_t (SubBytesIns_Inst_Sbox_7_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L6), .B0_t (SubBytesIns_Inst_Sbox_7_L10), .Z0_t (SubBytesIns_Inst_Sbox_7_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L7), .B0_t (SubBytesIns_Inst_Sbox_7_L9), .Z0_t (SubBytesIns_Inst_Sbox_7_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L8), .B0_t (SubBytesIns_Inst_Sbox_7_L10), .Z0_t (SubBytesIns_Inst_Sbox_7_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L11), .B0_t (SubBytesIns_Inst_Sbox_7_L14), .Z0_t (SubBytesIns_Inst_Sbox_7_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L11), .B0_t (SubBytesIns_Inst_Sbox_7_L17), .Z0_t (SubBytesIns_Inst_Sbox_7_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L6), .B0_t (SubBytesIns_Inst_Sbox_7_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L16), .B0_t (SubBytesIns_Inst_Sbox_7_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L19), .B0_t (SubBytesIns_Inst_Sbox_7_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L6), .B0_t (SubBytesIns_Inst_Sbox_7_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L20), .B0_t (SubBytesIns_Inst_Sbox_7_L22), .Z0_t (MixColumnsInput[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L25), .B0_t (SubBytesIns_Inst_Sbox_7_L29), .Z0_t (MixColumnsInput[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L13), .B0_t (SubBytesIns_Inst_Sbox_7_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_7_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_7_L6), .B0_t (SubBytesIns_Inst_Sbox_7_L23), .Z0_t (MixColumnsInput[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T1_U1 ( .A0_t (ciphertext[71]), .B0_t (ciphertext[68]), .Z0_t (SubBytesIns_Inst_Sbox_8_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T2_U1 ( .A0_t (ciphertext[71]), .B0_t (ciphertext[66]), .Z0_t (SubBytesIns_Inst_Sbox_8_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T3_U1 ( .A0_t (ciphertext[71]), .B0_t (ciphertext[65]), .Z0_t (SubBytesIns_Inst_Sbox_8_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T4_U1 ( .A0_t (ciphertext[68]), .B0_t (ciphertext[66]), .Z0_t (SubBytesIns_Inst_Sbox_8_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T5_U1 ( .A0_t (ciphertext[67]), .B0_t (ciphertext[65]), .Z0_t (SubBytesIns_Inst_Sbox_8_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T1), .B0_t (SubBytesIns_Inst_Sbox_8_T5), .Z0_t (SubBytesIns_Inst_Sbox_8_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T7_U1 ( .A0_t (ciphertext[70]), .B0_t (ciphertext[69]), .Z0_t (SubBytesIns_Inst_Sbox_8_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T8_U1 ( .A0_t (ciphertext[64]), .B0_t (SubBytesIns_Inst_Sbox_8_T6), .Z0_t (SubBytesIns_Inst_Sbox_8_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T9_U1 ( .A0_t (ciphertext[64]), .B0_t (SubBytesIns_Inst_Sbox_8_T7), .Z0_t (SubBytesIns_Inst_Sbox_8_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T6), .B0_t (SubBytesIns_Inst_Sbox_8_T7), .Z0_t (SubBytesIns_Inst_Sbox_8_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T11_U1 ( .A0_t (ciphertext[70]), .B0_t (ciphertext[66]), .Z0_t (SubBytesIns_Inst_Sbox_8_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T12_U1 ( .A0_t (ciphertext[69]), .B0_t (ciphertext[66]), .Z0_t (SubBytesIns_Inst_Sbox_8_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T3), .B0_t (SubBytesIns_Inst_Sbox_8_T4), .Z0_t (SubBytesIns_Inst_Sbox_8_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T6), .B0_t (SubBytesIns_Inst_Sbox_8_T11), .Z0_t (SubBytesIns_Inst_Sbox_8_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T5), .B0_t (SubBytesIns_Inst_Sbox_8_T11), .Z0_t (SubBytesIns_Inst_Sbox_8_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T5), .B0_t (SubBytesIns_Inst_Sbox_8_T12), .Z0_t (SubBytesIns_Inst_Sbox_8_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T9), .B0_t (SubBytesIns_Inst_Sbox_8_T16), .Z0_t (SubBytesIns_Inst_Sbox_8_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T18_U1 ( .A0_t (ciphertext[68]), .B0_t (ciphertext[64]), .Z0_t (SubBytesIns_Inst_Sbox_8_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T7), .B0_t (SubBytesIns_Inst_Sbox_8_T18), .Z0_t (SubBytesIns_Inst_Sbox_8_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T1), .B0_t (SubBytesIns_Inst_Sbox_8_T19), .Z0_t (SubBytesIns_Inst_Sbox_8_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T21_U1 ( .A0_t (ciphertext[65]), .B0_t (ciphertext[64]), .Z0_t (SubBytesIns_Inst_Sbox_8_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T7), .B0_t (SubBytesIns_Inst_Sbox_8_T21), .Z0_t (SubBytesIns_Inst_Sbox_8_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T2), .B0_t (SubBytesIns_Inst_Sbox_8_T22), .Z0_t (SubBytesIns_Inst_Sbox_8_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T2), .B0_t (SubBytesIns_Inst_Sbox_8_T10), .Z0_t (SubBytesIns_Inst_Sbox_8_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T20), .B0_t (SubBytesIns_Inst_Sbox_8_T17), .Z0_t (SubBytesIns_Inst_Sbox_8_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T3), .B0_t (SubBytesIns_Inst_Sbox_8_T16), .Z0_t (SubBytesIns_Inst_Sbox_8_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T1), .B0_t (SubBytesIns_Inst_Sbox_8_T12), .Z0_t (SubBytesIns_Inst_Sbox_8_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T13), .B0_t (SubBytesIns_Inst_Sbox_8_T6), .Z0_t (SubBytesIns_Inst_Sbox_8_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T23), .B0_t (SubBytesIns_Inst_Sbox_8_T8), .Z0_t (SubBytesIns_Inst_Sbox_8_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T14), .B0_t (SubBytesIns_Inst_Sbox_8_M1), .Z0_t (SubBytesIns_Inst_Sbox_8_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T19), .B0_t (ciphertext[64]), .Z0_t (SubBytesIns_Inst_Sbox_8_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M4), .B0_t (SubBytesIns_Inst_Sbox_8_M1), .Z0_t (SubBytesIns_Inst_Sbox_8_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T3), .B0_t (SubBytesIns_Inst_Sbox_8_T16), .Z0_t (SubBytesIns_Inst_Sbox_8_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T22), .B0_t (SubBytesIns_Inst_Sbox_8_T9), .Z0_t (SubBytesIns_Inst_Sbox_8_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T26), .B0_t (SubBytesIns_Inst_Sbox_8_M6), .Z0_t (SubBytesIns_Inst_Sbox_8_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T20), .B0_t (SubBytesIns_Inst_Sbox_8_T17), .Z0_t (SubBytesIns_Inst_Sbox_8_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M9), .B0_t (SubBytesIns_Inst_Sbox_8_M6), .Z0_t (SubBytesIns_Inst_Sbox_8_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T1), .B0_t (SubBytesIns_Inst_Sbox_8_T15), .Z0_t (SubBytesIns_Inst_Sbox_8_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T4), .B0_t (SubBytesIns_Inst_Sbox_8_T27), .Z0_t (SubBytesIns_Inst_Sbox_8_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M12), .B0_t (SubBytesIns_Inst_Sbox_8_M11), .Z0_t (SubBytesIns_Inst_Sbox_8_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_T2), .B0_t (SubBytesIns_Inst_Sbox_8_T10), .Z0_t (SubBytesIns_Inst_Sbox_8_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M14), .B0_t (SubBytesIns_Inst_Sbox_8_M11), .Z0_t (SubBytesIns_Inst_Sbox_8_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M3), .B0_t (SubBytesIns_Inst_Sbox_8_M2), .Z0_t (SubBytesIns_Inst_Sbox_8_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M5), .B0_t (SubBytesIns_Inst_Sbox_8_T24), .Z0_t (SubBytesIns_Inst_Sbox_8_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M8), .B0_t (SubBytesIns_Inst_Sbox_8_M7), .Z0_t (SubBytesIns_Inst_Sbox_8_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M10), .B0_t (SubBytesIns_Inst_Sbox_8_M15), .Z0_t (SubBytesIns_Inst_Sbox_8_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M16), .B0_t (SubBytesIns_Inst_Sbox_8_M13), .Z0_t (SubBytesIns_Inst_Sbox_8_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M17), .B0_t (SubBytesIns_Inst_Sbox_8_M15), .Z0_t (SubBytesIns_Inst_Sbox_8_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M18), .B0_t (SubBytesIns_Inst_Sbox_8_M13), .Z0_t (SubBytesIns_Inst_Sbox_8_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M19), .B0_t (SubBytesIns_Inst_Sbox_8_T25), .Z0_t (SubBytesIns_Inst_Sbox_8_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M22), .B0_t (SubBytesIns_Inst_Sbox_8_M23), .Z0_t (SubBytesIns_Inst_Sbox_8_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M22), .B0_t (SubBytesIns_Inst_Sbox_8_M20), .Z0_t (SubBytesIns_Inst_Sbox_8_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M21), .B0_t (SubBytesIns_Inst_Sbox_8_M25), .Z0_t (SubBytesIns_Inst_Sbox_8_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M20), .B0_t (SubBytesIns_Inst_Sbox_8_M21), .Z0_t (SubBytesIns_Inst_Sbox_8_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M23), .B0_t (SubBytesIns_Inst_Sbox_8_M25), .Z0_t (SubBytesIns_Inst_Sbox_8_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M28), .B0_t (SubBytesIns_Inst_Sbox_8_M27), .Z0_t (SubBytesIns_Inst_Sbox_8_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M26), .B0_t (SubBytesIns_Inst_Sbox_8_M24), .Z0_t (SubBytesIns_Inst_Sbox_8_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M20), .B0_t (SubBytesIns_Inst_Sbox_8_M23), .Z0_t (SubBytesIns_Inst_Sbox_8_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M27), .B0_t (SubBytesIns_Inst_Sbox_8_M31), .Z0_t (SubBytesIns_Inst_Sbox_8_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M27), .B0_t (SubBytesIns_Inst_Sbox_8_M25), .Z0_t (SubBytesIns_Inst_Sbox_8_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M21), .B0_t (SubBytesIns_Inst_Sbox_8_M22), .Z0_t (SubBytesIns_Inst_Sbox_8_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M24), .B0_t (SubBytesIns_Inst_Sbox_8_M34), .Z0_t (SubBytesIns_Inst_Sbox_8_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M24), .B0_t (SubBytesIns_Inst_Sbox_8_M25), .Z0_t (SubBytesIns_Inst_Sbox_8_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M21), .B0_t (SubBytesIns_Inst_Sbox_8_M29), .Z0_t (SubBytesIns_Inst_Sbox_8_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M32), .B0_t (SubBytesIns_Inst_Sbox_8_M33), .Z0_t (SubBytesIns_Inst_Sbox_8_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M23), .B0_t (SubBytesIns_Inst_Sbox_8_M30), .Z0_t (SubBytesIns_Inst_Sbox_8_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M35), .B0_t (SubBytesIns_Inst_Sbox_8_M36), .Z0_t (SubBytesIns_Inst_Sbox_8_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M38), .B0_t (SubBytesIns_Inst_Sbox_8_M40), .Z0_t (SubBytesIns_Inst_Sbox_8_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M37), .B0_t (SubBytesIns_Inst_Sbox_8_M39), .Z0_t (SubBytesIns_Inst_Sbox_8_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M37), .B0_t (SubBytesIns_Inst_Sbox_8_M38), .Z0_t (SubBytesIns_Inst_Sbox_8_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M39), .B0_t (SubBytesIns_Inst_Sbox_8_M40), .Z0_t (SubBytesIns_Inst_Sbox_8_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M42), .B0_t (SubBytesIns_Inst_Sbox_8_M41), .Z0_t (SubBytesIns_Inst_Sbox_8_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M44), .B0_t (SubBytesIns_Inst_Sbox_8_T6), .Z0_t (SubBytesIns_Inst_Sbox_8_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M40), .B0_t (SubBytesIns_Inst_Sbox_8_T8), .Z0_t (SubBytesIns_Inst_Sbox_8_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M39), .B0_t (ciphertext[64]), .Z0_t (SubBytesIns_Inst_Sbox_8_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M43), .B0_t (SubBytesIns_Inst_Sbox_8_T16), .Z0_t (SubBytesIns_Inst_Sbox_8_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M38), .B0_t (SubBytesIns_Inst_Sbox_8_T9), .Z0_t (SubBytesIns_Inst_Sbox_8_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M37), .B0_t (SubBytesIns_Inst_Sbox_8_T17), .Z0_t (SubBytesIns_Inst_Sbox_8_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M42), .B0_t (SubBytesIns_Inst_Sbox_8_T15), .Z0_t (SubBytesIns_Inst_Sbox_8_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M45), .B0_t (SubBytesIns_Inst_Sbox_8_T27), .Z0_t (SubBytesIns_Inst_Sbox_8_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M41), .B0_t (SubBytesIns_Inst_Sbox_8_T10), .Z0_t (SubBytesIns_Inst_Sbox_8_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M44), .B0_t (SubBytesIns_Inst_Sbox_8_T13), .Z0_t (SubBytesIns_Inst_Sbox_8_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M40), .B0_t (SubBytesIns_Inst_Sbox_8_T23), .Z0_t (SubBytesIns_Inst_Sbox_8_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M39), .B0_t (SubBytesIns_Inst_Sbox_8_T19), .Z0_t (SubBytesIns_Inst_Sbox_8_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M43), .B0_t (SubBytesIns_Inst_Sbox_8_T3), .Z0_t (SubBytesIns_Inst_Sbox_8_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M38), .B0_t (SubBytesIns_Inst_Sbox_8_T22), .Z0_t (SubBytesIns_Inst_Sbox_8_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M37), .B0_t (SubBytesIns_Inst_Sbox_8_T20), .Z0_t (SubBytesIns_Inst_Sbox_8_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M42), .B0_t (SubBytesIns_Inst_Sbox_8_T1), .Z0_t (SubBytesIns_Inst_Sbox_8_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M45), .B0_t (SubBytesIns_Inst_Sbox_8_T4), .Z0_t (SubBytesIns_Inst_Sbox_8_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M41), .B0_t (SubBytesIns_Inst_Sbox_8_T2), .Z0_t (SubBytesIns_Inst_Sbox_8_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M61), .B0_t (SubBytesIns_Inst_Sbox_8_M62), .Z0_t (SubBytesIns_Inst_Sbox_8_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M50), .B0_t (SubBytesIns_Inst_Sbox_8_M56), .Z0_t (SubBytesIns_Inst_Sbox_8_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M46), .B0_t (SubBytesIns_Inst_Sbox_8_M48), .Z0_t (SubBytesIns_Inst_Sbox_8_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M47), .B0_t (SubBytesIns_Inst_Sbox_8_M55), .Z0_t (SubBytesIns_Inst_Sbox_8_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M54), .B0_t (SubBytesIns_Inst_Sbox_8_M58), .Z0_t (SubBytesIns_Inst_Sbox_8_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M49), .B0_t (SubBytesIns_Inst_Sbox_8_M61), .Z0_t (SubBytesIns_Inst_Sbox_8_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M62), .B0_t (SubBytesIns_Inst_Sbox_8_L5), .Z0_t (SubBytesIns_Inst_Sbox_8_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M46), .B0_t (SubBytesIns_Inst_Sbox_8_L3), .Z0_t (SubBytesIns_Inst_Sbox_8_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M51), .B0_t (SubBytesIns_Inst_Sbox_8_M59), .Z0_t (SubBytesIns_Inst_Sbox_8_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M52), .B0_t (SubBytesIns_Inst_Sbox_8_M53), .Z0_t (SubBytesIns_Inst_Sbox_8_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M53), .B0_t (SubBytesIns_Inst_Sbox_8_L4), .Z0_t (SubBytesIns_Inst_Sbox_8_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M60), .B0_t (SubBytesIns_Inst_Sbox_8_L2), .Z0_t (SubBytesIns_Inst_Sbox_8_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M48), .B0_t (SubBytesIns_Inst_Sbox_8_M51), .Z0_t (SubBytesIns_Inst_Sbox_8_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M50), .B0_t (SubBytesIns_Inst_Sbox_8_L0), .Z0_t (SubBytesIns_Inst_Sbox_8_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M52), .B0_t (SubBytesIns_Inst_Sbox_8_M61), .Z0_t (SubBytesIns_Inst_Sbox_8_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M55), .B0_t (SubBytesIns_Inst_Sbox_8_L1), .Z0_t (SubBytesIns_Inst_Sbox_8_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M56), .B0_t (SubBytesIns_Inst_Sbox_8_L0), .Z0_t (SubBytesIns_Inst_Sbox_8_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M57), .B0_t (SubBytesIns_Inst_Sbox_8_L1), .Z0_t (SubBytesIns_Inst_Sbox_8_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M58), .B0_t (SubBytesIns_Inst_Sbox_8_L8), .Z0_t (SubBytesIns_Inst_Sbox_8_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_M63), .B0_t (SubBytesIns_Inst_Sbox_8_L4), .Z0_t (SubBytesIns_Inst_Sbox_8_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L0), .B0_t (SubBytesIns_Inst_Sbox_8_L1), .Z0_t (SubBytesIns_Inst_Sbox_8_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L1), .B0_t (SubBytesIns_Inst_Sbox_8_L7), .Z0_t (SubBytesIns_Inst_Sbox_8_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L3), .B0_t (SubBytesIns_Inst_Sbox_8_L12), .Z0_t (SubBytesIns_Inst_Sbox_8_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L18), .B0_t (SubBytesIns_Inst_Sbox_8_L2), .Z0_t (SubBytesIns_Inst_Sbox_8_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L15), .B0_t (SubBytesIns_Inst_Sbox_8_L9), .Z0_t (SubBytesIns_Inst_Sbox_8_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L6), .B0_t (SubBytesIns_Inst_Sbox_8_L10), .Z0_t (SubBytesIns_Inst_Sbox_8_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L7), .B0_t (SubBytesIns_Inst_Sbox_8_L9), .Z0_t (SubBytesIns_Inst_Sbox_8_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L8), .B0_t (SubBytesIns_Inst_Sbox_8_L10), .Z0_t (SubBytesIns_Inst_Sbox_8_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L11), .B0_t (SubBytesIns_Inst_Sbox_8_L14), .Z0_t (SubBytesIns_Inst_Sbox_8_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L11), .B0_t (SubBytesIns_Inst_Sbox_8_L17), .Z0_t (SubBytesIns_Inst_Sbox_8_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L6), .B0_t (SubBytesIns_Inst_Sbox_8_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L16), .B0_t (SubBytesIns_Inst_Sbox_8_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L19), .B0_t (SubBytesIns_Inst_Sbox_8_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L6), .B0_t (SubBytesIns_Inst_Sbox_8_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L20), .B0_t (SubBytesIns_Inst_Sbox_8_L22), .Z0_t (MixColumnsInput[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L25), .B0_t (SubBytesIns_Inst_Sbox_8_L29), .Z0_t (MixColumnsInput[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L13), .B0_t (SubBytesIns_Inst_Sbox_8_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_8_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_8_L6), .B0_t (SubBytesIns_Inst_Sbox_8_L23), .Z0_t (MixColumnsInput[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T1_U1 ( .A0_t (ciphertext[79]), .B0_t (ciphertext[76]), .Z0_t (SubBytesIns_Inst_Sbox_9_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T2_U1 ( .A0_t (ciphertext[79]), .B0_t (ciphertext[74]), .Z0_t (SubBytesIns_Inst_Sbox_9_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T3_U1 ( .A0_t (ciphertext[79]), .B0_t (ciphertext[73]), .Z0_t (SubBytesIns_Inst_Sbox_9_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T4_U1 ( .A0_t (ciphertext[76]), .B0_t (ciphertext[74]), .Z0_t (SubBytesIns_Inst_Sbox_9_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T5_U1 ( .A0_t (ciphertext[75]), .B0_t (ciphertext[73]), .Z0_t (SubBytesIns_Inst_Sbox_9_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T1), .B0_t (SubBytesIns_Inst_Sbox_9_T5), .Z0_t (SubBytesIns_Inst_Sbox_9_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T7_U1 ( .A0_t (ciphertext[78]), .B0_t (ciphertext[77]), .Z0_t (SubBytesIns_Inst_Sbox_9_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T8_U1 ( .A0_t (ciphertext[72]), .B0_t (SubBytesIns_Inst_Sbox_9_T6), .Z0_t (SubBytesIns_Inst_Sbox_9_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T9_U1 ( .A0_t (ciphertext[72]), .B0_t (SubBytesIns_Inst_Sbox_9_T7), .Z0_t (SubBytesIns_Inst_Sbox_9_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T6), .B0_t (SubBytesIns_Inst_Sbox_9_T7), .Z0_t (SubBytesIns_Inst_Sbox_9_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T11_U1 ( .A0_t (ciphertext[78]), .B0_t (ciphertext[74]), .Z0_t (SubBytesIns_Inst_Sbox_9_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T12_U1 ( .A0_t (ciphertext[77]), .B0_t (ciphertext[74]), .Z0_t (SubBytesIns_Inst_Sbox_9_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T3), .B0_t (SubBytesIns_Inst_Sbox_9_T4), .Z0_t (SubBytesIns_Inst_Sbox_9_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T6), .B0_t (SubBytesIns_Inst_Sbox_9_T11), .Z0_t (SubBytesIns_Inst_Sbox_9_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T5), .B0_t (SubBytesIns_Inst_Sbox_9_T11), .Z0_t (SubBytesIns_Inst_Sbox_9_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T5), .B0_t (SubBytesIns_Inst_Sbox_9_T12), .Z0_t (SubBytesIns_Inst_Sbox_9_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T9), .B0_t (SubBytesIns_Inst_Sbox_9_T16), .Z0_t (SubBytesIns_Inst_Sbox_9_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T18_U1 ( .A0_t (ciphertext[76]), .B0_t (ciphertext[72]), .Z0_t (SubBytesIns_Inst_Sbox_9_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T7), .B0_t (SubBytesIns_Inst_Sbox_9_T18), .Z0_t (SubBytesIns_Inst_Sbox_9_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T1), .B0_t (SubBytesIns_Inst_Sbox_9_T19), .Z0_t (SubBytesIns_Inst_Sbox_9_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T21_U1 ( .A0_t (ciphertext[73]), .B0_t (ciphertext[72]), .Z0_t (SubBytesIns_Inst_Sbox_9_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T7), .B0_t (SubBytesIns_Inst_Sbox_9_T21), .Z0_t (SubBytesIns_Inst_Sbox_9_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T2), .B0_t (SubBytesIns_Inst_Sbox_9_T22), .Z0_t (SubBytesIns_Inst_Sbox_9_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T2), .B0_t (SubBytesIns_Inst_Sbox_9_T10), .Z0_t (SubBytesIns_Inst_Sbox_9_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T20), .B0_t (SubBytesIns_Inst_Sbox_9_T17), .Z0_t (SubBytesIns_Inst_Sbox_9_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T3), .B0_t (SubBytesIns_Inst_Sbox_9_T16), .Z0_t (SubBytesIns_Inst_Sbox_9_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T1), .B0_t (SubBytesIns_Inst_Sbox_9_T12), .Z0_t (SubBytesIns_Inst_Sbox_9_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T13), .B0_t (SubBytesIns_Inst_Sbox_9_T6), .Z0_t (SubBytesIns_Inst_Sbox_9_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T23), .B0_t (SubBytesIns_Inst_Sbox_9_T8), .Z0_t (SubBytesIns_Inst_Sbox_9_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T14), .B0_t (SubBytesIns_Inst_Sbox_9_M1), .Z0_t (SubBytesIns_Inst_Sbox_9_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T19), .B0_t (ciphertext[72]), .Z0_t (SubBytesIns_Inst_Sbox_9_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M4), .B0_t (SubBytesIns_Inst_Sbox_9_M1), .Z0_t (SubBytesIns_Inst_Sbox_9_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T3), .B0_t (SubBytesIns_Inst_Sbox_9_T16), .Z0_t (SubBytesIns_Inst_Sbox_9_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T22), .B0_t (SubBytesIns_Inst_Sbox_9_T9), .Z0_t (SubBytesIns_Inst_Sbox_9_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T26), .B0_t (SubBytesIns_Inst_Sbox_9_M6), .Z0_t (SubBytesIns_Inst_Sbox_9_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T20), .B0_t (SubBytesIns_Inst_Sbox_9_T17), .Z0_t (SubBytesIns_Inst_Sbox_9_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M9), .B0_t (SubBytesIns_Inst_Sbox_9_M6), .Z0_t (SubBytesIns_Inst_Sbox_9_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T1), .B0_t (SubBytesIns_Inst_Sbox_9_T15), .Z0_t (SubBytesIns_Inst_Sbox_9_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T4), .B0_t (SubBytesIns_Inst_Sbox_9_T27), .Z0_t (SubBytesIns_Inst_Sbox_9_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M12), .B0_t (SubBytesIns_Inst_Sbox_9_M11), .Z0_t (SubBytesIns_Inst_Sbox_9_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_T2), .B0_t (SubBytesIns_Inst_Sbox_9_T10), .Z0_t (SubBytesIns_Inst_Sbox_9_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M14), .B0_t (SubBytesIns_Inst_Sbox_9_M11), .Z0_t (SubBytesIns_Inst_Sbox_9_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M3), .B0_t (SubBytesIns_Inst_Sbox_9_M2), .Z0_t (SubBytesIns_Inst_Sbox_9_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M5), .B0_t (SubBytesIns_Inst_Sbox_9_T24), .Z0_t (SubBytesIns_Inst_Sbox_9_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M8), .B0_t (SubBytesIns_Inst_Sbox_9_M7), .Z0_t (SubBytesIns_Inst_Sbox_9_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M10), .B0_t (SubBytesIns_Inst_Sbox_9_M15), .Z0_t (SubBytesIns_Inst_Sbox_9_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M16), .B0_t (SubBytesIns_Inst_Sbox_9_M13), .Z0_t (SubBytesIns_Inst_Sbox_9_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M17), .B0_t (SubBytesIns_Inst_Sbox_9_M15), .Z0_t (SubBytesIns_Inst_Sbox_9_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M18), .B0_t (SubBytesIns_Inst_Sbox_9_M13), .Z0_t (SubBytesIns_Inst_Sbox_9_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M19), .B0_t (SubBytesIns_Inst_Sbox_9_T25), .Z0_t (SubBytesIns_Inst_Sbox_9_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M22), .B0_t (SubBytesIns_Inst_Sbox_9_M23), .Z0_t (SubBytesIns_Inst_Sbox_9_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M22), .B0_t (SubBytesIns_Inst_Sbox_9_M20), .Z0_t (SubBytesIns_Inst_Sbox_9_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M21), .B0_t (SubBytesIns_Inst_Sbox_9_M25), .Z0_t (SubBytesIns_Inst_Sbox_9_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M20), .B0_t (SubBytesIns_Inst_Sbox_9_M21), .Z0_t (SubBytesIns_Inst_Sbox_9_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M23), .B0_t (SubBytesIns_Inst_Sbox_9_M25), .Z0_t (SubBytesIns_Inst_Sbox_9_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M28), .B0_t (SubBytesIns_Inst_Sbox_9_M27), .Z0_t (SubBytesIns_Inst_Sbox_9_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M26), .B0_t (SubBytesIns_Inst_Sbox_9_M24), .Z0_t (SubBytesIns_Inst_Sbox_9_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M20), .B0_t (SubBytesIns_Inst_Sbox_9_M23), .Z0_t (SubBytesIns_Inst_Sbox_9_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M27), .B0_t (SubBytesIns_Inst_Sbox_9_M31), .Z0_t (SubBytesIns_Inst_Sbox_9_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M27), .B0_t (SubBytesIns_Inst_Sbox_9_M25), .Z0_t (SubBytesIns_Inst_Sbox_9_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M21), .B0_t (SubBytesIns_Inst_Sbox_9_M22), .Z0_t (SubBytesIns_Inst_Sbox_9_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M24), .B0_t (SubBytesIns_Inst_Sbox_9_M34), .Z0_t (SubBytesIns_Inst_Sbox_9_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M24), .B0_t (SubBytesIns_Inst_Sbox_9_M25), .Z0_t (SubBytesIns_Inst_Sbox_9_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M21), .B0_t (SubBytesIns_Inst_Sbox_9_M29), .Z0_t (SubBytesIns_Inst_Sbox_9_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M32), .B0_t (SubBytesIns_Inst_Sbox_9_M33), .Z0_t (SubBytesIns_Inst_Sbox_9_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M23), .B0_t (SubBytesIns_Inst_Sbox_9_M30), .Z0_t (SubBytesIns_Inst_Sbox_9_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M35), .B0_t (SubBytesIns_Inst_Sbox_9_M36), .Z0_t (SubBytesIns_Inst_Sbox_9_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M38), .B0_t (SubBytesIns_Inst_Sbox_9_M40), .Z0_t (SubBytesIns_Inst_Sbox_9_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M37), .B0_t (SubBytesIns_Inst_Sbox_9_M39), .Z0_t (SubBytesIns_Inst_Sbox_9_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M37), .B0_t (SubBytesIns_Inst_Sbox_9_M38), .Z0_t (SubBytesIns_Inst_Sbox_9_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M39), .B0_t (SubBytesIns_Inst_Sbox_9_M40), .Z0_t (SubBytesIns_Inst_Sbox_9_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M42), .B0_t (SubBytesIns_Inst_Sbox_9_M41), .Z0_t (SubBytesIns_Inst_Sbox_9_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M44), .B0_t (SubBytesIns_Inst_Sbox_9_T6), .Z0_t (SubBytesIns_Inst_Sbox_9_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M40), .B0_t (SubBytesIns_Inst_Sbox_9_T8), .Z0_t (SubBytesIns_Inst_Sbox_9_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M39), .B0_t (ciphertext[72]), .Z0_t (SubBytesIns_Inst_Sbox_9_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M43), .B0_t (SubBytesIns_Inst_Sbox_9_T16), .Z0_t (SubBytesIns_Inst_Sbox_9_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M38), .B0_t (SubBytesIns_Inst_Sbox_9_T9), .Z0_t (SubBytesIns_Inst_Sbox_9_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M37), .B0_t (SubBytesIns_Inst_Sbox_9_T17), .Z0_t (SubBytesIns_Inst_Sbox_9_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M42), .B0_t (SubBytesIns_Inst_Sbox_9_T15), .Z0_t (SubBytesIns_Inst_Sbox_9_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M45), .B0_t (SubBytesIns_Inst_Sbox_9_T27), .Z0_t (SubBytesIns_Inst_Sbox_9_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M41), .B0_t (SubBytesIns_Inst_Sbox_9_T10), .Z0_t (SubBytesIns_Inst_Sbox_9_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M44), .B0_t (SubBytesIns_Inst_Sbox_9_T13), .Z0_t (SubBytesIns_Inst_Sbox_9_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M40), .B0_t (SubBytesIns_Inst_Sbox_9_T23), .Z0_t (SubBytesIns_Inst_Sbox_9_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M39), .B0_t (SubBytesIns_Inst_Sbox_9_T19), .Z0_t (SubBytesIns_Inst_Sbox_9_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M43), .B0_t (SubBytesIns_Inst_Sbox_9_T3), .Z0_t (SubBytesIns_Inst_Sbox_9_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M38), .B0_t (SubBytesIns_Inst_Sbox_9_T22), .Z0_t (SubBytesIns_Inst_Sbox_9_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M37), .B0_t (SubBytesIns_Inst_Sbox_9_T20), .Z0_t (SubBytesIns_Inst_Sbox_9_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M42), .B0_t (SubBytesIns_Inst_Sbox_9_T1), .Z0_t (SubBytesIns_Inst_Sbox_9_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M45), .B0_t (SubBytesIns_Inst_Sbox_9_T4), .Z0_t (SubBytesIns_Inst_Sbox_9_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M41), .B0_t (SubBytesIns_Inst_Sbox_9_T2), .Z0_t (SubBytesIns_Inst_Sbox_9_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M61), .B0_t (SubBytesIns_Inst_Sbox_9_M62), .Z0_t (SubBytesIns_Inst_Sbox_9_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M50), .B0_t (SubBytesIns_Inst_Sbox_9_M56), .Z0_t (SubBytesIns_Inst_Sbox_9_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M46), .B0_t (SubBytesIns_Inst_Sbox_9_M48), .Z0_t (SubBytesIns_Inst_Sbox_9_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M47), .B0_t (SubBytesIns_Inst_Sbox_9_M55), .Z0_t (SubBytesIns_Inst_Sbox_9_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M54), .B0_t (SubBytesIns_Inst_Sbox_9_M58), .Z0_t (SubBytesIns_Inst_Sbox_9_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M49), .B0_t (SubBytesIns_Inst_Sbox_9_M61), .Z0_t (SubBytesIns_Inst_Sbox_9_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M62), .B0_t (SubBytesIns_Inst_Sbox_9_L5), .Z0_t (SubBytesIns_Inst_Sbox_9_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M46), .B0_t (SubBytesIns_Inst_Sbox_9_L3), .Z0_t (SubBytesIns_Inst_Sbox_9_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M51), .B0_t (SubBytesIns_Inst_Sbox_9_M59), .Z0_t (SubBytesIns_Inst_Sbox_9_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M52), .B0_t (SubBytesIns_Inst_Sbox_9_M53), .Z0_t (SubBytesIns_Inst_Sbox_9_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M53), .B0_t (SubBytesIns_Inst_Sbox_9_L4), .Z0_t (SubBytesIns_Inst_Sbox_9_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M60), .B0_t (SubBytesIns_Inst_Sbox_9_L2), .Z0_t (SubBytesIns_Inst_Sbox_9_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M48), .B0_t (SubBytesIns_Inst_Sbox_9_M51), .Z0_t (SubBytesIns_Inst_Sbox_9_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M50), .B0_t (SubBytesIns_Inst_Sbox_9_L0), .Z0_t (SubBytesIns_Inst_Sbox_9_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M52), .B0_t (SubBytesIns_Inst_Sbox_9_M61), .Z0_t (SubBytesIns_Inst_Sbox_9_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M55), .B0_t (SubBytesIns_Inst_Sbox_9_L1), .Z0_t (SubBytesIns_Inst_Sbox_9_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M56), .B0_t (SubBytesIns_Inst_Sbox_9_L0), .Z0_t (SubBytesIns_Inst_Sbox_9_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M57), .B0_t (SubBytesIns_Inst_Sbox_9_L1), .Z0_t (SubBytesIns_Inst_Sbox_9_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M58), .B0_t (SubBytesIns_Inst_Sbox_9_L8), .Z0_t (SubBytesIns_Inst_Sbox_9_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_M63), .B0_t (SubBytesIns_Inst_Sbox_9_L4), .Z0_t (SubBytesIns_Inst_Sbox_9_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L0), .B0_t (SubBytesIns_Inst_Sbox_9_L1), .Z0_t (SubBytesIns_Inst_Sbox_9_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L1), .B0_t (SubBytesIns_Inst_Sbox_9_L7), .Z0_t (SubBytesIns_Inst_Sbox_9_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L3), .B0_t (SubBytesIns_Inst_Sbox_9_L12), .Z0_t (SubBytesIns_Inst_Sbox_9_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L18), .B0_t (SubBytesIns_Inst_Sbox_9_L2), .Z0_t (SubBytesIns_Inst_Sbox_9_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L15), .B0_t (SubBytesIns_Inst_Sbox_9_L9), .Z0_t (SubBytesIns_Inst_Sbox_9_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L6), .B0_t (SubBytesIns_Inst_Sbox_9_L10), .Z0_t (SubBytesIns_Inst_Sbox_9_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L7), .B0_t (SubBytesIns_Inst_Sbox_9_L9), .Z0_t (SubBytesIns_Inst_Sbox_9_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L8), .B0_t (SubBytesIns_Inst_Sbox_9_L10), .Z0_t (SubBytesIns_Inst_Sbox_9_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L11), .B0_t (SubBytesIns_Inst_Sbox_9_L14), .Z0_t (SubBytesIns_Inst_Sbox_9_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L11), .B0_t (SubBytesIns_Inst_Sbox_9_L17), .Z0_t (SubBytesIns_Inst_Sbox_9_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L6), .B0_t (SubBytesIns_Inst_Sbox_9_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L16), .B0_t (SubBytesIns_Inst_Sbox_9_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L19), .B0_t (SubBytesIns_Inst_Sbox_9_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L6), .B0_t (SubBytesIns_Inst_Sbox_9_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L20), .B0_t (SubBytesIns_Inst_Sbox_9_L22), .Z0_t (MixColumnsInput[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L25), .B0_t (SubBytesIns_Inst_Sbox_9_L29), .Z0_t (MixColumnsInput[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L13), .B0_t (SubBytesIns_Inst_Sbox_9_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_9_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_9_L6), .B0_t (SubBytesIns_Inst_Sbox_9_L23), .Z0_t (MixColumnsInput[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T1_U1 ( .A0_t (ciphertext[87]), .B0_t (ciphertext[84]), .Z0_t (SubBytesIns_Inst_Sbox_10_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T2_U1 ( .A0_t (ciphertext[87]), .B0_t (ciphertext[82]), .Z0_t (SubBytesIns_Inst_Sbox_10_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T3_U1 ( .A0_t (ciphertext[87]), .B0_t (ciphertext[81]), .Z0_t (SubBytesIns_Inst_Sbox_10_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T4_U1 ( .A0_t (ciphertext[84]), .B0_t (ciphertext[82]), .Z0_t (SubBytesIns_Inst_Sbox_10_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T5_U1 ( .A0_t (ciphertext[83]), .B0_t (ciphertext[81]), .Z0_t (SubBytesIns_Inst_Sbox_10_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T1), .B0_t (SubBytesIns_Inst_Sbox_10_T5), .Z0_t (SubBytesIns_Inst_Sbox_10_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T7_U1 ( .A0_t (ciphertext[86]), .B0_t (ciphertext[85]), .Z0_t (SubBytesIns_Inst_Sbox_10_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T8_U1 ( .A0_t (ciphertext[80]), .B0_t (SubBytesIns_Inst_Sbox_10_T6), .Z0_t (SubBytesIns_Inst_Sbox_10_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T9_U1 ( .A0_t (ciphertext[80]), .B0_t (SubBytesIns_Inst_Sbox_10_T7), .Z0_t (SubBytesIns_Inst_Sbox_10_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T6), .B0_t (SubBytesIns_Inst_Sbox_10_T7), .Z0_t (SubBytesIns_Inst_Sbox_10_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T11_U1 ( .A0_t (ciphertext[86]), .B0_t (ciphertext[82]), .Z0_t (SubBytesIns_Inst_Sbox_10_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T12_U1 ( .A0_t (ciphertext[85]), .B0_t (ciphertext[82]), .Z0_t (SubBytesIns_Inst_Sbox_10_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T3), .B0_t (SubBytesIns_Inst_Sbox_10_T4), .Z0_t (SubBytesIns_Inst_Sbox_10_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T6), .B0_t (SubBytesIns_Inst_Sbox_10_T11), .Z0_t (SubBytesIns_Inst_Sbox_10_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T5), .B0_t (SubBytesIns_Inst_Sbox_10_T11), .Z0_t (SubBytesIns_Inst_Sbox_10_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T5), .B0_t (SubBytesIns_Inst_Sbox_10_T12), .Z0_t (SubBytesIns_Inst_Sbox_10_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T9), .B0_t (SubBytesIns_Inst_Sbox_10_T16), .Z0_t (SubBytesIns_Inst_Sbox_10_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T18_U1 ( .A0_t (ciphertext[84]), .B0_t (ciphertext[80]), .Z0_t (SubBytesIns_Inst_Sbox_10_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T7), .B0_t (SubBytesIns_Inst_Sbox_10_T18), .Z0_t (SubBytesIns_Inst_Sbox_10_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T1), .B0_t (SubBytesIns_Inst_Sbox_10_T19), .Z0_t (SubBytesIns_Inst_Sbox_10_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T21_U1 ( .A0_t (ciphertext[81]), .B0_t (ciphertext[80]), .Z0_t (SubBytesIns_Inst_Sbox_10_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T7), .B0_t (SubBytesIns_Inst_Sbox_10_T21), .Z0_t (SubBytesIns_Inst_Sbox_10_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T2), .B0_t (SubBytesIns_Inst_Sbox_10_T22), .Z0_t (SubBytesIns_Inst_Sbox_10_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T2), .B0_t (SubBytesIns_Inst_Sbox_10_T10), .Z0_t (SubBytesIns_Inst_Sbox_10_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T20), .B0_t (SubBytesIns_Inst_Sbox_10_T17), .Z0_t (SubBytesIns_Inst_Sbox_10_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T3), .B0_t (SubBytesIns_Inst_Sbox_10_T16), .Z0_t (SubBytesIns_Inst_Sbox_10_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T1), .B0_t (SubBytesIns_Inst_Sbox_10_T12), .Z0_t (SubBytesIns_Inst_Sbox_10_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T13), .B0_t (SubBytesIns_Inst_Sbox_10_T6), .Z0_t (SubBytesIns_Inst_Sbox_10_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T23), .B0_t (SubBytesIns_Inst_Sbox_10_T8), .Z0_t (SubBytesIns_Inst_Sbox_10_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T14), .B0_t (SubBytesIns_Inst_Sbox_10_M1), .Z0_t (SubBytesIns_Inst_Sbox_10_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T19), .B0_t (ciphertext[80]), .Z0_t (SubBytesIns_Inst_Sbox_10_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M4), .B0_t (SubBytesIns_Inst_Sbox_10_M1), .Z0_t (SubBytesIns_Inst_Sbox_10_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T3), .B0_t (SubBytesIns_Inst_Sbox_10_T16), .Z0_t (SubBytesIns_Inst_Sbox_10_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T22), .B0_t (SubBytesIns_Inst_Sbox_10_T9), .Z0_t (SubBytesIns_Inst_Sbox_10_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T26), .B0_t (SubBytesIns_Inst_Sbox_10_M6), .Z0_t (SubBytesIns_Inst_Sbox_10_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T20), .B0_t (SubBytesIns_Inst_Sbox_10_T17), .Z0_t (SubBytesIns_Inst_Sbox_10_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M9), .B0_t (SubBytesIns_Inst_Sbox_10_M6), .Z0_t (SubBytesIns_Inst_Sbox_10_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T1), .B0_t (SubBytesIns_Inst_Sbox_10_T15), .Z0_t (SubBytesIns_Inst_Sbox_10_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T4), .B0_t (SubBytesIns_Inst_Sbox_10_T27), .Z0_t (SubBytesIns_Inst_Sbox_10_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M12), .B0_t (SubBytesIns_Inst_Sbox_10_M11), .Z0_t (SubBytesIns_Inst_Sbox_10_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_T2), .B0_t (SubBytesIns_Inst_Sbox_10_T10), .Z0_t (SubBytesIns_Inst_Sbox_10_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M14), .B0_t (SubBytesIns_Inst_Sbox_10_M11), .Z0_t (SubBytesIns_Inst_Sbox_10_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M3), .B0_t (SubBytesIns_Inst_Sbox_10_M2), .Z0_t (SubBytesIns_Inst_Sbox_10_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M5), .B0_t (SubBytesIns_Inst_Sbox_10_T24), .Z0_t (SubBytesIns_Inst_Sbox_10_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M8), .B0_t (SubBytesIns_Inst_Sbox_10_M7), .Z0_t (SubBytesIns_Inst_Sbox_10_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M10), .B0_t (SubBytesIns_Inst_Sbox_10_M15), .Z0_t (SubBytesIns_Inst_Sbox_10_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M16), .B0_t (SubBytesIns_Inst_Sbox_10_M13), .Z0_t (SubBytesIns_Inst_Sbox_10_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M17), .B0_t (SubBytesIns_Inst_Sbox_10_M15), .Z0_t (SubBytesIns_Inst_Sbox_10_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M18), .B0_t (SubBytesIns_Inst_Sbox_10_M13), .Z0_t (SubBytesIns_Inst_Sbox_10_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M19), .B0_t (SubBytesIns_Inst_Sbox_10_T25), .Z0_t (SubBytesIns_Inst_Sbox_10_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M22), .B0_t (SubBytesIns_Inst_Sbox_10_M23), .Z0_t (SubBytesIns_Inst_Sbox_10_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M22), .B0_t (SubBytesIns_Inst_Sbox_10_M20), .Z0_t (SubBytesIns_Inst_Sbox_10_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M21), .B0_t (SubBytesIns_Inst_Sbox_10_M25), .Z0_t (SubBytesIns_Inst_Sbox_10_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M20), .B0_t (SubBytesIns_Inst_Sbox_10_M21), .Z0_t (SubBytesIns_Inst_Sbox_10_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M23), .B0_t (SubBytesIns_Inst_Sbox_10_M25), .Z0_t (SubBytesIns_Inst_Sbox_10_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M28), .B0_t (SubBytesIns_Inst_Sbox_10_M27), .Z0_t (SubBytesIns_Inst_Sbox_10_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M26), .B0_t (SubBytesIns_Inst_Sbox_10_M24), .Z0_t (SubBytesIns_Inst_Sbox_10_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M20), .B0_t (SubBytesIns_Inst_Sbox_10_M23), .Z0_t (SubBytesIns_Inst_Sbox_10_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M27), .B0_t (SubBytesIns_Inst_Sbox_10_M31), .Z0_t (SubBytesIns_Inst_Sbox_10_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M27), .B0_t (SubBytesIns_Inst_Sbox_10_M25), .Z0_t (SubBytesIns_Inst_Sbox_10_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M21), .B0_t (SubBytesIns_Inst_Sbox_10_M22), .Z0_t (SubBytesIns_Inst_Sbox_10_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M24), .B0_t (SubBytesIns_Inst_Sbox_10_M34), .Z0_t (SubBytesIns_Inst_Sbox_10_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M24), .B0_t (SubBytesIns_Inst_Sbox_10_M25), .Z0_t (SubBytesIns_Inst_Sbox_10_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M21), .B0_t (SubBytesIns_Inst_Sbox_10_M29), .Z0_t (SubBytesIns_Inst_Sbox_10_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M32), .B0_t (SubBytesIns_Inst_Sbox_10_M33), .Z0_t (SubBytesIns_Inst_Sbox_10_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M23), .B0_t (SubBytesIns_Inst_Sbox_10_M30), .Z0_t (SubBytesIns_Inst_Sbox_10_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M35), .B0_t (SubBytesIns_Inst_Sbox_10_M36), .Z0_t (SubBytesIns_Inst_Sbox_10_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M38), .B0_t (SubBytesIns_Inst_Sbox_10_M40), .Z0_t (SubBytesIns_Inst_Sbox_10_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M37), .B0_t (SubBytesIns_Inst_Sbox_10_M39), .Z0_t (SubBytesIns_Inst_Sbox_10_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M37), .B0_t (SubBytesIns_Inst_Sbox_10_M38), .Z0_t (SubBytesIns_Inst_Sbox_10_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M39), .B0_t (SubBytesIns_Inst_Sbox_10_M40), .Z0_t (SubBytesIns_Inst_Sbox_10_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M42), .B0_t (SubBytesIns_Inst_Sbox_10_M41), .Z0_t (SubBytesIns_Inst_Sbox_10_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M44), .B0_t (SubBytesIns_Inst_Sbox_10_T6), .Z0_t (SubBytesIns_Inst_Sbox_10_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M40), .B0_t (SubBytesIns_Inst_Sbox_10_T8), .Z0_t (SubBytesIns_Inst_Sbox_10_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M39), .B0_t (ciphertext[80]), .Z0_t (SubBytesIns_Inst_Sbox_10_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M43), .B0_t (SubBytesIns_Inst_Sbox_10_T16), .Z0_t (SubBytesIns_Inst_Sbox_10_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M38), .B0_t (SubBytesIns_Inst_Sbox_10_T9), .Z0_t (SubBytesIns_Inst_Sbox_10_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M37), .B0_t (SubBytesIns_Inst_Sbox_10_T17), .Z0_t (SubBytesIns_Inst_Sbox_10_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M42), .B0_t (SubBytesIns_Inst_Sbox_10_T15), .Z0_t (SubBytesIns_Inst_Sbox_10_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M45), .B0_t (SubBytesIns_Inst_Sbox_10_T27), .Z0_t (SubBytesIns_Inst_Sbox_10_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M41), .B0_t (SubBytesIns_Inst_Sbox_10_T10), .Z0_t (SubBytesIns_Inst_Sbox_10_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M44), .B0_t (SubBytesIns_Inst_Sbox_10_T13), .Z0_t (SubBytesIns_Inst_Sbox_10_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M40), .B0_t (SubBytesIns_Inst_Sbox_10_T23), .Z0_t (SubBytesIns_Inst_Sbox_10_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M39), .B0_t (SubBytesIns_Inst_Sbox_10_T19), .Z0_t (SubBytesIns_Inst_Sbox_10_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M43), .B0_t (SubBytesIns_Inst_Sbox_10_T3), .Z0_t (SubBytesIns_Inst_Sbox_10_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M38), .B0_t (SubBytesIns_Inst_Sbox_10_T22), .Z0_t (SubBytesIns_Inst_Sbox_10_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M37), .B0_t (SubBytesIns_Inst_Sbox_10_T20), .Z0_t (SubBytesIns_Inst_Sbox_10_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M42), .B0_t (SubBytesIns_Inst_Sbox_10_T1), .Z0_t (SubBytesIns_Inst_Sbox_10_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M45), .B0_t (SubBytesIns_Inst_Sbox_10_T4), .Z0_t (SubBytesIns_Inst_Sbox_10_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M41), .B0_t (SubBytesIns_Inst_Sbox_10_T2), .Z0_t (SubBytesIns_Inst_Sbox_10_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M61), .B0_t (SubBytesIns_Inst_Sbox_10_M62), .Z0_t (SubBytesIns_Inst_Sbox_10_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M50), .B0_t (SubBytesIns_Inst_Sbox_10_M56), .Z0_t (SubBytesIns_Inst_Sbox_10_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M46), .B0_t (SubBytesIns_Inst_Sbox_10_M48), .Z0_t (SubBytesIns_Inst_Sbox_10_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M47), .B0_t (SubBytesIns_Inst_Sbox_10_M55), .Z0_t (SubBytesIns_Inst_Sbox_10_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M54), .B0_t (SubBytesIns_Inst_Sbox_10_M58), .Z0_t (SubBytesIns_Inst_Sbox_10_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M49), .B0_t (SubBytesIns_Inst_Sbox_10_M61), .Z0_t (SubBytesIns_Inst_Sbox_10_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M62), .B0_t (SubBytesIns_Inst_Sbox_10_L5), .Z0_t (SubBytesIns_Inst_Sbox_10_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M46), .B0_t (SubBytesIns_Inst_Sbox_10_L3), .Z0_t (SubBytesIns_Inst_Sbox_10_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M51), .B0_t (SubBytesIns_Inst_Sbox_10_M59), .Z0_t (SubBytesIns_Inst_Sbox_10_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M52), .B0_t (SubBytesIns_Inst_Sbox_10_M53), .Z0_t (SubBytesIns_Inst_Sbox_10_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M53), .B0_t (SubBytesIns_Inst_Sbox_10_L4), .Z0_t (SubBytesIns_Inst_Sbox_10_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M60), .B0_t (SubBytesIns_Inst_Sbox_10_L2), .Z0_t (SubBytesIns_Inst_Sbox_10_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M48), .B0_t (SubBytesIns_Inst_Sbox_10_M51), .Z0_t (SubBytesIns_Inst_Sbox_10_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M50), .B0_t (SubBytesIns_Inst_Sbox_10_L0), .Z0_t (SubBytesIns_Inst_Sbox_10_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M52), .B0_t (SubBytesIns_Inst_Sbox_10_M61), .Z0_t (SubBytesIns_Inst_Sbox_10_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M55), .B0_t (SubBytesIns_Inst_Sbox_10_L1), .Z0_t (SubBytesIns_Inst_Sbox_10_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M56), .B0_t (SubBytesIns_Inst_Sbox_10_L0), .Z0_t (SubBytesIns_Inst_Sbox_10_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M57), .B0_t (SubBytesIns_Inst_Sbox_10_L1), .Z0_t (SubBytesIns_Inst_Sbox_10_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M58), .B0_t (SubBytesIns_Inst_Sbox_10_L8), .Z0_t (SubBytesIns_Inst_Sbox_10_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_M63), .B0_t (SubBytesIns_Inst_Sbox_10_L4), .Z0_t (SubBytesIns_Inst_Sbox_10_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L0), .B0_t (SubBytesIns_Inst_Sbox_10_L1), .Z0_t (SubBytesIns_Inst_Sbox_10_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L1), .B0_t (SubBytesIns_Inst_Sbox_10_L7), .Z0_t (SubBytesIns_Inst_Sbox_10_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L3), .B0_t (SubBytesIns_Inst_Sbox_10_L12), .Z0_t (SubBytesIns_Inst_Sbox_10_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L18), .B0_t (SubBytesIns_Inst_Sbox_10_L2), .Z0_t (SubBytesIns_Inst_Sbox_10_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L15), .B0_t (SubBytesIns_Inst_Sbox_10_L9), .Z0_t (SubBytesIns_Inst_Sbox_10_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L6), .B0_t (SubBytesIns_Inst_Sbox_10_L10), .Z0_t (SubBytesIns_Inst_Sbox_10_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L7), .B0_t (SubBytesIns_Inst_Sbox_10_L9), .Z0_t (SubBytesIns_Inst_Sbox_10_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L8), .B0_t (SubBytesIns_Inst_Sbox_10_L10), .Z0_t (SubBytesIns_Inst_Sbox_10_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L11), .B0_t (SubBytesIns_Inst_Sbox_10_L14), .Z0_t (SubBytesIns_Inst_Sbox_10_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L11), .B0_t (SubBytesIns_Inst_Sbox_10_L17), .Z0_t (SubBytesIns_Inst_Sbox_10_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L6), .B0_t (SubBytesIns_Inst_Sbox_10_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L16), .B0_t (SubBytesIns_Inst_Sbox_10_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L19), .B0_t (SubBytesIns_Inst_Sbox_10_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L6), .B0_t (SubBytesIns_Inst_Sbox_10_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L20), .B0_t (SubBytesIns_Inst_Sbox_10_L22), .Z0_t (MixColumnsInput[115]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L25), .B0_t (SubBytesIns_Inst_Sbox_10_L29), .Z0_t (MixColumnsInput[114]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L13), .B0_t (SubBytesIns_Inst_Sbox_10_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_10_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_10_L6), .B0_t (SubBytesIns_Inst_Sbox_10_L23), .Z0_t (MixColumnsInput[112]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T1_U1 ( .A0_t (ciphertext[95]), .B0_t (ciphertext[92]), .Z0_t (SubBytesIns_Inst_Sbox_11_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T2_U1 ( .A0_t (ciphertext[95]), .B0_t (ciphertext[90]), .Z0_t (SubBytesIns_Inst_Sbox_11_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T3_U1 ( .A0_t (ciphertext[95]), .B0_t (ciphertext[89]), .Z0_t (SubBytesIns_Inst_Sbox_11_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T4_U1 ( .A0_t (ciphertext[92]), .B0_t (ciphertext[90]), .Z0_t (SubBytesIns_Inst_Sbox_11_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T5_U1 ( .A0_t (ciphertext[91]), .B0_t (ciphertext[89]), .Z0_t (SubBytesIns_Inst_Sbox_11_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T1), .B0_t (SubBytesIns_Inst_Sbox_11_T5), .Z0_t (SubBytesIns_Inst_Sbox_11_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T7_U1 ( .A0_t (ciphertext[94]), .B0_t (ciphertext[93]), .Z0_t (SubBytesIns_Inst_Sbox_11_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T8_U1 ( .A0_t (ciphertext[88]), .B0_t (SubBytesIns_Inst_Sbox_11_T6), .Z0_t (SubBytesIns_Inst_Sbox_11_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T9_U1 ( .A0_t (ciphertext[88]), .B0_t (SubBytesIns_Inst_Sbox_11_T7), .Z0_t (SubBytesIns_Inst_Sbox_11_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T6), .B0_t (SubBytesIns_Inst_Sbox_11_T7), .Z0_t (SubBytesIns_Inst_Sbox_11_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T11_U1 ( .A0_t (ciphertext[94]), .B0_t (ciphertext[90]), .Z0_t (SubBytesIns_Inst_Sbox_11_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T12_U1 ( .A0_t (ciphertext[93]), .B0_t (ciphertext[90]), .Z0_t (SubBytesIns_Inst_Sbox_11_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T3), .B0_t (SubBytesIns_Inst_Sbox_11_T4), .Z0_t (SubBytesIns_Inst_Sbox_11_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T6), .B0_t (SubBytesIns_Inst_Sbox_11_T11), .Z0_t (SubBytesIns_Inst_Sbox_11_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T5), .B0_t (SubBytesIns_Inst_Sbox_11_T11), .Z0_t (SubBytesIns_Inst_Sbox_11_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T5), .B0_t (SubBytesIns_Inst_Sbox_11_T12), .Z0_t (SubBytesIns_Inst_Sbox_11_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T9), .B0_t (SubBytesIns_Inst_Sbox_11_T16), .Z0_t (SubBytesIns_Inst_Sbox_11_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T18_U1 ( .A0_t (ciphertext[92]), .B0_t (ciphertext[88]), .Z0_t (SubBytesIns_Inst_Sbox_11_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T7), .B0_t (SubBytesIns_Inst_Sbox_11_T18), .Z0_t (SubBytesIns_Inst_Sbox_11_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T1), .B0_t (SubBytesIns_Inst_Sbox_11_T19), .Z0_t (SubBytesIns_Inst_Sbox_11_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T21_U1 ( .A0_t (ciphertext[89]), .B0_t (ciphertext[88]), .Z0_t (SubBytesIns_Inst_Sbox_11_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T7), .B0_t (SubBytesIns_Inst_Sbox_11_T21), .Z0_t (SubBytesIns_Inst_Sbox_11_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T2), .B0_t (SubBytesIns_Inst_Sbox_11_T22), .Z0_t (SubBytesIns_Inst_Sbox_11_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T2), .B0_t (SubBytesIns_Inst_Sbox_11_T10), .Z0_t (SubBytesIns_Inst_Sbox_11_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T20), .B0_t (SubBytesIns_Inst_Sbox_11_T17), .Z0_t (SubBytesIns_Inst_Sbox_11_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T3), .B0_t (SubBytesIns_Inst_Sbox_11_T16), .Z0_t (SubBytesIns_Inst_Sbox_11_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T1), .B0_t (SubBytesIns_Inst_Sbox_11_T12), .Z0_t (SubBytesIns_Inst_Sbox_11_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T13), .B0_t (SubBytesIns_Inst_Sbox_11_T6), .Z0_t (SubBytesIns_Inst_Sbox_11_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T23), .B0_t (SubBytesIns_Inst_Sbox_11_T8), .Z0_t (SubBytesIns_Inst_Sbox_11_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T14), .B0_t (SubBytesIns_Inst_Sbox_11_M1), .Z0_t (SubBytesIns_Inst_Sbox_11_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T19), .B0_t (ciphertext[88]), .Z0_t (SubBytesIns_Inst_Sbox_11_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M4), .B0_t (SubBytesIns_Inst_Sbox_11_M1), .Z0_t (SubBytesIns_Inst_Sbox_11_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T3), .B0_t (SubBytesIns_Inst_Sbox_11_T16), .Z0_t (SubBytesIns_Inst_Sbox_11_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T22), .B0_t (SubBytesIns_Inst_Sbox_11_T9), .Z0_t (SubBytesIns_Inst_Sbox_11_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T26), .B0_t (SubBytesIns_Inst_Sbox_11_M6), .Z0_t (SubBytesIns_Inst_Sbox_11_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T20), .B0_t (SubBytesIns_Inst_Sbox_11_T17), .Z0_t (SubBytesIns_Inst_Sbox_11_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M9), .B0_t (SubBytesIns_Inst_Sbox_11_M6), .Z0_t (SubBytesIns_Inst_Sbox_11_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T1), .B0_t (SubBytesIns_Inst_Sbox_11_T15), .Z0_t (SubBytesIns_Inst_Sbox_11_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T4), .B0_t (SubBytesIns_Inst_Sbox_11_T27), .Z0_t (SubBytesIns_Inst_Sbox_11_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M12), .B0_t (SubBytesIns_Inst_Sbox_11_M11), .Z0_t (SubBytesIns_Inst_Sbox_11_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_T2), .B0_t (SubBytesIns_Inst_Sbox_11_T10), .Z0_t (SubBytesIns_Inst_Sbox_11_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M14), .B0_t (SubBytesIns_Inst_Sbox_11_M11), .Z0_t (SubBytesIns_Inst_Sbox_11_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M3), .B0_t (SubBytesIns_Inst_Sbox_11_M2), .Z0_t (SubBytesIns_Inst_Sbox_11_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M5), .B0_t (SubBytesIns_Inst_Sbox_11_T24), .Z0_t (SubBytesIns_Inst_Sbox_11_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M8), .B0_t (SubBytesIns_Inst_Sbox_11_M7), .Z0_t (SubBytesIns_Inst_Sbox_11_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M10), .B0_t (SubBytesIns_Inst_Sbox_11_M15), .Z0_t (SubBytesIns_Inst_Sbox_11_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M16), .B0_t (SubBytesIns_Inst_Sbox_11_M13), .Z0_t (SubBytesIns_Inst_Sbox_11_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M17), .B0_t (SubBytesIns_Inst_Sbox_11_M15), .Z0_t (SubBytesIns_Inst_Sbox_11_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M18), .B0_t (SubBytesIns_Inst_Sbox_11_M13), .Z0_t (SubBytesIns_Inst_Sbox_11_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M19), .B0_t (SubBytesIns_Inst_Sbox_11_T25), .Z0_t (SubBytesIns_Inst_Sbox_11_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M22), .B0_t (SubBytesIns_Inst_Sbox_11_M23), .Z0_t (SubBytesIns_Inst_Sbox_11_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M22), .B0_t (SubBytesIns_Inst_Sbox_11_M20), .Z0_t (SubBytesIns_Inst_Sbox_11_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M21), .B0_t (SubBytesIns_Inst_Sbox_11_M25), .Z0_t (SubBytesIns_Inst_Sbox_11_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M20), .B0_t (SubBytesIns_Inst_Sbox_11_M21), .Z0_t (SubBytesIns_Inst_Sbox_11_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M23), .B0_t (SubBytesIns_Inst_Sbox_11_M25), .Z0_t (SubBytesIns_Inst_Sbox_11_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M28), .B0_t (SubBytesIns_Inst_Sbox_11_M27), .Z0_t (SubBytesIns_Inst_Sbox_11_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M26), .B0_t (SubBytesIns_Inst_Sbox_11_M24), .Z0_t (SubBytesIns_Inst_Sbox_11_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M20), .B0_t (SubBytesIns_Inst_Sbox_11_M23), .Z0_t (SubBytesIns_Inst_Sbox_11_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M27), .B0_t (SubBytesIns_Inst_Sbox_11_M31), .Z0_t (SubBytesIns_Inst_Sbox_11_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M27), .B0_t (SubBytesIns_Inst_Sbox_11_M25), .Z0_t (SubBytesIns_Inst_Sbox_11_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M21), .B0_t (SubBytesIns_Inst_Sbox_11_M22), .Z0_t (SubBytesIns_Inst_Sbox_11_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M24), .B0_t (SubBytesIns_Inst_Sbox_11_M34), .Z0_t (SubBytesIns_Inst_Sbox_11_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M24), .B0_t (SubBytesIns_Inst_Sbox_11_M25), .Z0_t (SubBytesIns_Inst_Sbox_11_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M21), .B0_t (SubBytesIns_Inst_Sbox_11_M29), .Z0_t (SubBytesIns_Inst_Sbox_11_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M32), .B0_t (SubBytesIns_Inst_Sbox_11_M33), .Z0_t (SubBytesIns_Inst_Sbox_11_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M23), .B0_t (SubBytesIns_Inst_Sbox_11_M30), .Z0_t (SubBytesIns_Inst_Sbox_11_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M35), .B0_t (SubBytesIns_Inst_Sbox_11_M36), .Z0_t (SubBytesIns_Inst_Sbox_11_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M38), .B0_t (SubBytesIns_Inst_Sbox_11_M40), .Z0_t (SubBytesIns_Inst_Sbox_11_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M37), .B0_t (SubBytesIns_Inst_Sbox_11_M39), .Z0_t (SubBytesIns_Inst_Sbox_11_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M37), .B0_t (SubBytesIns_Inst_Sbox_11_M38), .Z0_t (SubBytesIns_Inst_Sbox_11_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M39), .B0_t (SubBytesIns_Inst_Sbox_11_M40), .Z0_t (SubBytesIns_Inst_Sbox_11_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M42), .B0_t (SubBytesIns_Inst_Sbox_11_M41), .Z0_t (SubBytesIns_Inst_Sbox_11_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M44), .B0_t (SubBytesIns_Inst_Sbox_11_T6), .Z0_t (SubBytesIns_Inst_Sbox_11_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M40), .B0_t (SubBytesIns_Inst_Sbox_11_T8), .Z0_t (SubBytesIns_Inst_Sbox_11_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M39), .B0_t (ciphertext[88]), .Z0_t (SubBytesIns_Inst_Sbox_11_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M43), .B0_t (SubBytesIns_Inst_Sbox_11_T16), .Z0_t (SubBytesIns_Inst_Sbox_11_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M38), .B0_t (SubBytesIns_Inst_Sbox_11_T9), .Z0_t (SubBytesIns_Inst_Sbox_11_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M37), .B0_t (SubBytesIns_Inst_Sbox_11_T17), .Z0_t (SubBytesIns_Inst_Sbox_11_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M42), .B0_t (SubBytesIns_Inst_Sbox_11_T15), .Z0_t (SubBytesIns_Inst_Sbox_11_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M45), .B0_t (SubBytesIns_Inst_Sbox_11_T27), .Z0_t (SubBytesIns_Inst_Sbox_11_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M41), .B0_t (SubBytesIns_Inst_Sbox_11_T10), .Z0_t (SubBytesIns_Inst_Sbox_11_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M44), .B0_t (SubBytesIns_Inst_Sbox_11_T13), .Z0_t (SubBytesIns_Inst_Sbox_11_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M40), .B0_t (SubBytesIns_Inst_Sbox_11_T23), .Z0_t (SubBytesIns_Inst_Sbox_11_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M39), .B0_t (SubBytesIns_Inst_Sbox_11_T19), .Z0_t (SubBytesIns_Inst_Sbox_11_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M43), .B0_t (SubBytesIns_Inst_Sbox_11_T3), .Z0_t (SubBytesIns_Inst_Sbox_11_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M38), .B0_t (SubBytesIns_Inst_Sbox_11_T22), .Z0_t (SubBytesIns_Inst_Sbox_11_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M37), .B0_t (SubBytesIns_Inst_Sbox_11_T20), .Z0_t (SubBytesIns_Inst_Sbox_11_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M42), .B0_t (SubBytesIns_Inst_Sbox_11_T1), .Z0_t (SubBytesIns_Inst_Sbox_11_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M45), .B0_t (SubBytesIns_Inst_Sbox_11_T4), .Z0_t (SubBytesIns_Inst_Sbox_11_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M41), .B0_t (SubBytesIns_Inst_Sbox_11_T2), .Z0_t (SubBytesIns_Inst_Sbox_11_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M61), .B0_t (SubBytesIns_Inst_Sbox_11_M62), .Z0_t (SubBytesIns_Inst_Sbox_11_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M50), .B0_t (SubBytesIns_Inst_Sbox_11_M56), .Z0_t (SubBytesIns_Inst_Sbox_11_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M46), .B0_t (SubBytesIns_Inst_Sbox_11_M48), .Z0_t (SubBytesIns_Inst_Sbox_11_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M47), .B0_t (SubBytesIns_Inst_Sbox_11_M55), .Z0_t (SubBytesIns_Inst_Sbox_11_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M54), .B0_t (SubBytesIns_Inst_Sbox_11_M58), .Z0_t (SubBytesIns_Inst_Sbox_11_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M49), .B0_t (SubBytesIns_Inst_Sbox_11_M61), .Z0_t (SubBytesIns_Inst_Sbox_11_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M62), .B0_t (SubBytesIns_Inst_Sbox_11_L5), .Z0_t (SubBytesIns_Inst_Sbox_11_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M46), .B0_t (SubBytesIns_Inst_Sbox_11_L3), .Z0_t (SubBytesIns_Inst_Sbox_11_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M51), .B0_t (SubBytesIns_Inst_Sbox_11_M59), .Z0_t (SubBytesIns_Inst_Sbox_11_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M52), .B0_t (SubBytesIns_Inst_Sbox_11_M53), .Z0_t (SubBytesIns_Inst_Sbox_11_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M53), .B0_t (SubBytesIns_Inst_Sbox_11_L4), .Z0_t (SubBytesIns_Inst_Sbox_11_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M60), .B0_t (SubBytesIns_Inst_Sbox_11_L2), .Z0_t (SubBytesIns_Inst_Sbox_11_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M48), .B0_t (SubBytesIns_Inst_Sbox_11_M51), .Z0_t (SubBytesIns_Inst_Sbox_11_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M50), .B0_t (SubBytesIns_Inst_Sbox_11_L0), .Z0_t (SubBytesIns_Inst_Sbox_11_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M52), .B0_t (SubBytesIns_Inst_Sbox_11_M61), .Z0_t (SubBytesIns_Inst_Sbox_11_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M55), .B0_t (SubBytesIns_Inst_Sbox_11_L1), .Z0_t (SubBytesIns_Inst_Sbox_11_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M56), .B0_t (SubBytesIns_Inst_Sbox_11_L0), .Z0_t (SubBytesIns_Inst_Sbox_11_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M57), .B0_t (SubBytesIns_Inst_Sbox_11_L1), .Z0_t (SubBytesIns_Inst_Sbox_11_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M58), .B0_t (SubBytesIns_Inst_Sbox_11_L8), .Z0_t (SubBytesIns_Inst_Sbox_11_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_M63), .B0_t (SubBytesIns_Inst_Sbox_11_L4), .Z0_t (SubBytesIns_Inst_Sbox_11_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L0), .B0_t (SubBytesIns_Inst_Sbox_11_L1), .Z0_t (SubBytesIns_Inst_Sbox_11_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L1), .B0_t (SubBytesIns_Inst_Sbox_11_L7), .Z0_t (SubBytesIns_Inst_Sbox_11_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L3), .B0_t (SubBytesIns_Inst_Sbox_11_L12), .Z0_t (SubBytesIns_Inst_Sbox_11_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L18), .B0_t (SubBytesIns_Inst_Sbox_11_L2), .Z0_t (SubBytesIns_Inst_Sbox_11_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L15), .B0_t (SubBytesIns_Inst_Sbox_11_L9), .Z0_t (SubBytesIns_Inst_Sbox_11_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L6), .B0_t (SubBytesIns_Inst_Sbox_11_L10), .Z0_t (SubBytesIns_Inst_Sbox_11_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L7), .B0_t (SubBytesIns_Inst_Sbox_11_L9), .Z0_t (SubBytesIns_Inst_Sbox_11_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L8), .B0_t (SubBytesIns_Inst_Sbox_11_L10), .Z0_t (SubBytesIns_Inst_Sbox_11_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L11), .B0_t (SubBytesIns_Inst_Sbox_11_L14), .Z0_t (SubBytesIns_Inst_Sbox_11_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L11), .B0_t (SubBytesIns_Inst_Sbox_11_L17), .Z0_t (SubBytesIns_Inst_Sbox_11_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L6), .B0_t (SubBytesIns_Inst_Sbox_11_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L16), .B0_t (SubBytesIns_Inst_Sbox_11_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L19), .B0_t (SubBytesIns_Inst_Sbox_11_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L6), .B0_t (SubBytesIns_Inst_Sbox_11_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L20), .B0_t (SubBytesIns_Inst_Sbox_11_L22), .Z0_t (MixColumnsInput[91]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L25), .B0_t (SubBytesIns_Inst_Sbox_11_L29), .Z0_t (MixColumnsInput[90]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L13), .B0_t (SubBytesIns_Inst_Sbox_11_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_11_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_11_L6), .B0_t (SubBytesIns_Inst_Sbox_11_L23), .Z0_t (MixColumnsInput[88]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T1_U1 ( .A0_t (ciphertext[103]), .B0_t (ciphertext[100]), .Z0_t (SubBytesIns_Inst_Sbox_12_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T2_U1 ( .A0_t (ciphertext[103]), .B0_t (ciphertext[98]), .Z0_t (SubBytesIns_Inst_Sbox_12_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T3_U1 ( .A0_t (ciphertext[103]), .B0_t (ciphertext[97]), .Z0_t (SubBytesIns_Inst_Sbox_12_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T4_U1 ( .A0_t (ciphertext[100]), .B0_t (ciphertext[98]), .Z0_t (SubBytesIns_Inst_Sbox_12_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T5_U1 ( .A0_t (ciphertext[99]), .B0_t (ciphertext[97]), .Z0_t (SubBytesIns_Inst_Sbox_12_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T1), .B0_t (SubBytesIns_Inst_Sbox_12_T5), .Z0_t (SubBytesIns_Inst_Sbox_12_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T7_U1 ( .A0_t (ciphertext[102]), .B0_t (ciphertext[101]), .Z0_t (SubBytesIns_Inst_Sbox_12_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T8_U1 ( .A0_t (ciphertext[96]), .B0_t (SubBytesIns_Inst_Sbox_12_T6), .Z0_t (SubBytesIns_Inst_Sbox_12_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T9_U1 ( .A0_t (ciphertext[96]), .B0_t (SubBytesIns_Inst_Sbox_12_T7), .Z0_t (SubBytesIns_Inst_Sbox_12_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T6), .B0_t (SubBytesIns_Inst_Sbox_12_T7), .Z0_t (SubBytesIns_Inst_Sbox_12_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T11_U1 ( .A0_t (ciphertext[102]), .B0_t (ciphertext[98]), .Z0_t (SubBytesIns_Inst_Sbox_12_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T12_U1 ( .A0_t (ciphertext[101]), .B0_t (ciphertext[98]), .Z0_t (SubBytesIns_Inst_Sbox_12_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T3), .B0_t (SubBytesIns_Inst_Sbox_12_T4), .Z0_t (SubBytesIns_Inst_Sbox_12_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T6), .B0_t (SubBytesIns_Inst_Sbox_12_T11), .Z0_t (SubBytesIns_Inst_Sbox_12_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T5), .B0_t (SubBytesIns_Inst_Sbox_12_T11), .Z0_t (SubBytesIns_Inst_Sbox_12_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T5), .B0_t (SubBytesIns_Inst_Sbox_12_T12), .Z0_t (SubBytesIns_Inst_Sbox_12_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T9), .B0_t (SubBytesIns_Inst_Sbox_12_T16), .Z0_t (SubBytesIns_Inst_Sbox_12_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T18_U1 ( .A0_t (ciphertext[100]), .B0_t (ciphertext[96]), .Z0_t (SubBytesIns_Inst_Sbox_12_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T7), .B0_t (SubBytesIns_Inst_Sbox_12_T18), .Z0_t (SubBytesIns_Inst_Sbox_12_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T1), .B0_t (SubBytesIns_Inst_Sbox_12_T19), .Z0_t (SubBytesIns_Inst_Sbox_12_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T21_U1 ( .A0_t (ciphertext[97]), .B0_t (ciphertext[96]), .Z0_t (SubBytesIns_Inst_Sbox_12_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T7), .B0_t (SubBytesIns_Inst_Sbox_12_T21), .Z0_t (SubBytesIns_Inst_Sbox_12_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T2), .B0_t (SubBytesIns_Inst_Sbox_12_T22), .Z0_t (SubBytesIns_Inst_Sbox_12_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T2), .B0_t (SubBytesIns_Inst_Sbox_12_T10), .Z0_t (SubBytesIns_Inst_Sbox_12_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T20), .B0_t (SubBytesIns_Inst_Sbox_12_T17), .Z0_t (SubBytesIns_Inst_Sbox_12_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T3), .B0_t (SubBytesIns_Inst_Sbox_12_T16), .Z0_t (SubBytesIns_Inst_Sbox_12_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T1), .B0_t (SubBytesIns_Inst_Sbox_12_T12), .Z0_t (SubBytesIns_Inst_Sbox_12_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T13), .B0_t (SubBytesIns_Inst_Sbox_12_T6), .Z0_t (SubBytesIns_Inst_Sbox_12_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T23), .B0_t (SubBytesIns_Inst_Sbox_12_T8), .Z0_t (SubBytesIns_Inst_Sbox_12_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T14), .B0_t (SubBytesIns_Inst_Sbox_12_M1), .Z0_t (SubBytesIns_Inst_Sbox_12_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T19), .B0_t (ciphertext[96]), .Z0_t (SubBytesIns_Inst_Sbox_12_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M4), .B0_t (SubBytesIns_Inst_Sbox_12_M1), .Z0_t (SubBytesIns_Inst_Sbox_12_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T3), .B0_t (SubBytesIns_Inst_Sbox_12_T16), .Z0_t (SubBytesIns_Inst_Sbox_12_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T22), .B0_t (SubBytesIns_Inst_Sbox_12_T9), .Z0_t (SubBytesIns_Inst_Sbox_12_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T26), .B0_t (SubBytesIns_Inst_Sbox_12_M6), .Z0_t (SubBytesIns_Inst_Sbox_12_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T20), .B0_t (SubBytesIns_Inst_Sbox_12_T17), .Z0_t (SubBytesIns_Inst_Sbox_12_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M9), .B0_t (SubBytesIns_Inst_Sbox_12_M6), .Z0_t (SubBytesIns_Inst_Sbox_12_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T1), .B0_t (SubBytesIns_Inst_Sbox_12_T15), .Z0_t (SubBytesIns_Inst_Sbox_12_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T4), .B0_t (SubBytesIns_Inst_Sbox_12_T27), .Z0_t (SubBytesIns_Inst_Sbox_12_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M12), .B0_t (SubBytesIns_Inst_Sbox_12_M11), .Z0_t (SubBytesIns_Inst_Sbox_12_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_T2), .B0_t (SubBytesIns_Inst_Sbox_12_T10), .Z0_t (SubBytesIns_Inst_Sbox_12_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M14), .B0_t (SubBytesIns_Inst_Sbox_12_M11), .Z0_t (SubBytesIns_Inst_Sbox_12_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M3), .B0_t (SubBytesIns_Inst_Sbox_12_M2), .Z0_t (SubBytesIns_Inst_Sbox_12_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M5), .B0_t (SubBytesIns_Inst_Sbox_12_T24), .Z0_t (SubBytesIns_Inst_Sbox_12_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M8), .B0_t (SubBytesIns_Inst_Sbox_12_M7), .Z0_t (SubBytesIns_Inst_Sbox_12_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M10), .B0_t (SubBytesIns_Inst_Sbox_12_M15), .Z0_t (SubBytesIns_Inst_Sbox_12_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M16), .B0_t (SubBytesIns_Inst_Sbox_12_M13), .Z0_t (SubBytesIns_Inst_Sbox_12_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M17), .B0_t (SubBytesIns_Inst_Sbox_12_M15), .Z0_t (SubBytesIns_Inst_Sbox_12_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M18), .B0_t (SubBytesIns_Inst_Sbox_12_M13), .Z0_t (SubBytesIns_Inst_Sbox_12_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M19), .B0_t (SubBytesIns_Inst_Sbox_12_T25), .Z0_t (SubBytesIns_Inst_Sbox_12_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M22), .B0_t (SubBytesIns_Inst_Sbox_12_M23), .Z0_t (SubBytesIns_Inst_Sbox_12_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M22), .B0_t (SubBytesIns_Inst_Sbox_12_M20), .Z0_t (SubBytesIns_Inst_Sbox_12_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M21), .B0_t (SubBytesIns_Inst_Sbox_12_M25), .Z0_t (SubBytesIns_Inst_Sbox_12_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M20), .B0_t (SubBytesIns_Inst_Sbox_12_M21), .Z0_t (SubBytesIns_Inst_Sbox_12_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M23), .B0_t (SubBytesIns_Inst_Sbox_12_M25), .Z0_t (SubBytesIns_Inst_Sbox_12_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M28), .B0_t (SubBytesIns_Inst_Sbox_12_M27), .Z0_t (SubBytesIns_Inst_Sbox_12_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M26), .B0_t (SubBytesIns_Inst_Sbox_12_M24), .Z0_t (SubBytesIns_Inst_Sbox_12_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M20), .B0_t (SubBytesIns_Inst_Sbox_12_M23), .Z0_t (SubBytesIns_Inst_Sbox_12_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M27), .B0_t (SubBytesIns_Inst_Sbox_12_M31), .Z0_t (SubBytesIns_Inst_Sbox_12_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M27), .B0_t (SubBytesIns_Inst_Sbox_12_M25), .Z0_t (SubBytesIns_Inst_Sbox_12_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M21), .B0_t (SubBytesIns_Inst_Sbox_12_M22), .Z0_t (SubBytesIns_Inst_Sbox_12_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M24), .B0_t (SubBytesIns_Inst_Sbox_12_M34), .Z0_t (SubBytesIns_Inst_Sbox_12_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M24), .B0_t (SubBytesIns_Inst_Sbox_12_M25), .Z0_t (SubBytesIns_Inst_Sbox_12_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M21), .B0_t (SubBytesIns_Inst_Sbox_12_M29), .Z0_t (SubBytesIns_Inst_Sbox_12_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M32), .B0_t (SubBytesIns_Inst_Sbox_12_M33), .Z0_t (SubBytesIns_Inst_Sbox_12_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M23), .B0_t (SubBytesIns_Inst_Sbox_12_M30), .Z0_t (SubBytesIns_Inst_Sbox_12_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M35), .B0_t (SubBytesIns_Inst_Sbox_12_M36), .Z0_t (SubBytesIns_Inst_Sbox_12_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M38), .B0_t (SubBytesIns_Inst_Sbox_12_M40), .Z0_t (SubBytesIns_Inst_Sbox_12_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M37), .B0_t (SubBytesIns_Inst_Sbox_12_M39), .Z0_t (SubBytesIns_Inst_Sbox_12_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M37), .B0_t (SubBytesIns_Inst_Sbox_12_M38), .Z0_t (SubBytesIns_Inst_Sbox_12_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M39), .B0_t (SubBytesIns_Inst_Sbox_12_M40), .Z0_t (SubBytesIns_Inst_Sbox_12_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M42), .B0_t (SubBytesIns_Inst_Sbox_12_M41), .Z0_t (SubBytesIns_Inst_Sbox_12_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M44), .B0_t (SubBytesIns_Inst_Sbox_12_T6), .Z0_t (SubBytesIns_Inst_Sbox_12_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M40), .B0_t (SubBytesIns_Inst_Sbox_12_T8), .Z0_t (SubBytesIns_Inst_Sbox_12_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M39), .B0_t (ciphertext[96]), .Z0_t (SubBytesIns_Inst_Sbox_12_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M43), .B0_t (SubBytesIns_Inst_Sbox_12_T16), .Z0_t (SubBytesIns_Inst_Sbox_12_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M38), .B0_t (SubBytesIns_Inst_Sbox_12_T9), .Z0_t (SubBytesIns_Inst_Sbox_12_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M37), .B0_t (SubBytesIns_Inst_Sbox_12_T17), .Z0_t (SubBytesIns_Inst_Sbox_12_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M42), .B0_t (SubBytesIns_Inst_Sbox_12_T15), .Z0_t (SubBytesIns_Inst_Sbox_12_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M45), .B0_t (SubBytesIns_Inst_Sbox_12_T27), .Z0_t (SubBytesIns_Inst_Sbox_12_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M41), .B0_t (SubBytesIns_Inst_Sbox_12_T10), .Z0_t (SubBytesIns_Inst_Sbox_12_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M44), .B0_t (SubBytesIns_Inst_Sbox_12_T13), .Z0_t (SubBytesIns_Inst_Sbox_12_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M40), .B0_t (SubBytesIns_Inst_Sbox_12_T23), .Z0_t (SubBytesIns_Inst_Sbox_12_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M39), .B0_t (SubBytesIns_Inst_Sbox_12_T19), .Z0_t (SubBytesIns_Inst_Sbox_12_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M43), .B0_t (SubBytesIns_Inst_Sbox_12_T3), .Z0_t (SubBytesIns_Inst_Sbox_12_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M38), .B0_t (SubBytesIns_Inst_Sbox_12_T22), .Z0_t (SubBytesIns_Inst_Sbox_12_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M37), .B0_t (SubBytesIns_Inst_Sbox_12_T20), .Z0_t (SubBytesIns_Inst_Sbox_12_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M42), .B0_t (SubBytesIns_Inst_Sbox_12_T1), .Z0_t (SubBytesIns_Inst_Sbox_12_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M45), .B0_t (SubBytesIns_Inst_Sbox_12_T4), .Z0_t (SubBytesIns_Inst_Sbox_12_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M41), .B0_t (SubBytesIns_Inst_Sbox_12_T2), .Z0_t (SubBytesIns_Inst_Sbox_12_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M61), .B0_t (SubBytesIns_Inst_Sbox_12_M62), .Z0_t (SubBytesIns_Inst_Sbox_12_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M50), .B0_t (SubBytesIns_Inst_Sbox_12_M56), .Z0_t (SubBytesIns_Inst_Sbox_12_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M46), .B0_t (SubBytesIns_Inst_Sbox_12_M48), .Z0_t (SubBytesIns_Inst_Sbox_12_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M47), .B0_t (SubBytesIns_Inst_Sbox_12_M55), .Z0_t (SubBytesIns_Inst_Sbox_12_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M54), .B0_t (SubBytesIns_Inst_Sbox_12_M58), .Z0_t (SubBytesIns_Inst_Sbox_12_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M49), .B0_t (SubBytesIns_Inst_Sbox_12_M61), .Z0_t (SubBytesIns_Inst_Sbox_12_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M62), .B0_t (SubBytesIns_Inst_Sbox_12_L5), .Z0_t (SubBytesIns_Inst_Sbox_12_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M46), .B0_t (SubBytesIns_Inst_Sbox_12_L3), .Z0_t (SubBytesIns_Inst_Sbox_12_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M51), .B0_t (SubBytesIns_Inst_Sbox_12_M59), .Z0_t (SubBytesIns_Inst_Sbox_12_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M52), .B0_t (SubBytesIns_Inst_Sbox_12_M53), .Z0_t (SubBytesIns_Inst_Sbox_12_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M53), .B0_t (SubBytesIns_Inst_Sbox_12_L4), .Z0_t (SubBytesIns_Inst_Sbox_12_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M60), .B0_t (SubBytesIns_Inst_Sbox_12_L2), .Z0_t (SubBytesIns_Inst_Sbox_12_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M48), .B0_t (SubBytesIns_Inst_Sbox_12_M51), .Z0_t (SubBytesIns_Inst_Sbox_12_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M50), .B0_t (SubBytesIns_Inst_Sbox_12_L0), .Z0_t (SubBytesIns_Inst_Sbox_12_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M52), .B0_t (SubBytesIns_Inst_Sbox_12_M61), .Z0_t (SubBytesIns_Inst_Sbox_12_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M55), .B0_t (SubBytesIns_Inst_Sbox_12_L1), .Z0_t (SubBytesIns_Inst_Sbox_12_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M56), .B0_t (SubBytesIns_Inst_Sbox_12_L0), .Z0_t (SubBytesIns_Inst_Sbox_12_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M57), .B0_t (SubBytesIns_Inst_Sbox_12_L1), .Z0_t (SubBytesIns_Inst_Sbox_12_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M58), .B0_t (SubBytesIns_Inst_Sbox_12_L8), .Z0_t (SubBytesIns_Inst_Sbox_12_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_M63), .B0_t (SubBytesIns_Inst_Sbox_12_L4), .Z0_t (SubBytesIns_Inst_Sbox_12_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L0), .B0_t (SubBytesIns_Inst_Sbox_12_L1), .Z0_t (SubBytesIns_Inst_Sbox_12_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L1), .B0_t (SubBytesIns_Inst_Sbox_12_L7), .Z0_t (SubBytesIns_Inst_Sbox_12_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L3), .B0_t (SubBytesIns_Inst_Sbox_12_L12), .Z0_t (SubBytesIns_Inst_Sbox_12_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L18), .B0_t (SubBytesIns_Inst_Sbox_12_L2), .Z0_t (SubBytesIns_Inst_Sbox_12_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L15), .B0_t (SubBytesIns_Inst_Sbox_12_L9), .Z0_t (SubBytesIns_Inst_Sbox_12_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L6), .B0_t (SubBytesIns_Inst_Sbox_12_L10), .Z0_t (SubBytesIns_Inst_Sbox_12_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L7), .B0_t (SubBytesIns_Inst_Sbox_12_L9), .Z0_t (SubBytesIns_Inst_Sbox_12_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L8), .B0_t (SubBytesIns_Inst_Sbox_12_L10), .Z0_t (SubBytesIns_Inst_Sbox_12_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L11), .B0_t (SubBytesIns_Inst_Sbox_12_L14), .Z0_t (SubBytesIns_Inst_Sbox_12_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L11), .B0_t (SubBytesIns_Inst_Sbox_12_L17), .Z0_t (SubBytesIns_Inst_Sbox_12_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L6), .B0_t (SubBytesIns_Inst_Sbox_12_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L16), .B0_t (SubBytesIns_Inst_Sbox_12_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L19), .B0_t (SubBytesIns_Inst_Sbox_12_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L6), .B0_t (SubBytesIns_Inst_Sbox_12_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L20), .B0_t (SubBytesIns_Inst_Sbox_12_L22), .Z0_t (MixColumnsInput[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L25), .B0_t (SubBytesIns_Inst_Sbox_12_L29), .Z0_t (MixColumnsInput[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L13), .B0_t (SubBytesIns_Inst_Sbox_12_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_12_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_12_L6), .B0_t (SubBytesIns_Inst_Sbox_12_L23), .Z0_t (MixColumnsInput[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T1_U1 ( .A0_t (ciphertext[111]), .B0_t (ciphertext[108]), .Z0_t (SubBytesIns_Inst_Sbox_13_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T2_U1 ( .A0_t (ciphertext[111]), .B0_t (ciphertext[106]), .Z0_t (SubBytesIns_Inst_Sbox_13_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T3_U1 ( .A0_t (ciphertext[111]), .B0_t (ciphertext[105]), .Z0_t (SubBytesIns_Inst_Sbox_13_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T4_U1 ( .A0_t (ciphertext[108]), .B0_t (ciphertext[106]), .Z0_t (SubBytesIns_Inst_Sbox_13_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T5_U1 ( .A0_t (ciphertext[107]), .B0_t (ciphertext[105]), .Z0_t (SubBytesIns_Inst_Sbox_13_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T1), .B0_t (SubBytesIns_Inst_Sbox_13_T5), .Z0_t (SubBytesIns_Inst_Sbox_13_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T7_U1 ( .A0_t (ciphertext[110]), .B0_t (ciphertext[109]), .Z0_t (SubBytesIns_Inst_Sbox_13_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T8_U1 ( .A0_t (ciphertext[104]), .B0_t (SubBytesIns_Inst_Sbox_13_T6), .Z0_t (SubBytesIns_Inst_Sbox_13_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T9_U1 ( .A0_t (ciphertext[104]), .B0_t (SubBytesIns_Inst_Sbox_13_T7), .Z0_t (SubBytesIns_Inst_Sbox_13_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T6), .B0_t (SubBytesIns_Inst_Sbox_13_T7), .Z0_t (SubBytesIns_Inst_Sbox_13_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T11_U1 ( .A0_t (ciphertext[110]), .B0_t (ciphertext[106]), .Z0_t (SubBytesIns_Inst_Sbox_13_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T12_U1 ( .A0_t (ciphertext[109]), .B0_t (ciphertext[106]), .Z0_t (SubBytesIns_Inst_Sbox_13_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T3), .B0_t (SubBytesIns_Inst_Sbox_13_T4), .Z0_t (SubBytesIns_Inst_Sbox_13_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T6), .B0_t (SubBytesIns_Inst_Sbox_13_T11), .Z0_t (SubBytesIns_Inst_Sbox_13_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T5), .B0_t (SubBytesIns_Inst_Sbox_13_T11), .Z0_t (SubBytesIns_Inst_Sbox_13_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T5), .B0_t (SubBytesIns_Inst_Sbox_13_T12), .Z0_t (SubBytesIns_Inst_Sbox_13_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T9), .B0_t (SubBytesIns_Inst_Sbox_13_T16), .Z0_t (SubBytesIns_Inst_Sbox_13_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T18_U1 ( .A0_t (ciphertext[108]), .B0_t (ciphertext[104]), .Z0_t (SubBytesIns_Inst_Sbox_13_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T7), .B0_t (SubBytesIns_Inst_Sbox_13_T18), .Z0_t (SubBytesIns_Inst_Sbox_13_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T1), .B0_t (SubBytesIns_Inst_Sbox_13_T19), .Z0_t (SubBytesIns_Inst_Sbox_13_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T21_U1 ( .A0_t (ciphertext[105]), .B0_t (ciphertext[104]), .Z0_t (SubBytesIns_Inst_Sbox_13_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T7), .B0_t (SubBytesIns_Inst_Sbox_13_T21), .Z0_t (SubBytesIns_Inst_Sbox_13_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T2), .B0_t (SubBytesIns_Inst_Sbox_13_T22), .Z0_t (SubBytesIns_Inst_Sbox_13_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T2), .B0_t (SubBytesIns_Inst_Sbox_13_T10), .Z0_t (SubBytesIns_Inst_Sbox_13_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T20), .B0_t (SubBytesIns_Inst_Sbox_13_T17), .Z0_t (SubBytesIns_Inst_Sbox_13_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T3), .B0_t (SubBytesIns_Inst_Sbox_13_T16), .Z0_t (SubBytesIns_Inst_Sbox_13_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T1), .B0_t (SubBytesIns_Inst_Sbox_13_T12), .Z0_t (SubBytesIns_Inst_Sbox_13_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T13), .B0_t (SubBytesIns_Inst_Sbox_13_T6), .Z0_t (SubBytesIns_Inst_Sbox_13_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T23), .B0_t (SubBytesIns_Inst_Sbox_13_T8), .Z0_t (SubBytesIns_Inst_Sbox_13_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T14), .B0_t (SubBytesIns_Inst_Sbox_13_M1), .Z0_t (SubBytesIns_Inst_Sbox_13_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T19), .B0_t (ciphertext[104]), .Z0_t (SubBytesIns_Inst_Sbox_13_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M4), .B0_t (SubBytesIns_Inst_Sbox_13_M1), .Z0_t (SubBytesIns_Inst_Sbox_13_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T3), .B0_t (SubBytesIns_Inst_Sbox_13_T16), .Z0_t (SubBytesIns_Inst_Sbox_13_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T22), .B0_t (SubBytesIns_Inst_Sbox_13_T9), .Z0_t (SubBytesIns_Inst_Sbox_13_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T26), .B0_t (SubBytesIns_Inst_Sbox_13_M6), .Z0_t (SubBytesIns_Inst_Sbox_13_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T20), .B0_t (SubBytesIns_Inst_Sbox_13_T17), .Z0_t (SubBytesIns_Inst_Sbox_13_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M9), .B0_t (SubBytesIns_Inst_Sbox_13_M6), .Z0_t (SubBytesIns_Inst_Sbox_13_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T1), .B0_t (SubBytesIns_Inst_Sbox_13_T15), .Z0_t (SubBytesIns_Inst_Sbox_13_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T4), .B0_t (SubBytesIns_Inst_Sbox_13_T27), .Z0_t (SubBytesIns_Inst_Sbox_13_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M12), .B0_t (SubBytesIns_Inst_Sbox_13_M11), .Z0_t (SubBytesIns_Inst_Sbox_13_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_T2), .B0_t (SubBytesIns_Inst_Sbox_13_T10), .Z0_t (SubBytesIns_Inst_Sbox_13_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M14), .B0_t (SubBytesIns_Inst_Sbox_13_M11), .Z0_t (SubBytesIns_Inst_Sbox_13_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M3), .B0_t (SubBytesIns_Inst_Sbox_13_M2), .Z0_t (SubBytesIns_Inst_Sbox_13_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M5), .B0_t (SubBytesIns_Inst_Sbox_13_T24), .Z0_t (SubBytesIns_Inst_Sbox_13_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M8), .B0_t (SubBytesIns_Inst_Sbox_13_M7), .Z0_t (SubBytesIns_Inst_Sbox_13_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M10), .B0_t (SubBytesIns_Inst_Sbox_13_M15), .Z0_t (SubBytesIns_Inst_Sbox_13_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M16), .B0_t (SubBytesIns_Inst_Sbox_13_M13), .Z0_t (SubBytesIns_Inst_Sbox_13_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M17), .B0_t (SubBytesIns_Inst_Sbox_13_M15), .Z0_t (SubBytesIns_Inst_Sbox_13_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M18), .B0_t (SubBytesIns_Inst_Sbox_13_M13), .Z0_t (SubBytesIns_Inst_Sbox_13_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M19), .B0_t (SubBytesIns_Inst_Sbox_13_T25), .Z0_t (SubBytesIns_Inst_Sbox_13_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M22), .B0_t (SubBytesIns_Inst_Sbox_13_M23), .Z0_t (SubBytesIns_Inst_Sbox_13_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M22), .B0_t (SubBytesIns_Inst_Sbox_13_M20), .Z0_t (SubBytesIns_Inst_Sbox_13_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M21), .B0_t (SubBytesIns_Inst_Sbox_13_M25), .Z0_t (SubBytesIns_Inst_Sbox_13_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M20), .B0_t (SubBytesIns_Inst_Sbox_13_M21), .Z0_t (SubBytesIns_Inst_Sbox_13_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M23), .B0_t (SubBytesIns_Inst_Sbox_13_M25), .Z0_t (SubBytesIns_Inst_Sbox_13_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M28), .B0_t (SubBytesIns_Inst_Sbox_13_M27), .Z0_t (SubBytesIns_Inst_Sbox_13_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M26), .B0_t (SubBytesIns_Inst_Sbox_13_M24), .Z0_t (SubBytesIns_Inst_Sbox_13_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M20), .B0_t (SubBytesIns_Inst_Sbox_13_M23), .Z0_t (SubBytesIns_Inst_Sbox_13_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M27), .B0_t (SubBytesIns_Inst_Sbox_13_M31), .Z0_t (SubBytesIns_Inst_Sbox_13_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M27), .B0_t (SubBytesIns_Inst_Sbox_13_M25), .Z0_t (SubBytesIns_Inst_Sbox_13_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M21), .B0_t (SubBytesIns_Inst_Sbox_13_M22), .Z0_t (SubBytesIns_Inst_Sbox_13_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M24), .B0_t (SubBytesIns_Inst_Sbox_13_M34), .Z0_t (SubBytesIns_Inst_Sbox_13_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M24), .B0_t (SubBytesIns_Inst_Sbox_13_M25), .Z0_t (SubBytesIns_Inst_Sbox_13_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M21), .B0_t (SubBytesIns_Inst_Sbox_13_M29), .Z0_t (SubBytesIns_Inst_Sbox_13_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M32), .B0_t (SubBytesIns_Inst_Sbox_13_M33), .Z0_t (SubBytesIns_Inst_Sbox_13_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M23), .B0_t (SubBytesIns_Inst_Sbox_13_M30), .Z0_t (SubBytesIns_Inst_Sbox_13_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M35), .B0_t (SubBytesIns_Inst_Sbox_13_M36), .Z0_t (SubBytesIns_Inst_Sbox_13_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M38), .B0_t (SubBytesIns_Inst_Sbox_13_M40), .Z0_t (SubBytesIns_Inst_Sbox_13_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M37), .B0_t (SubBytesIns_Inst_Sbox_13_M39), .Z0_t (SubBytesIns_Inst_Sbox_13_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M37), .B0_t (SubBytesIns_Inst_Sbox_13_M38), .Z0_t (SubBytesIns_Inst_Sbox_13_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M39), .B0_t (SubBytesIns_Inst_Sbox_13_M40), .Z0_t (SubBytesIns_Inst_Sbox_13_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M42), .B0_t (SubBytesIns_Inst_Sbox_13_M41), .Z0_t (SubBytesIns_Inst_Sbox_13_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M44), .B0_t (SubBytesIns_Inst_Sbox_13_T6), .Z0_t (SubBytesIns_Inst_Sbox_13_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M40), .B0_t (SubBytesIns_Inst_Sbox_13_T8), .Z0_t (SubBytesIns_Inst_Sbox_13_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M39), .B0_t (ciphertext[104]), .Z0_t (SubBytesIns_Inst_Sbox_13_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M43), .B0_t (SubBytesIns_Inst_Sbox_13_T16), .Z0_t (SubBytesIns_Inst_Sbox_13_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M38), .B0_t (SubBytesIns_Inst_Sbox_13_T9), .Z0_t (SubBytesIns_Inst_Sbox_13_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M37), .B0_t (SubBytesIns_Inst_Sbox_13_T17), .Z0_t (SubBytesIns_Inst_Sbox_13_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M42), .B0_t (SubBytesIns_Inst_Sbox_13_T15), .Z0_t (SubBytesIns_Inst_Sbox_13_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M45), .B0_t (SubBytesIns_Inst_Sbox_13_T27), .Z0_t (SubBytesIns_Inst_Sbox_13_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M41), .B0_t (SubBytesIns_Inst_Sbox_13_T10), .Z0_t (SubBytesIns_Inst_Sbox_13_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M44), .B0_t (SubBytesIns_Inst_Sbox_13_T13), .Z0_t (SubBytesIns_Inst_Sbox_13_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M40), .B0_t (SubBytesIns_Inst_Sbox_13_T23), .Z0_t (SubBytesIns_Inst_Sbox_13_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M39), .B0_t (SubBytesIns_Inst_Sbox_13_T19), .Z0_t (SubBytesIns_Inst_Sbox_13_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M43), .B0_t (SubBytesIns_Inst_Sbox_13_T3), .Z0_t (SubBytesIns_Inst_Sbox_13_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M38), .B0_t (SubBytesIns_Inst_Sbox_13_T22), .Z0_t (SubBytesIns_Inst_Sbox_13_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M37), .B0_t (SubBytesIns_Inst_Sbox_13_T20), .Z0_t (SubBytesIns_Inst_Sbox_13_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M42), .B0_t (SubBytesIns_Inst_Sbox_13_T1), .Z0_t (SubBytesIns_Inst_Sbox_13_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M45), .B0_t (SubBytesIns_Inst_Sbox_13_T4), .Z0_t (SubBytesIns_Inst_Sbox_13_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M41), .B0_t (SubBytesIns_Inst_Sbox_13_T2), .Z0_t (SubBytesIns_Inst_Sbox_13_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M61), .B0_t (SubBytesIns_Inst_Sbox_13_M62), .Z0_t (SubBytesIns_Inst_Sbox_13_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M50), .B0_t (SubBytesIns_Inst_Sbox_13_M56), .Z0_t (SubBytesIns_Inst_Sbox_13_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M46), .B0_t (SubBytesIns_Inst_Sbox_13_M48), .Z0_t (SubBytesIns_Inst_Sbox_13_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M47), .B0_t (SubBytesIns_Inst_Sbox_13_M55), .Z0_t (SubBytesIns_Inst_Sbox_13_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M54), .B0_t (SubBytesIns_Inst_Sbox_13_M58), .Z0_t (SubBytesIns_Inst_Sbox_13_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M49), .B0_t (SubBytesIns_Inst_Sbox_13_M61), .Z0_t (SubBytesIns_Inst_Sbox_13_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M62), .B0_t (SubBytesIns_Inst_Sbox_13_L5), .Z0_t (SubBytesIns_Inst_Sbox_13_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M46), .B0_t (SubBytesIns_Inst_Sbox_13_L3), .Z0_t (SubBytesIns_Inst_Sbox_13_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M51), .B0_t (SubBytesIns_Inst_Sbox_13_M59), .Z0_t (SubBytesIns_Inst_Sbox_13_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M52), .B0_t (SubBytesIns_Inst_Sbox_13_M53), .Z0_t (SubBytesIns_Inst_Sbox_13_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M53), .B0_t (SubBytesIns_Inst_Sbox_13_L4), .Z0_t (SubBytesIns_Inst_Sbox_13_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M60), .B0_t (SubBytesIns_Inst_Sbox_13_L2), .Z0_t (SubBytesIns_Inst_Sbox_13_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M48), .B0_t (SubBytesIns_Inst_Sbox_13_M51), .Z0_t (SubBytesIns_Inst_Sbox_13_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M50), .B0_t (SubBytesIns_Inst_Sbox_13_L0), .Z0_t (SubBytesIns_Inst_Sbox_13_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M52), .B0_t (SubBytesIns_Inst_Sbox_13_M61), .Z0_t (SubBytesIns_Inst_Sbox_13_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M55), .B0_t (SubBytesIns_Inst_Sbox_13_L1), .Z0_t (SubBytesIns_Inst_Sbox_13_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M56), .B0_t (SubBytesIns_Inst_Sbox_13_L0), .Z0_t (SubBytesIns_Inst_Sbox_13_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M57), .B0_t (SubBytesIns_Inst_Sbox_13_L1), .Z0_t (SubBytesIns_Inst_Sbox_13_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M58), .B0_t (SubBytesIns_Inst_Sbox_13_L8), .Z0_t (SubBytesIns_Inst_Sbox_13_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_M63), .B0_t (SubBytesIns_Inst_Sbox_13_L4), .Z0_t (SubBytesIns_Inst_Sbox_13_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L0), .B0_t (SubBytesIns_Inst_Sbox_13_L1), .Z0_t (SubBytesIns_Inst_Sbox_13_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L1), .B0_t (SubBytesIns_Inst_Sbox_13_L7), .Z0_t (SubBytesIns_Inst_Sbox_13_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L3), .B0_t (SubBytesIns_Inst_Sbox_13_L12), .Z0_t (SubBytesIns_Inst_Sbox_13_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L18), .B0_t (SubBytesIns_Inst_Sbox_13_L2), .Z0_t (SubBytesIns_Inst_Sbox_13_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L15), .B0_t (SubBytesIns_Inst_Sbox_13_L9), .Z0_t (SubBytesIns_Inst_Sbox_13_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L6), .B0_t (SubBytesIns_Inst_Sbox_13_L10), .Z0_t (SubBytesIns_Inst_Sbox_13_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L7), .B0_t (SubBytesIns_Inst_Sbox_13_L9), .Z0_t (SubBytesIns_Inst_Sbox_13_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L8), .B0_t (SubBytesIns_Inst_Sbox_13_L10), .Z0_t (SubBytesIns_Inst_Sbox_13_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L11), .B0_t (SubBytesIns_Inst_Sbox_13_L14), .Z0_t (SubBytesIns_Inst_Sbox_13_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L11), .B0_t (SubBytesIns_Inst_Sbox_13_L17), .Z0_t (SubBytesIns_Inst_Sbox_13_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L6), .B0_t (SubBytesIns_Inst_Sbox_13_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L16), .B0_t (SubBytesIns_Inst_Sbox_13_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L19), .B0_t (SubBytesIns_Inst_Sbox_13_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L6), .B0_t (SubBytesIns_Inst_Sbox_13_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L20), .B0_t (SubBytesIns_Inst_Sbox_13_L22), .Z0_t (MixColumnsInput[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L25), .B0_t (SubBytesIns_Inst_Sbox_13_L29), .Z0_t (MixColumnsInput[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L13), .B0_t (SubBytesIns_Inst_Sbox_13_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_13_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_13_L6), .B0_t (SubBytesIns_Inst_Sbox_13_L23), .Z0_t (MixColumnsInput[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T1_U1 ( .A0_t (ciphertext[119]), .B0_t (ciphertext[116]), .Z0_t (SubBytesIns_Inst_Sbox_14_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T2_U1 ( .A0_t (ciphertext[119]), .B0_t (ciphertext[114]), .Z0_t (SubBytesIns_Inst_Sbox_14_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T3_U1 ( .A0_t (ciphertext[119]), .B0_t (ciphertext[113]), .Z0_t (SubBytesIns_Inst_Sbox_14_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T4_U1 ( .A0_t (ciphertext[116]), .B0_t (ciphertext[114]), .Z0_t (SubBytesIns_Inst_Sbox_14_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T5_U1 ( .A0_t (ciphertext[115]), .B0_t (ciphertext[113]), .Z0_t (SubBytesIns_Inst_Sbox_14_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T1), .B0_t (SubBytesIns_Inst_Sbox_14_T5), .Z0_t (SubBytesIns_Inst_Sbox_14_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T7_U1 ( .A0_t (ciphertext[118]), .B0_t (ciphertext[117]), .Z0_t (SubBytesIns_Inst_Sbox_14_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T8_U1 ( .A0_t (ciphertext[112]), .B0_t (SubBytesIns_Inst_Sbox_14_T6), .Z0_t (SubBytesIns_Inst_Sbox_14_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T9_U1 ( .A0_t (ciphertext[112]), .B0_t (SubBytesIns_Inst_Sbox_14_T7), .Z0_t (SubBytesIns_Inst_Sbox_14_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T6), .B0_t (SubBytesIns_Inst_Sbox_14_T7), .Z0_t (SubBytesIns_Inst_Sbox_14_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T11_U1 ( .A0_t (ciphertext[118]), .B0_t (ciphertext[114]), .Z0_t (SubBytesIns_Inst_Sbox_14_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T12_U1 ( .A0_t (ciphertext[117]), .B0_t (ciphertext[114]), .Z0_t (SubBytesIns_Inst_Sbox_14_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T3), .B0_t (SubBytesIns_Inst_Sbox_14_T4), .Z0_t (SubBytesIns_Inst_Sbox_14_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T6), .B0_t (SubBytesIns_Inst_Sbox_14_T11), .Z0_t (SubBytesIns_Inst_Sbox_14_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T5), .B0_t (SubBytesIns_Inst_Sbox_14_T11), .Z0_t (SubBytesIns_Inst_Sbox_14_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T5), .B0_t (SubBytesIns_Inst_Sbox_14_T12), .Z0_t (SubBytesIns_Inst_Sbox_14_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T9), .B0_t (SubBytesIns_Inst_Sbox_14_T16), .Z0_t (SubBytesIns_Inst_Sbox_14_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T18_U1 ( .A0_t (ciphertext[116]), .B0_t (ciphertext[112]), .Z0_t (SubBytesIns_Inst_Sbox_14_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T7), .B0_t (SubBytesIns_Inst_Sbox_14_T18), .Z0_t (SubBytesIns_Inst_Sbox_14_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T1), .B0_t (SubBytesIns_Inst_Sbox_14_T19), .Z0_t (SubBytesIns_Inst_Sbox_14_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T21_U1 ( .A0_t (ciphertext[113]), .B0_t (ciphertext[112]), .Z0_t (SubBytesIns_Inst_Sbox_14_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T7), .B0_t (SubBytesIns_Inst_Sbox_14_T21), .Z0_t (SubBytesIns_Inst_Sbox_14_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T2), .B0_t (SubBytesIns_Inst_Sbox_14_T22), .Z0_t (SubBytesIns_Inst_Sbox_14_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T2), .B0_t (SubBytesIns_Inst_Sbox_14_T10), .Z0_t (SubBytesIns_Inst_Sbox_14_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T20), .B0_t (SubBytesIns_Inst_Sbox_14_T17), .Z0_t (SubBytesIns_Inst_Sbox_14_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T3), .B0_t (SubBytesIns_Inst_Sbox_14_T16), .Z0_t (SubBytesIns_Inst_Sbox_14_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T1), .B0_t (SubBytesIns_Inst_Sbox_14_T12), .Z0_t (SubBytesIns_Inst_Sbox_14_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T13), .B0_t (SubBytesIns_Inst_Sbox_14_T6), .Z0_t (SubBytesIns_Inst_Sbox_14_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T23), .B0_t (SubBytesIns_Inst_Sbox_14_T8), .Z0_t (SubBytesIns_Inst_Sbox_14_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T14), .B0_t (SubBytesIns_Inst_Sbox_14_M1), .Z0_t (SubBytesIns_Inst_Sbox_14_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T19), .B0_t (ciphertext[112]), .Z0_t (SubBytesIns_Inst_Sbox_14_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M4), .B0_t (SubBytesIns_Inst_Sbox_14_M1), .Z0_t (SubBytesIns_Inst_Sbox_14_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T3), .B0_t (SubBytesIns_Inst_Sbox_14_T16), .Z0_t (SubBytesIns_Inst_Sbox_14_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T22), .B0_t (SubBytesIns_Inst_Sbox_14_T9), .Z0_t (SubBytesIns_Inst_Sbox_14_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T26), .B0_t (SubBytesIns_Inst_Sbox_14_M6), .Z0_t (SubBytesIns_Inst_Sbox_14_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T20), .B0_t (SubBytesIns_Inst_Sbox_14_T17), .Z0_t (SubBytesIns_Inst_Sbox_14_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M9), .B0_t (SubBytesIns_Inst_Sbox_14_M6), .Z0_t (SubBytesIns_Inst_Sbox_14_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T1), .B0_t (SubBytesIns_Inst_Sbox_14_T15), .Z0_t (SubBytesIns_Inst_Sbox_14_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T4), .B0_t (SubBytesIns_Inst_Sbox_14_T27), .Z0_t (SubBytesIns_Inst_Sbox_14_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M12), .B0_t (SubBytesIns_Inst_Sbox_14_M11), .Z0_t (SubBytesIns_Inst_Sbox_14_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_T2), .B0_t (SubBytesIns_Inst_Sbox_14_T10), .Z0_t (SubBytesIns_Inst_Sbox_14_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M14), .B0_t (SubBytesIns_Inst_Sbox_14_M11), .Z0_t (SubBytesIns_Inst_Sbox_14_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M3), .B0_t (SubBytesIns_Inst_Sbox_14_M2), .Z0_t (SubBytesIns_Inst_Sbox_14_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M5), .B0_t (SubBytesIns_Inst_Sbox_14_T24), .Z0_t (SubBytesIns_Inst_Sbox_14_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M8), .B0_t (SubBytesIns_Inst_Sbox_14_M7), .Z0_t (SubBytesIns_Inst_Sbox_14_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M10), .B0_t (SubBytesIns_Inst_Sbox_14_M15), .Z0_t (SubBytesIns_Inst_Sbox_14_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M16), .B0_t (SubBytesIns_Inst_Sbox_14_M13), .Z0_t (SubBytesIns_Inst_Sbox_14_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M17), .B0_t (SubBytesIns_Inst_Sbox_14_M15), .Z0_t (SubBytesIns_Inst_Sbox_14_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M18), .B0_t (SubBytesIns_Inst_Sbox_14_M13), .Z0_t (SubBytesIns_Inst_Sbox_14_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M19), .B0_t (SubBytesIns_Inst_Sbox_14_T25), .Z0_t (SubBytesIns_Inst_Sbox_14_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M22), .B0_t (SubBytesIns_Inst_Sbox_14_M23), .Z0_t (SubBytesIns_Inst_Sbox_14_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M22), .B0_t (SubBytesIns_Inst_Sbox_14_M20), .Z0_t (SubBytesIns_Inst_Sbox_14_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M21), .B0_t (SubBytesIns_Inst_Sbox_14_M25), .Z0_t (SubBytesIns_Inst_Sbox_14_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M20), .B0_t (SubBytesIns_Inst_Sbox_14_M21), .Z0_t (SubBytesIns_Inst_Sbox_14_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M23), .B0_t (SubBytesIns_Inst_Sbox_14_M25), .Z0_t (SubBytesIns_Inst_Sbox_14_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M28), .B0_t (SubBytesIns_Inst_Sbox_14_M27), .Z0_t (SubBytesIns_Inst_Sbox_14_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M26), .B0_t (SubBytesIns_Inst_Sbox_14_M24), .Z0_t (SubBytesIns_Inst_Sbox_14_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M20), .B0_t (SubBytesIns_Inst_Sbox_14_M23), .Z0_t (SubBytesIns_Inst_Sbox_14_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M27), .B0_t (SubBytesIns_Inst_Sbox_14_M31), .Z0_t (SubBytesIns_Inst_Sbox_14_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M27), .B0_t (SubBytesIns_Inst_Sbox_14_M25), .Z0_t (SubBytesIns_Inst_Sbox_14_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M21), .B0_t (SubBytesIns_Inst_Sbox_14_M22), .Z0_t (SubBytesIns_Inst_Sbox_14_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M24), .B0_t (SubBytesIns_Inst_Sbox_14_M34), .Z0_t (SubBytesIns_Inst_Sbox_14_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M24), .B0_t (SubBytesIns_Inst_Sbox_14_M25), .Z0_t (SubBytesIns_Inst_Sbox_14_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M21), .B0_t (SubBytesIns_Inst_Sbox_14_M29), .Z0_t (SubBytesIns_Inst_Sbox_14_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M32), .B0_t (SubBytesIns_Inst_Sbox_14_M33), .Z0_t (SubBytesIns_Inst_Sbox_14_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M23), .B0_t (SubBytesIns_Inst_Sbox_14_M30), .Z0_t (SubBytesIns_Inst_Sbox_14_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M35), .B0_t (SubBytesIns_Inst_Sbox_14_M36), .Z0_t (SubBytesIns_Inst_Sbox_14_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M38), .B0_t (SubBytesIns_Inst_Sbox_14_M40), .Z0_t (SubBytesIns_Inst_Sbox_14_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M37), .B0_t (SubBytesIns_Inst_Sbox_14_M39), .Z0_t (SubBytesIns_Inst_Sbox_14_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M37), .B0_t (SubBytesIns_Inst_Sbox_14_M38), .Z0_t (SubBytesIns_Inst_Sbox_14_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M39), .B0_t (SubBytesIns_Inst_Sbox_14_M40), .Z0_t (SubBytesIns_Inst_Sbox_14_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M42), .B0_t (SubBytesIns_Inst_Sbox_14_M41), .Z0_t (SubBytesIns_Inst_Sbox_14_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M44), .B0_t (SubBytesIns_Inst_Sbox_14_T6), .Z0_t (SubBytesIns_Inst_Sbox_14_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M40), .B0_t (SubBytesIns_Inst_Sbox_14_T8), .Z0_t (SubBytesIns_Inst_Sbox_14_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M39), .B0_t (ciphertext[112]), .Z0_t (SubBytesIns_Inst_Sbox_14_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M43), .B0_t (SubBytesIns_Inst_Sbox_14_T16), .Z0_t (SubBytesIns_Inst_Sbox_14_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M38), .B0_t (SubBytesIns_Inst_Sbox_14_T9), .Z0_t (SubBytesIns_Inst_Sbox_14_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M37), .B0_t (SubBytesIns_Inst_Sbox_14_T17), .Z0_t (SubBytesIns_Inst_Sbox_14_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M42), .B0_t (SubBytesIns_Inst_Sbox_14_T15), .Z0_t (SubBytesIns_Inst_Sbox_14_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M45), .B0_t (SubBytesIns_Inst_Sbox_14_T27), .Z0_t (SubBytesIns_Inst_Sbox_14_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M41), .B0_t (SubBytesIns_Inst_Sbox_14_T10), .Z0_t (SubBytesIns_Inst_Sbox_14_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M44), .B0_t (SubBytesIns_Inst_Sbox_14_T13), .Z0_t (SubBytesIns_Inst_Sbox_14_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M40), .B0_t (SubBytesIns_Inst_Sbox_14_T23), .Z0_t (SubBytesIns_Inst_Sbox_14_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M39), .B0_t (SubBytesIns_Inst_Sbox_14_T19), .Z0_t (SubBytesIns_Inst_Sbox_14_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M43), .B0_t (SubBytesIns_Inst_Sbox_14_T3), .Z0_t (SubBytesIns_Inst_Sbox_14_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M38), .B0_t (SubBytesIns_Inst_Sbox_14_T22), .Z0_t (SubBytesIns_Inst_Sbox_14_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M37), .B0_t (SubBytesIns_Inst_Sbox_14_T20), .Z0_t (SubBytesIns_Inst_Sbox_14_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M42), .B0_t (SubBytesIns_Inst_Sbox_14_T1), .Z0_t (SubBytesIns_Inst_Sbox_14_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M45), .B0_t (SubBytesIns_Inst_Sbox_14_T4), .Z0_t (SubBytesIns_Inst_Sbox_14_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M41), .B0_t (SubBytesIns_Inst_Sbox_14_T2), .Z0_t (SubBytesIns_Inst_Sbox_14_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M61), .B0_t (SubBytesIns_Inst_Sbox_14_M62), .Z0_t (SubBytesIns_Inst_Sbox_14_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M50), .B0_t (SubBytesIns_Inst_Sbox_14_M56), .Z0_t (SubBytesIns_Inst_Sbox_14_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M46), .B0_t (SubBytesIns_Inst_Sbox_14_M48), .Z0_t (SubBytesIns_Inst_Sbox_14_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M47), .B0_t (SubBytesIns_Inst_Sbox_14_M55), .Z0_t (SubBytesIns_Inst_Sbox_14_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M54), .B0_t (SubBytesIns_Inst_Sbox_14_M58), .Z0_t (SubBytesIns_Inst_Sbox_14_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M49), .B0_t (SubBytesIns_Inst_Sbox_14_M61), .Z0_t (SubBytesIns_Inst_Sbox_14_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M62), .B0_t (SubBytesIns_Inst_Sbox_14_L5), .Z0_t (SubBytesIns_Inst_Sbox_14_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M46), .B0_t (SubBytesIns_Inst_Sbox_14_L3), .Z0_t (SubBytesIns_Inst_Sbox_14_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M51), .B0_t (SubBytesIns_Inst_Sbox_14_M59), .Z0_t (SubBytesIns_Inst_Sbox_14_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M52), .B0_t (SubBytesIns_Inst_Sbox_14_M53), .Z0_t (SubBytesIns_Inst_Sbox_14_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M53), .B0_t (SubBytesIns_Inst_Sbox_14_L4), .Z0_t (SubBytesIns_Inst_Sbox_14_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M60), .B0_t (SubBytesIns_Inst_Sbox_14_L2), .Z0_t (SubBytesIns_Inst_Sbox_14_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M48), .B0_t (SubBytesIns_Inst_Sbox_14_M51), .Z0_t (SubBytesIns_Inst_Sbox_14_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M50), .B0_t (SubBytesIns_Inst_Sbox_14_L0), .Z0_t (SubBytesIns_Inst_Sbox_14_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M52), .B0_t (SubBytesIns_Inst_Sbox_14_M61), .Z0_t (SubBytesIns_Inst_Sbox_14_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M55), .B0_t (SubBytesIns_Inst_Sbox_14_L1), .Z0_t (SubBytesIns_Inst_Sbox_14_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M56), .B0_t (SubBytesIns_Inst_Sbox_14_L0), .Z0_t (SubBytesIns_Inst_Sbox_14_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M57), .B0_t (SubBytesIns_Inst_Sbox_14_L1), .Z0_t (SubBytesIns_Inst_Sbox_14_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M58), .B0_t (SubBytesIns_Inst_Sbox_14_L8), .Z0_t (SubBytesIns_Inst_Sbox_14_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_M63), .B0_t (SubBytesIns_Inst_Sbox_14_L4), .Z0_t (SubBytesIns_Inst_Sbox_14_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L0), .B0_t (SubBytesIns_Inst_Sbox_14_L1), .Z0_t (SubBytesIns_Inst_Sbox_14_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L1), .B0_t (SubBytesIns_Inst_Sbox_14_L7), .Z0_t (SubBytesIns_Inst_Sbox_14_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L3), .B0_t (SubBytesIns_Inst_Sbox_14_L12), .Z0_t (SubBytesIns_Inst_Sbox_14_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L18), .B0_t (SubBytesIns_Inst_Sbox_14_L2), .Z0_t (SubBytesIns_Inst_Sbox_14_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L15), .B0_t (SubBytesIns_Inst_Sbox_14_L9), .Z0_t (SubBytesIns_Inst_Sbox_14_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L6), .B0_t (SubBytesIns_Inst_Sbox_14_L10), .Z0_t (SubBytesIns_Inst_Sbox_14_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L7), .B0_t (SubBytesIns_Inst_Sbox_14_L9), .Z0_t (SubBytesIns_Inst_Sbox_14_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L8), .B0_t (SubBytesIns_Inst_Sbox_14_L10), .Z0_t (SubBytesIns_Inst_Sbox_14_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L11), .B0_t (SubBytesIns_Inst_Sbox_14_L14), .Z0_t (SubBytesIns_Inst_Sbox_14_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L11), .B0_t (SubBytesIns_Inst_Sbox_14_L17), .Z0_t (SubBytesIns_Inst_Sbox_14_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L6), .B0_t (SubBytesIns_Inst_Sbox_14_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L16), .B0_t (SubBytesIns_Inst_Sbox_14_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L19), .B0_t (SubBytesIns_Inst_Sbox_14_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L6), .B0_t (SubBytesIns_Inst_Sbox_14_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L20), .B0_t (SubBytesIns_Inst_Sbox_14_L22), .Z0_t (MixColumnsInput[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L25), .B0_t (SubBytesIns_Inst_Sbox_14_L29), .Z0_t (MixColumnsInput[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L13), .B0_t (SubBytesIns_Inst_Sbox_14_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_14_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_14_L6), .B0_t (SubBytesIns_Inst_Sbox_14_L23), .Z0_t (MixColumnsInput[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T1_U1 ( .A0_t (ciphertext[127]), .B0_t (ciphertext[124]), .Z0_t (SubBytesIns_Inst_Sbox_15_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T2_U1 ( .A0_t (ciphertext[127]), .B0_t (ciphertext[122]), .Z0_t (SubBytesIns_Inst_Sbox_15_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T3_U1 ( .A0_t (ciphertext[127]), .B0_t (ciphertext[121]), .Z0_t (SubBytesIns_Inst_Sbox_15_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T4_U1 ( .A0_t (ciphertext[124]), .B0_t (ciphertext[122]), .Z0_t (SubBytesIns_Inst_Sbox_15_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T5_U1 ( .A0_t (ciphertext[123]), .B0_t (ciphertext[121]), .Z0_t (SubBytesIns_Inst_Sbox_15_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T1), .B0_t (SubBytesIns_Inst_Sbox_15_T5), .Z0_t (SubBytesIns_Inst_Sbox_15_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T7_U1 ( .A0_t (ciphertext[126]), .B0_t (ciphertext[125]), .Z0_t (SubBytesIns_Inst_Sbox_15_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T8_U1 ( .A0_t (ciphertext[120]), .B0_t (SubBytesIns_Inst_Sbox_15_T6), .Z0_t (SubBytesIns_Inst_Sbox_15_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T9_U1 ( .A0_t (ciphertext[120]), .B0_t (SubBytesIns_Inst_Sbox_15_T7), .Z0_t (SubBytesIns_Inst_Sbox_15_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T6), .B0_t (SubBytesIns_Inst_Sbox_15_T7), .Z0_t (SubBytesIns_Inst_Sbox_15_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T11_U1 ( .A0_t (ciphertext[126]), .B0_t (ciphertext[122]), .Z0_t (SubBytesIns_Inst_Sbox_15_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T12_U1 ( .A0_t (ciphertext[125]), .B0_t (ciphertext[122]), .Z0_t (SubBytesIns_Inst_Sbox_15_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T3), .B0_t (SubBytesIns_Inst_Sbox_15_T4), .Z0_t (SubBytesIns_Inst_Sbox_15_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T6), .B0_t (SubBytesIns_Inst_Sbox_15_T11), .Z0_t (SubBytesIns_Inst_Sbox_15_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T5), .B0_t (SubBytesIns_Inst_Sbox_15_T11), .Z0_t (SubBytesIns_Inst_Sbox_15_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T5), .B0_t (SubBytesIns_Inst_Sbox_15_T12), .Z0_t (SubBytesIns_Inst_Sbox_15_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T9), .B0_t (SubBytesIns_Inst_Sbox_15_T16), .Z0_t (SubBytesIns_Inst_Sbox_15_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T18_U1 ( .A0_t (ciphertext[124]), .B0_t (ciphertext[120]), .Z0_t (SubBytesIns_Inst_Sbox_15_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T7), .B0_t (SubBytesIns_Inst_Sbox_15_T18), .Z0_t (SubBytesIns_Inst_Sbox_15_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T1), .B0_t (SubBytesIns_Inst_Sbox_15_T19), .Z0_t (SubBytesIns_Inst_Sbox_15_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T21_U1 ( .A0_t (ciphertext[121]), .B0_t (ciphertext[120]), .Z0_t (SubBytesIns_Inst_Sbox_15_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T7), .B0_t (SubBytesIns_Inst_Sbox_15_T21), .Z0_t (SubBytesIns_Inst_Sbox_15_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T2), .B0_t (SubBytesIns_Inst_Sbox_15_T22), .Z0_t (SubBytesIns_Inst_Sbox_15_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T2), .B0_t (SubBytesIns_Inst_Sbox_15_T10), .Z0_t (SubBytesIns_Inst_Sbox_15_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T20), .B0_t (SubBytesIns_Inst_Sbox_15_T17), .Z0_t (SubBytesIns_Inst_Sbox_15_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T3), .B0_t (SubBytesIns_Inst_Sbox_15_T16), .Z0_t (SubBytesIns_Inst_Sbox_15_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_T27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T1), .B0_t (SubBytesIns_Inst_Sbox_15_T12), .Z0_t (SubBytesIns_Inst_Sbox_15_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T13), .B0_t (SubBytesIns_Inst_Sbox_15_T6), .Z0_t (SubBytesIns_Inst_Sbox_15_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T23), .B0_t (SubBytesIns_Inst_Sbox_15_T8), .Z0_t (SubBytesIns_Inst_Sbox_15_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T14), .B0_t (SubBytesIns_Inst_Sbox_15_M1), .Z0_t (SubBytesIns_Inst_Sbox_15_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T19), .B0_t (ciphertext[120]), .Z0_t (SubBytesIns_Inst_Sbox_15_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M4), .B0_t (SubBytesIns_Inst_Sbox_15_M1), .Z0_t (SubBytesIns_Inst_Sbox_15_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T3), .B0_t (SubBytesIns_Inst_Sbox_15_T16), .Z0_t (SubBytesIns_Inst_Sbox_15_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T22), .B0_t (SubBytesIns_Inst_Sbox_15_T9), .Z0_t (SubBytesIns_Inst_Sbox_15_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T26), .B0_t (SubBytesIns_Inst_Sbox_15_M6), .Z0_t (SubBytesIns_Inst_Sbox_15_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T20), .B0_t (SubBytesIns_Inst_Sbox_15_T17), .Z0_t (SubBytesIns_Inst_Sbox_15_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M9), .B0_t (SubBytesIns_Inst_Sbox_15_M6), .Z0_t (SubBytesIns_Inst_Sbox_15_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T1), .B0_t (SubBytesIns_Inst_Sbox_15_T15), .Z0_t (SubBytesIns_Inst_Sbox_15_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T4), .B0_t (SubBytesIns_Inst_Sbox_15_T27), .Z0_t (SubBytesIns_Inst_Sbox_15_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M12), .B0_t (SubBytesIns_Inst_Sbox_15_M11), .Z0_t (SubBytesIns_Inst_Sbox_15_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_T2), .B0_t (SubBytesIns_Inst_Sbox_15_T10), .Z0_t (SubBytesIns_Inst_Sbox_15_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M14), .B0_t (SubBytesIns_Inst_Sbox_15_M11), .Z0_t (SubBytesIns_Inst_Sbox_15_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M3), .B0_t (SubBytesIns_Inst_Sbox_15_M2), .Z0_t (SubBytesIns_Inst_Sbox_15_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M5), .B0_t (SubBytesIns_Inst_Sbox_15_T24), .Z0_t (SubBytesIns_Inst_Sbox_15_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M8), .B0_t (SubBytesIns_Inst_Sbox_15_M7), .Z0_t (SubBytesIns_Inst_Sbox_15_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M10), .B0_t (SubBytesIns_Inst_Sbox_15_M15), .Z0_t (SubBytesIns_Inst_Sbox_15_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M16), .B0_t (SubBytesIns_Inst_Sbox_15_M13), .Z0_t (SubBytesIns_Inst_Sbox_15_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M17), .B0_t (SubBytesIns_Inst_Sbox_15_M15), .Z0_t (SubBytesIns_Inst_Sbox_15_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M18), .B0_t (SubBytesIns_Inst_Sbox_15_M13), .Z0_t (SubBytesIns_Inst_Sbox_15_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M19), .B0_t (SubBytesIns_Inst_Sbox_15_T25), .Z0_t (SubBytesIns_Inst_Sbox_15_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M22), .B0_t (SubBytesIns_Inst_Sbox_15_M23), .Z0_t (SubBytesIns_Inst_Sbox_15_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M22), .B0_t (SubBytesIns_Inst_Sbox_15_M20), .Z0_t (SubBytesIns_Inst_Sbox_15_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M21), .B0_t (SubBytesIns_Inst_Sbox_15_M25), .Z0_t (SubBytesIns_Inst_Sbox_15_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M20), .B0_t (SubBytesIns_Inst_Sbox_15_M21), .Z0_t (SubBytesIns_Inst_Sbox_15_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M23), .B0_t (SubBytesIns_Inst_Sbox_15_M25), .Z0_t (SubBytesIns_Inst_Sbox_15_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M28), .B0_t (SubBytesIns_Inst_Sbox_15_M27), .Z0_t (SubBytesIns_Inst_Sbox_15_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M30_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M26), .B0_t (SubBytesIns_Inst_Sbox_15_M24), .Z0_t (SubBytesIns_Inst_Sbox_15_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M31_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M20), .B0_t (SubBytesIns_Inst_Sbox_15_M23), .Z0_t (SubBytesIns_Inst_Sbox_15_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M32_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M27), .B0_t (SubBytesIns_Inst_Sbox_15_M31), .Z0_t (SubBytesIns_Inst_Sbox_15_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M33_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M27), .B0_t (SubBytesIns_Inst_Sbox_15_M25), .Z0_t (SubBytesIns_Inst_Sbox_15_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M34_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M21), .B0_t (SubBytesIns_Inst_Sbox_15_M22), .Z0_t (SubBytesIns_Inst_Sbox_15_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M35_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M24), .B0_t (SubBytesIns_Inst_Sbox_15_M34), .Z0_t (SubBytesIns_Inst_Sbox_15_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M36_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M24), .B0_t (SubBytesIns_Inst_Sbox_15_M25), .Z0_t (SubBytesIns_Inst_Sbox_15_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M37_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M21), .B0_t (SubBytesIns_Inst_Sbox_15_M29), .Z0_t (SubBytesIns_Inst_Sbox_15_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M38_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M32), .B0_t (SubBytesIns_Inst_Sbox_15_M33), .Z0_t (SubBytesIns_Inst_Sbox_15_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M39_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M23), .B0_t (SubBytesIns_Inst_Sbox_15_M30), .Z0_t (SubBytesIns_Inst_Sbox_15_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M40_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M35), .B0_t (SubBytesIns_Inst_Sbox_15_M36), .Z0_t (SubBytesIns_Inst_Sbox_15_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M41_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M38), .B0_t (SubBytesIns_Inst_Sbox_15_M40), .Z0_t (SubBytesIns_Inst_Sbox_15_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M42_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M37), .B0_t (SubBytesIns_Inst_Sbox_15_M39), .Z0_t (SubBytesIns_Inst_Sbox_15_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M43_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M37), .B0_t (SubBytesIns_Inst_Sbox_15_M38), .Z0_t (SubBytesIns_Inst_Sbox_15_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M44_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M39), .B0_t (SubBytesIns_Inst_Sbox_15_M40), .Z0_t (SubBytesIns_Inst_Sbox_15_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_M45_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M42), .B0_t (SubBytesIns_Inst_Sbox_15_M41), .Z0_t (SubBytesIns_Inst_Sbox_15_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M46_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M44), .B0_t (SubBytesIns_Inst_Sbox_15_T6), .Z0_t (SubBytesIns_Inst_Sbox_15_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M47_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M40), .B0_t (SubBytesIns_Inst_Sbox_15_T8), .Z0_t (SubBytesIns_Inst_Sbox_15_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M48_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M39), .B0_t (ciphertext[120]), .Z0_t (SubBytesIns_Inst_Sbox_15_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M49_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M43), .B0_t (SubBytesIns_Inst_Sbox_15_T16), .Z0_t (SubBytesIns_Inst_Sbox_15_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M50_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M38), .B0_t (SubBytesIns_Inst_Sbox_15_T9), .Z0_t (SubBytesIns_Inst_Sbox_15_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M51_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M37), .B0_t (SubBytesIns_Inst_Sbox_15_T17), .Z0_t (SubBytesIns_Inst_Sbox_15_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M52_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M42), .B0_t (SubBytesIns_Inst_Sbox_15_T15), .Z0_t (SubBytesIns_Inst_Sbox_15_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M53_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M45), .B0_t (SubBytesIns_Inst_Sbox_15_T27), .Z0_t (SubBytesIns_Inst_Sbox_15_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M54_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M41), .B0_t (SubBytesIns_Inst_Sbox_15_T10), .Z0_t (SubBytesIns_Inst_Sbox_15_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M55_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M44), .B0_t (SubBytesIns_Inst_Sbox_15_T13), .Z0_t (SubBytesIns_Inst_Sbox_15_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M56_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M40), .B0_t (SubBytesIns_Inst_Sbox_15_T23), .Z0_t (SubBytesIns_Inst_Sbox_15_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M57_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M39), .B0_t (SubBytesIns_Inst_Sbox_15_T19), .Z0_t (SubBytesIns_Inst_Sbox_15_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M58_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M43), .B0_t (SubBytesIns_Inst_Sbox_15_T3), .Z0_t (SubBytesIns_Inst_Sbox_15_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M59_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M38), .B0_t (SubBytesIns_Inst_Sbox_15_T22), .Z0_t (SubBytesIns_Inst_Sbox_15_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M60_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M37), .B0_t (SubBytesIns_Inst_Sbox_15_T20), .Z0_t (SubBytesIns_Inst_Sbox_15_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M61_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M42), .B0_t (SubBytesIns_Inst_Sbox_15_T1), .Z0_t (SubBytesIns_Inst_Sbox_15_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M62_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M45), .B0_t (SubBytesIns_Inst_Sbox_15_T4), .Z0_t (SubBytesIns_Inst_Sbox_15_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_AND_M63_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M41), .B0_t (SubBytesIns_Inst_Sbox_15_T2), .Z0_t (SubBytesIns_Inst_Sbox_15_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M61), .B0_t (SubBytesIns_Inst_Sbox_15_M62), .Z0_t (SubBytesIns_Inst_Sbox_15_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M50), .B0_t (SubBytesIns_Inst_Sbox_15_M56), .Z0_t (SubBytesIns_Inst_Sbox_15_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M46), .B0_t (SubBytesIns_Inst_Sbox_15_M48), .Z0_t (SubBytesIns_Inst_Sbox_15_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M47), .B0_t (SubBytesIns_Inst_Sbox_15_M55), .Z0_t (SubBytesIns_Inst_Sbox_15_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M54), .B0_t (SubBytesIns_Inst_Sbox_15_M58), .Z0_t (SubBytesIns_Inst_Sbox_15_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M49), .B0_t (SubBytesIns_Inst_Sbox_15_M61), .Z0_t (SubBytesIns_Inst_Sbox_15_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M62), .B0_t (SubBytesIns_Inst_Sbox_15_L5), .Z0_t (SubBytesIns_Inst_Sbox_15_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M46), .B0_t (SubBytesIns_Inst_Sbox_15_L3), .Z0_t (SubBytesIns_Inst_Sbox_15_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L8_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M51), .B0_t (SubBytesIns_Inst_Sbox_15_M59), .Z0_t (SubBytesIns_Inst_Sbox_15_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L9_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M52), .B0_t (SubBytesIns_Inst_Sbox_15_M53), .Z0_t (SubBytesIns_Inst_Sbox_15_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L10_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M53), .B0_t (SubBytesIns_Inst_Sbox_15_L4), .Z0_t (SubBytesIns_Inst_Sbox_15_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L11_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M60), .B0_t (SubBytesIns_Inst_Sbox_15_L2), .Z0_t (SubBytesIns_Inst_Sbox_15_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L12_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M48), .B0_t (SubBytesIns_Inst_Sbox_15_M51), .Z0_t (SubBytesIns_Inst_Sbox_15_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L13_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M50), .B0_t (SubBytesIns_Inst_Sbox_15_L0), .Z0_t (SubBytesIns_Inst_Sbox_15_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L14_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M52), .B0_t (SubBytesIns_Inst_Sbox_15_M61), .Z0_t (SubBytesIns_Inst_Sbox_15_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L15_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M55), .B0_t (SubBytesIns_Inst_Sbox_15_L1), .Z0_t (SubBytesIns_Inst_Sbox_15_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L16_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M56), .B0_t (SubBytesIns_Inst_Sbox_15_L0), .Z0_t (SubBytesIns_Inst_Sbox_15_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L17_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M57), .B0_t (SubBytesIns_Inst_Sbox_15_L1), .Z0_t (SubBytesIns_Inst_Sbox_15_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L18_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M58), .B0_t (SubBytesIns_Inst_Sbox_15_L8), .Z0_t (SubBytesIns_Inst_Sbox_15_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L19_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_M63), .B0_t (SubBytesIns_Inst_Sbox_15_L4), .Z0_t (SubBytesIns_Inst_Sbox_15_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L20_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L0), .B0_t (SubBytesIns_Inst_Sbox_15_L1), .Z0_t (SubBytesIns_Inst_Sbox_15_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L21_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L1), .B0_t (SubBytesIns_Inst_Sbox_15_L7), .Z0_t (SubBytesIns_Inst_Sbox_15_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L22_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L3), .B0_t (SubBytesIns_Inst_Sbox_15_L12), .Z0_t (SubBytesIns_Inst_Sbox_15_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L23_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L18), .B0_t (SubBytesIns_Inst_Sbox_15_L2), .Z0_t (SubBytesIns_Inst_Sbox_15_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L24_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L15), .B0_t (SubBytesIns_Inst_Sbox_15_L9), .Z0_t (SubBytesIns_Inst_Sbox_15_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L25_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L6), .B0_t (SubBytesIns_Inst_Sbox_15_L10), .Z0_t (SubBytesIns_Inst_Sbox_15_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L26_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L7), .B0_t (SubBytesIns_Inst_Sbox_15_L9), .Z0_t (SubBytesIns_Inst_Sbox_15_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L27_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L8), .B0_t (SubBytesIns_Inst_Sbox_15_L10), .Z0_t (SubBytesIns_Inst_Sbox_15_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L28_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L11), .B0_t (SubBytesIns_Inst_Sbox_15_L14), .Z0_t (SubBytesIns_Inst_Sbox_15_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_L29_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L11), .B0_t (SubBytesIns_Inst_Sbox_15_L17), .Z0_t (SubBytesIns_Inst_Sbox_15_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S0_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L6), .B0_t (SubBytesIns_Inst_Sbox_15_L24), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S1_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L16), .B0_t (SubBytesIns_Inst_Sbox_15_L26), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S2_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L19), .B0_t (SubBytesIns_Inst_Sbox_15_L28), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S3_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L6), .B0_t (SubBytesIns_Inst_Sbox_15_L21), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S4_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L20), .B0_t (SubBytesIns_Inst_Sbox_15_L22), .Z0_t (MixColumnsInput[123]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S5_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L25), .B0_t (SubBytesIns_Inst_Sbox_15_L29), .Z0_t (MixColumnsInput[122]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S6_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L13), .B0_t (SubBytesIns_Inst_Sbox_15_L27), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubBytesIns_Inst_Sbox_15_XOR_S7_U1 ( .A0_t (SubBytesIns_Inst_Sbox_15_L6), .B0_t (SubBytesIns_Inst_Sbox_15_L23), .Z0_t (MixColumnsInput[120]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U96 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n192), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .Z0_t (MixColumnsOutput[105]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U95 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n191), .B0_t (MixColumnsIns_MixOneColumnInst_0_n190), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U94 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n189), .B0_t (MixColumnsIns_MixOneColumnInst_0_n188), .Z0_t (MixColumnsOutput[104]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U93 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n187), .B0_t (MixColumnsInput[112]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U92 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n186), .B0_t (MixColumnsIns_MixOneColumnInst_0_n185), .Z0_t (MixColumnsOutput[103]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U91 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n184), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U90 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n183), .B0_t (MixColumnsIns_MixOneColumnInst_0_n182), .Z0_t (MixColumnsOutput[102]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U89 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n181), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U88 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n180), .B0_t (MixColumnsIns_MixOneColumnInst_0_n179), .Z0_t (MixColumnsOutput[101]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U87 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n178), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U86 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n177), .B0_t (MixColumnsIns_MixOneColumnInst_0_n176), .Z0_t (MixColumnsOutput[100]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U85 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n175), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U84 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n174), .B0_t (MixColumnsIns_MixOneColumnInst_0_n173), .Z0_t (MixColumnsOutput[99]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U83 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n172), .B0_t (MixColumnsInput[107]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U82 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n171), .B0_t (MixColumnsIns_MixOneColumnInst_0_n185), .Z0_t (MixColumnsOutput[127]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U81 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U80 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n170), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U79 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n169), .B0_t (MixColumnsIns_MixOneColumnInst_0_n182), .Z0_t (MixColumnsOutput[126]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U78 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U77 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n168), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U76 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n167), .B0_t (MixColumnsIns_MixOneColumnInst_0_n166), .Z0_t (MixColumnsOutput[98]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U75 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n165), .B0_t (MixColumnsInput[106]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U74 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n164), .B0_t (MixColumnsIns_MixOneColumnInst_0_n179), .Z0_t (MixColumnsOutput[125]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U73 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U72 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n163), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U71 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n162), .B0_t (MixColumnsIns_MixOneColumnInst_0_n176), .Z0_t (MixColumnsOutput[124]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U70 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U69 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n161), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U68 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n160), .B0_t (MixColumnsIns_MixOneColumnInst_0_n173), .Z0_t (MixColumnsOutput[123]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U67 ( .A0_t (MixColumnsInput[115]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U66 ( .A0_t (MixColumnsInput[99]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n159), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U65 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n158), .B0_t (MixColumnsIns_MixOneColumnInst_0_n166), .Z0_t (MixColumnsOutput[122]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U64 ( .A0_t (MixColumnsInput[114]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U63 ( .A0_t (MixColumnsInput[98]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n157), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U62 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n156), .B0_t (MixColumnsIns_MixOneColumnInst_0_n155), .Z0_t (MixColumnsOutput[121]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U61 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n154), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U60 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n153), .B0_t (MixColumnsIns_MixOneColumnInst_0_n152), .Z0_t (MixColumnsOutput[120]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U59 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n151), .B0_t (MixColumnsInput[96]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U58 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n150), .B0_t (MixColumnsIns_MixOneColumnInst_0_n170), .Z0_t (MixColumnsOutput[119]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U57 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U56 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n149), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U55 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n148), .B0_t (MixColumnsIns_MixOneColumnInst_0_n168), .Z0_t (MixColumnsOutput[118]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U54 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U53 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n147), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U52 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n146), .B0_t (MixColumnsIns_MixOneColumnInst_0_n163), .Z0_t (MixColumnsOutput[117]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U51 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U50 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n145), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U49 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n144), .B0_t (MixColumnsIns_MixOneColumnInst_0_n161), .Z0_t (MixColumnsOutput[116]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U48 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U47 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n143), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U46 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n142), .B0_t (MixColumnsIns_MixOneColumnInst_0_n155), .Z0_t (MixColumnsOutput[97]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U45 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U44 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n190), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U43 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U42 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n141), .B0_t (MixColumnsIns_MixOneColumnInst_0_n159), .Z0_t (MixColumnsOutput[115]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U41 ( .A0_t (MixColumnsInput[107]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U40 ( .A0_t (MixColumnsInput[123]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n140), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U39 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n139), .B0_t (MixColumnsIns_MixOneColumnInst_0_n157), .Z0_t (MixColumnsOutput[114]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U38 ( .A0_t (MixColumnsInput[106]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U37 ( .A0_t (MixColumnsInput[122]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n138), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U36 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n137), .B0_t (MixColumnsIns_MixOneColumnInst_0_n154), .Z0_t (MixColumnsOutput[113]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U35 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U34 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n191), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U33 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U32 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n136), .B0_t (MixColumnsIns_MixOneColumnInst_0_n152), .Z0_t (MixColumnsOutput[112]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U31 ( .A0_t (MixColumnsInput[104]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U30 ( .A0_t (MixColumnsInput[120]), .B0_t (MixColumnsIns_MixOneColumnInst_0_n188), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U29 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B0_t (MixColumnsInput[96]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n188) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U28 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n135), .B0_t (MixColumnsIns_MixOneColumnInst_0_n149), .Z0_t (MixColumnsOutput[111]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U27 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U26 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n184), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U25 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U24 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n134), .B0_t (MixColumnsIns_MixOneColumnInst_0_n147), .Z0_t (MixColumnsOutput[110]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U23 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U22 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n181), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U21 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U20 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n133), .B0_t (MixColumnsIns_MixOneColumnInst_0_n145), .Z0_t (MixColumnsOutput[109]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U19 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U18 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n178), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U17 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U16 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n132), .B0_t (MixColumnsIns_MixOneColumnInst_0_n143), .Z0_t (MixColumnsOutput[108]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U15 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U14 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n175), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U13 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U12 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n131), .B0_t (MixColumnsIns_MixOneColumnInst_0_n140), .Z0_t (MixColumnsOutput[107]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U11 ( .A0_t (MixColumnsInput[99]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U10 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n172), .B0_t (MixColumnsInput[115]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U9 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]), .B0_t (MixColumnsInput[123]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U8 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n130), .B0_t (MixColumnsIns_MixOneColumnInst_0_n138), .Z0_t (MixColumnsOutput[106]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U7 ( .A0_t (MixColumnsInput[98]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U6 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n165), .B0_t (MixColumnsInput[114]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U5 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .B0_t (MixColumnsInput[122]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n129), .B0_t (MixColumnsInput[104]), .Z0_t (MixColumnsOutput[96]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_n187), .B0_t (MixColumnsIns_MixOneColumnInst_0_n151), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U2 ( .A0_t (MixColumnsInput[112]), .B0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_U1 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B0_t (MixColumnsInput[120]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_n187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B0_t (MixColumnsInput[123]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B0_t (MixColumnsInput[122]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B0_t (MixColumnsInput[120]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B0_t (MixColumnsInput[115]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B0_t (MixColumnsInput[114]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B0_t (MixColumnsInput[112]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B0_t (MixColumnsInput[107]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B0_t (MixColumnsInput[106]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B0_t (MixColumnsInput[104]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B0_t (MixColumnsInput[99]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B0_t (MixColumnsInput[98]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B0_t (MixColumnsInput[96]), .Z0_t (MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U96 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n192), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .Z0_t (MixColumnsOutput[73]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U95 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n191), .B0_t (MixColumnsIns_MixOneColumnInst_1_n190), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U94 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n189), .B0_t (MixColumnsIns_MixOneColumnInst_1_n188), .Z0_t (MixColumnsOutput[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U93 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n187), .B0_t (MixColumnsInput[80]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U92 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n186), .B0_t (MixColumnsIns_MixOneColumnInst_1_n185), .Z0_t (MixColumnsOutput[71]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U91 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n184), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U90 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n183), .B0_t (MixColumnsIns_MixOneColumnInst_1_n182), .Z0_t (MixColumnsOutput[70]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U89 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n181), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U88 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n180), .B0_t (MixColumnsIns_MixOneColumnInst_1_n179), .Z0_t (MixColumnsOutput[69]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U87 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n178), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U86 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n177), .B0_t (MixColumnsIns_MixOneColumnInst_1_n176), .Z0_t (MixColumnsOutput[68]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U85 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n175), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U84 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n174), .B0_t (MixColumnsIns_MixOneColumnInst_1_n173), .Z0_t (MixColumnsOutput[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U83 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n172), .B0_t (MixColumnsInput[75]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U82 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n171), .B0_t (MixColumnsIns_MixOneColumnInst_1_n185), .Z0_t (MixColumnsOutput[95]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U81 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U80 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n170), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U79 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n169), .B0_t (MixColumnsIns_MixOneColumnInst_1_n182), .Z0_t (MixColumnsOutput[94]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U78 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U77 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n168), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U76 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n167), .B0_t (MixColumnsIns_MixOneColumnInst_1_n166), .Z0_t (MixColumnsOutput[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U75 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n165), .B0_t (MixColumnsInput[74]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U74 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n164), .B0_t (MixColumnsIns_MixOneColumnInst_1_n179), .Z0_t (MixColumnsOutput[93]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U73 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U72 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n163), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U71 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n162), .B0_t (MixColumnsIns_MixOneColumnInst_1_n176), .Z0_t (MixColumnsOutput[92]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U70 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U69 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n161), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U68 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n160), .B0_t (MixColumnsIns_MixOneColumnInst_1_n173), .Z0_t (MixColumnsOutput[91]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U67 ( .A0_t (MixColumnsInput[83]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U66 ( .A0_t (MixColumnsInput[67]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n159), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U65 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n158), .B0_t (MixColumnsIns_MixOneColumnInst_1_n166), .Z0_t (MixColumnsOutput[90]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U64 ( .A0_t (MixColumnsInput[82]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U63 ( .A0_t (MixColumnsInput[66]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n157), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U62 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n156), .B0_t (MixColumnsIns_MixOneColumnInst_1_n155), .Z0_t (MixColumnsOutput[89]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U61 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n154), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U60 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n153), .B0_t (MixColumnsIns_MixOneColumnInst_1_n152), .Z0_t (MixColumnsOutput[88]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U59 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n151), .B0_t (MixColumnsInput[64]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U58 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n150), .B0_t (MixColumnsIns_MixOneColumnInst_1_n170), .Z0_t (MixColumnsOutput[87]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U57 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U56 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n149), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U55 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n148), .B0_t (MixColumnsIns_MixOneColumnInst_1_n168), .Z0_t (MixColumnsOutput[86]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U54 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U53 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n147), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U52 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n146), .B0_t (MixColumnsIns_MixOneColumnInst_1_n163), .Z0_t (MixColumnsOutput[85]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U51 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U50 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n145), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U49 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n144), .B0_t (MixColumnsIns_MixOneColumnInst_1_n161), .Z0_t (MixColumnsOutput[84]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U48 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U47 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n143), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U46 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n142), .B0_t (MixColumnsIns_MixOneColumnInst_1_n155), .Z0_t (MixColumnsOutput[65]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U45 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U44 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n190), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U43 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U42 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n141), .B0_t (MixColumnsIns_MixOneColumnInst_1_n159), .Z0_t (MixColumnsOutput[83]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U41 ( .A0_t (MixColumnsInput[75]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U40 ( .A0_t (MixColumnsInput[91]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n140), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U39 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n139), .B0_t (MixColumnsIns_MixOneColumnInst_1_n157), .Z0_t (MixColumnsOutput[82]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U38 ( .A0_t (MixColumnsInput[74]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U37 ( .A0_t (MixColumnsInput[90]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n138), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U36 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n137), .B0_t (MixColumnsIns_MixOneColumnInst_1_n154), .Z0_t (MixColumnsOutput[81]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U35 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U34 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n191), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U33 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U32 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n136), .B0_t (MixColumnsIns_MixOneColumnInst_1_n152), .Z0_t (MixColumnsOutput[80]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U31 ( .A0_t (MixColumnsInput[72]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U30 ( .A0_t (MixColumnsInput[88]), .B0_t (MixColumnsIns_MixOneColumnInst_1_n188), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U29 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B0_t (MixColumnsInput[64]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n188) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U28 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n135), .B0_t (MixColumnsIns_MixOneColumnInst_1_n149), .Z0_t (MixColumnsOutput[79]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U27 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U26 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n184), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U25 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U24 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n134), .B0_t (MixColumnsIns_MixOneColumnInst_1_n147), .Z0_t (MixColumnsOutput[78]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U23 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U22 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n181), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U21 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U20 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n133), .B0_t (MixColumnsIns_MixOneColumnInst_1_n145), .Z0_t (MixColumnsOutput[77]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U19 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U18 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n178), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U17 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U16 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n132), .B0_t (MixColumnsIns_MixOneColumnInst_1_n143), .Z0_t (MixColumnsOutput[76]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U15 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U14 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n175), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U13 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U12 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n131), .B0_t (MixColumnsIns_MixOneColumnInst_1_n140), .Z0_t (MixColumnsOutput[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U11 ( .A0_t (MixColumnsInput[67]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U10 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n172), .B0_t (MixColumnsInput[83]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U9 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]), .B0_t (MixColumnsInput[91]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U8 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n130), .B0_t (MixColumnsIns_MixOneColumnInst_1_n138), .Z0_t (MixColumnsOutput[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U7 ( .A0_t (MixColumnsInput[66]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U6 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n165), .B0_t (MixColumnsInput[82]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U5 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .B0_t (MixColumnsInput[90]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n129), .B0_t (MixColumnsInput[72]), .Z0_t (MixColumnsOutput[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_n187), .B0_t (MixColumnsIns_MixOneColumnInst_1_n151), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U2 ( .A0_t (MixColumnsInput[80]), .B0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_U1 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B0_t (MixColumnsInput[88]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_n187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B0_t (MixColumnsInput[91]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B0_t (MixColumnsInput[90]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B0_t (MixColumnsInput[88]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B0_t (MixColumnsInput[83]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B0_t (MixColumnsInput[82]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B0_t (MixColumnsInput[80]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B0_t (MixColumnsInput[75]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B0_t (MixColumnsInput[74]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B0_t (MixColumnsInput[72]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B0_t (MixColumnsInput[67]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B0_t (MixColumnsInput[66]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B0_t (MixColumnsInput[64]), .Z0_t (MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U96 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n192), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .Z0_t (MixColumnsOutput[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U95 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n191), .B0_t (MixColumnsIns_MixOneColumnInst_2_n190), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U94 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n189), .B0_t (MixColumnsIns_MixOneColumnInst_2_n188), .Z0_t (MixColumnsOutput[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U93 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n187), .B0_t (MixColumnsInput[48]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U92 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n186), .B0_t (MixColumnsIns_MixOneColumnInst_2_n185), .Z0_t (MixColumnsOutput[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U91 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n184), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U90 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n183), .B0_t (MixColumnsIns_MixOneColumnInst_2_n182), .Z0_t (MixColumnsOutput[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U89 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n181), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U88 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n180), .B0_t (MixColumnsIns_MixOneColumnInst_2_n179), .Z0_t (MixColumnsOutput[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U87 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n178), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U86 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n177), .B0_t (MixColumnsIns_MixOneColumnInst_2_n176), .Z0_t (MixColumnsOutput[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U85 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n175), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U84 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n174), .B0_t (MixColumnsIns_MixOneColumnInst_2_n173), .Z0_t (MixColumnsOutput[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U83 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n172), .B0_t (MixColumnsInput[43]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U82 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n171), .B0_t (MixColumnsIns_MixOneColumnInst_2_n185), .Z0_t (MixColumnsOutput[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U81 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U80 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n170), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U79 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n169), .B0_t (MixColumnsIns_MixOneColumnInst_2_n182), .Z0_t (MixColumnsOutput[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U78 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U77 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n168), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U76 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n167), .B0_t (MixColumnsIns_MixOneColumnInst_2_n166), .Z0_t (MixColumnsOutput[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U75 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n165), .B0_t (MixColumnsInput[42]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U74 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n164), .B0_t (MixColumnsIns_MixOneColumnInst_2_n179), .Z0_t (MixColumnsOutput[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U73 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U72 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n163), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U71 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n162), .B0_t (MixColumnsIns_MixOneColumnInst_2_n176), .Z0_t (MixColumnsOutput[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U70 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U69 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n161), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U68 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n160), .B0_t (MixColumnsIns_MixOneColumnInst_2_n173), .Z0_t (MixColumnsOutput[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U67 ( .A0_t (MixColumnsInput[51]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U66 ( .A0_t (MixColumnsInput[35]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n159), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U65 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n158), .B0_t (MixColumnsIns_MixOneColumnInst_2_n166), .Z0_t (MixColumnsOutput[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U64 ( .A0_t (MixColumnsInput[50]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U63 ( .A0_t (MixColumnsInput[34]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n157), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U62 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n156), .B0_t (MixColumnsIns_MixOneColumnInst_2_n155), .Z0_t (MixColumnsOutput[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U61 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n154), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U60 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n153), .B0_t (MixColumnsIns_MixOneColumnInst_2_n152), .Z0_t (MixColumnsOutput[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U59 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n151), .B0_t (MixColumnsInput[32]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U58 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n150), .B0_t (MixColumnsIns_MixOneColumnInst_2_n170), .Z0_t (MixColumnsOutput[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U57 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U56 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n149), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U55 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n148), .B0_t (MixColumnsIns_MixOneColumnInst_2_n168), .Z0_t (MixColumnsOutput[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U54 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U53 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n147), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U52 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n146), .B0_t (MixColumnsIns_MixOneColumnInst_2_n163), .Z0_t (MixColumnsOutput[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U51 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U50 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n145), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U49 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n144), .B0_t (MixColumnsIns_MixOneColumnInst_2_n161), .Z0_t (MixColumnsOutput[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U48 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U47 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n143), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U46 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n142), .B0_t (MixColumnsIns_MixOneColumnInst_2_n155), .Z0_t (MixColumnsOutput[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U45 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U44 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n190), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U43 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U42 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n141), .B0_t (MixColumnsIns_MixOneColumnInst_2_n159), .Z0_t (MixColumnsOutput[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U41 ( .A0_t (MixColumnsInput[43]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U40 ( .A0_t (MixColumnsInput[59]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n140), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U39 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n139), .B0_t (MixColumnsIns_MixOneColumnInst_2_n157), .Z0_t (MixColumnsOutput[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U38 ( .A0_t (MixColumnsInput[42]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U37 ( .A0_t (MixColumnsInput[58]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n138), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U36 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n137), .B0_t (MixColumnsIns_MixOneColumnInst_2_n154), .Z0_t (MixColumnsOutput[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U35 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U34 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n191), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U33 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U32 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n136), .B0_t (MixColumnsIns_MixOneColumnInst_2_n152), .Z0_t (MixColumnsOutput[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U31 ( .A0_t (MixColumnsInput[40]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U30 ( .A0_t (MixColumnsInput[56]), .B0_t (MixColumnsIns_MixOneColumnInst_2_n188), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U29 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B0_t (MixColumnsInput[32]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n188) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U28 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n135), .B0_t (MixColumnsIns_MixOneColumnInst_2_n149), .Z0_t (MixColumnsOutput[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U27 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U26 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n184), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U25 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U24 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n134), .B0_t (MixColumnsIns_MixOneColumnInst_2_n147), .Z0_t (MixColumnsOutput[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U23 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U22 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n181), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U21 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U20 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n133), .B0_t (MixColumnsIns_MixOneColumnInst_2_n145), .Z0_t (MixColumnsOutput[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U19 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U18 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n178), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U17 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U16 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n132), .B0_t (MixColumnsIns_MixOneColumnInst_2_n143), .Z0_t (MixColumnsOutput[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U15 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U14 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n175), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U13 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U12 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n131), .B0_t (MixColumnsIns_MixOneColumnInst_2_n140), .Z0_t (MixColumnsOutput[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U11 ( .A0_t (MixColumnsInput[35]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U10 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n172), .B0_t (MixColumnsInput[51]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U9 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]), .B0_t (MixColumnsInput[59]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U8 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n130), .B0_t (MixColumnsIns_MixOneColumnInst_2_n138), .Z0_t (MixColumnsOutput[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U7 ( .A0_t (MixColumnsInput[34]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U6 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n165), .B0_t (MixColumnsInput[50]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U5 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .B0_t (MixColumnsInput[58]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n129), .B0_t (MixColumnsInput[40]), .Z0_t (MixColumnsOutput[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_n187), .B0_t (MixColumnsIns_MixOneColumnInst_2_n151), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U2 ( .A0_t (MixColumnsInput[48]), .B0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_U1 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B0_t (MixColumnsInput[56]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_n187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B0_t (MixColumnsInput[59]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B0_t (MixColumnsInput[58]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B0_t (MixColumnsInput[56]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B0_t (MixColumnsInput[51]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B0_t (MixColumnsInput[50]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B0_t (MixColumnsInput[48]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B0_t (MixColumnsInput[43]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B0_t (MixColumnsInput[42]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B0_t (MixColumnsInput[40]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B0_t (MixColumnsInput[35]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B0_t (MixColumnsInput[34]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B0_t (MixColumnsInput[32]), .Z0_t (MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U96 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n192), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .Z0_t (MixColumnsOutput[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U95 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n191), .B0_t (MixColumnsIns_MixOneColumnInst_3_n190), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U94 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n189), .B0_t (MixColumnsIns_MixOneColumnInst_3_n188), .Z0_t (MixColumnsOutput[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U93 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n187), .B0_t (MixColumnsInput[16]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U92 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n186), .B0_t (MixColumnsIns_MixOneColumnInst_3_n185), .Z0_t (MixColumnsOutput[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U91 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n184), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U90 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n183), .B0_t (MixColumnsIns_MixOneColumnInst_3_n182), .Z0_t (MixColumnsOutput[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U89 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n181), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U88 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n180), .B0_t (MixColumnsIns_MixOneColumnInst_3_n179), .Z0_t (MixColumnsOutput[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U87 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n178), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U86 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n177), .B0_t (MixColumnsIns_MixOneColumnInst_3_n176), .Z0_t (MixColumnsOutput[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U85 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n175), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U84 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n174), .B0_t (MixColumnsIns_MixOneColumnInst_3_n173), .Z0_t (MixColumnsOutput[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U83 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n172), .B0_t (MixColumnsInput[11]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U82 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n171), .B0_t (MixColumnsIns_MixOneColumnInst_3_n185), .Z0_t (MixColumnsOutput[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U81 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U80 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n170), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U79 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n169), .B0_t (MixColumnsIns_MixOneColumnInst_3_n182), .Z0_t (MixColumnsOutput[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U78 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U77 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n168), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U76 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n167), .B0_t (MixColumnsIns_MixOneColumnInst_3_n166), .Z0_t (MixColumnsOutput[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U75 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n165), .B0_t (MixColumnsInput[10]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U74 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n164), .B0_t (MixColumnsIns_MixOneColumnInst_3_n179), .Z0_t (MixColumnsOutput[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U73 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U72 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n163), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U71 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n162), .B0_t (MixColumnsIns_MixOneColumnInst_3_n176), .Z0_t (MixColumnsOutput[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U70 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U69 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n161), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U68 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n160), .B0_t (MixColumnsIns_MixOneColumnInst_3_n173), .Z0_t (MixColumnsOutput[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U67 ( .A0_t (MixColumnsInput[19]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U66 ( .A0_t (MixColumnsInput[3]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n159), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U65 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n158), .B0_t (MixColumnsIns_MixOneColumnInst_3_n166), .Z0_t (MixColumnsOutput[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U64 ( .A0_t (MixColumnsInput[18]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U63 ( .A0_t (MixColumnsInput[2]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n157), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U62 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n156), .B0_t (MixColumnsIns_MixOneColumnInst_3_n155), .Z0_t (MixColumnsOutput[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U61 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n154), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U60 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n153), .B0_t (MixColumnsIns_MixOneColumnInst_3_n152), .Z0_t (MixColumnsOutput[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U59 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n151), .B0_t (MixColumnsInput[0]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U58 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n150), .B0_t (MixColumnsIns_MixOneColumnInst_3_n170), .Z0_t (MixColumnsOutput[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U57 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U56 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n149), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U55 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n148), .B0_t (MixColumnsIns_MixOneColumnInst_3_n168), .Z0_t (MixColumnsOutput[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U54 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U53 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n147), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U52 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n146), .B0_t (MixColumnsIns_MixOneColumnInst_3_n163), .Z0_t (MixColumnsOutput[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U51 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U50 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n145), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U49 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n144), .B0_t (MixColumnsIns_MixOneColumnInst_3_n161), .Z0_t (MixColumnsOutput[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U48 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U47 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n143), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U46 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n142), .B0_t (MixColumnsIns_MixOneColumnInst_3_n155), .Z0_t (MixColumnsOutput[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U45 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U44 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n190), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U43 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U42 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n141), .B0_t (MixColumnsIns_MixOneColumnInst_3_n159), .Z0_t (MixColumnsOutput[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U41 ( .A0_t (MixColumnsInput[11]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U40 ( .A0_t (MixColumnsInput[27]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n140), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U39 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n139), .B0_t (MixColumnsIns_MixOneColumnInst_3_n157), .Z0_t (MixColumnsOutput[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U38 ( .A0_t (MixColumnsInput[10]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U37 ( .A0_t (MixColumnsInput[26]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n138), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U36 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n137), .B0_t (MixColumnsIns_MixOneColumnInst_3_n154), .Z0_t (MixColumnsOutput[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U35 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U34 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n191), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U33 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U32 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n136), .B0_t (MixColumnsIns_MixOneColumnInst_3_n152), .Z0_t (MixColumnsOutput[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U31 ( .A0_t (MixColumnsInput[8]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U30 ( .A0_t (MixColumnsInput[24]), .B0_t (MixColumnsIns_MixOneColumnInst_3_n188), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U29 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B0_t (MixColumnsInput[0]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n188) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U28 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n135), .B0_t (MixColumnsIns_MixOneColumnInst_3_n149), .Z0_t (MixColumnsOutput[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U27 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U26 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n184), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U25 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U24 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n134), .B0_t (MixColumnsIns_MixOneColumnInst_3_n147), .Z0_t (MixColumnsOutput[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U23 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U22 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n181), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U21 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U20 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n133), .B0_t (MixColumnsIns_MixOneColumnInst_3_n145), .Z0_t (MixColumnsOutput[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U19 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U18 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n178), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U17 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U16 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n132), .B0_t (MixColumnsIns_MixOneColumnInst_3_n143), .Z0_t (MixColumnsOutput[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U15 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U14 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n175), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U13 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U12 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n131), .B0_t (MixColumnsIns_MixOneColumnInst_3_n140), .Z0_t (MixColumnsOutput[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U11 ( .A0_t (MixColumnsInput[3]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U10 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n172), .B0_t (MixColumnsInput[19]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U9 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]), .B0_t (MixColumnsInput[27]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U8 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n130), .B0_t (MixColumnsIns_MixOneColumnInst_3_n138), .Z0_t (MixColumnsOutput[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U7 ( .A0_t (MixColumnsInput[2]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U6 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n165), .B0_t (MixColumnsInput[18]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U5 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .B0_t (MixColumnsInput[26]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n129), .B0_t (MixColumnsInput[8]), .Z0_t (MixColumnsOutput[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_n187), .B0_t (MixColumnsIns_MixOneColumnInst_3_n151), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U2 ( .A0_t (MixColumnsInput[16]), .B0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_U1 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B0_t (MixColumnsInput[24]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_n187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B0_t (MixColumnsInput[27]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B0_t (MixColumnsInput[26]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B0_t (MixColumnsInput[24]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B0_t (MixColumnsInput[19]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B0_t (MixColumnsInput[18]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B0_t (MixColumnsInput[16]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B0_t (MixColumnsInput[11]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B0_t (MixColumnsInput[10]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B0_t (MixColumnsInput[8]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U4 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B0_t (MixColumnsInput[3]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U3 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B0_t (MixColumnsInput[2]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U2 ( .A0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B0_t (MixColumnsInput[0]), .Z0_t (MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_0_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[0]), .B0_t (key[0]), .Z0_t (KeyReg_Inst_ff_SDE_0_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_0_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_0_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_0_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_0_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_0_MUX_inst_Y), .B0_t (KeyExpansionOutput[0]), .Z0_t (RoundKey[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_1_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[1]), .B0_t (key[1]), .Z0_t (KeyReg_Inst_ff_SDE_1_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_1_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_1_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_1_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_1_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_1_MUX_inst_Y), .B0_t (KeyExpansionOutput[1]), .Z0_t (RoundKey[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_2_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[2]), .B0_t (key[2]), .Z0_t (KeyReg_Inst_ff_SDE_2_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_2_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_2_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_2_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_2_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_2_MUX_inst_Y), .B0_t (KeyExpansionOutput[2]), .Z0_t (RoundKey[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_3_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[3]), .B0_t (key[3]), .Z0_t (KeyReg_Inst_ff_SDE_3_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_3_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_3_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_3_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_3_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_3_MUX_inst_Y), .B0_t (KeyExpansionOutput[3]), .Z0_t (RoundKey[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_4_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[4]), .B0_t (key[4]), .Z0_t (KeyReg_Inst_ff_SDE_4_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_4_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_4_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_4_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_4_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_4_MUX_inst_Y), .B0_t (KeyExpansionOutput[4]), .Z0_t (RoundKey[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_5_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[5]), .B0_t (key[5]), .Z0_t (KeyReg_Inst_ff_SDE_5_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_5_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_5_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_5_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_5_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_5_MUX_inst_Y), .B0_t (KeyExpansionOutput[5]), .Z0_t (RoundKey[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_6_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[6]), .B0_t (key[6]), .Z0_t (KeyReg_Inst_ff_SDE_6_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_6_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_6_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_6_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_6_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_6_MUX_inst_Y), .B0_t (KeyExpansionOutput[6]), .Z0_t (RoundKey[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_7_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[7]), .B0_t (key[7]), .Z0_t (KeyReg_Inst_ff_SDE_7_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_7_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_7_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_7_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_7_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_7_MUX_inst_Y), .B0_t (KeyExpansionOutput[7]), .Z0_t (RoundKey[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_8_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[8]), .B0_t (key[8]), .Z0_t (KeyReg_Inst_ff_SDE_8_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_8_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_8_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_8_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_8_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_8_MUX_inst_Y), .B0_t (KeyExpansionOutput[8]), .Z0_t (RoundKey[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_9_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[9]), .B0_t (key[9]), .Z0_t (KeyReg_Inst_ff_SDE_9_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_9_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_9_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_9_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_9_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_9_MUX_inst_Y), .B0_t (KeyExpansionOutput[9]), .Z0_t (RoundKey[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_10_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[10]), .B0_t (key[10]), .Z0_t (KeyReg_Inst_ff_SDE_10_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_10_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_10_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_10_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_10_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_10_MUX_inst_Y), .B0_t (KeyExpansionOutput[10]), .Z0_t (RoundKey[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_11_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[11]), .B0_t (key[11]), .Z0_t (KeyReg_Inst_ff_SDE_11_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_11_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_11_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_11_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_11_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_11_MUX_inst_Y), .B0_t (KeyExpansionOutput[11]), .Z0_t (RoundKey[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_12_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[12]), .B0_t (key[12]), .Z0_t (KeyReg_Inst_ff_SDE_12_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_12_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_12_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_12_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_12_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_12_MUX_inst_Y), .B0_t (KeyExpansionOutput[12]), .Z0_t (RoundKey[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_13_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[13]), .B0_t (key[13]), .Z0_t (KeyReg_Inst_ff_SDE_13_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_13_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_13_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_13_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_13_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_13_MUX_inst_Y), .B0_t (KeyExpansionOutput[13]), .Z0_t (RoundKey[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_14_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[14]), .B0_t (key[14]), .Z0_t (KeyReg_Inst_ff_SDE_14_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_14_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_14_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_14_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_14_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_14_MUX_inst_Y), .B0_t (KeyExpansionOutput[14]), .Z0_t (RoundKey[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_15_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[15]), .B0_t (key[15]), .Z0_t (KeyReg_Inst_ff_SDE_15_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_15_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_15_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_15_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_15_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_15_MUX_inst_Y), .B0_t (KeyExpansionOutput[15]), .Z0_t (RoundKey[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_16_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[16]), .B0_t (key[16]), .Z0_t (KeyReg_Inst_ff_SDE_16_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_16_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_16_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_16_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_16_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_16_MUX_inst_Y), .B0_t (KeyExpansionOutput[16]), .Z0_t (RoundKey[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_17_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[17]), .B0_t (key[17]), .Z0_t (KeyReg_Inst_ff_SDE_17_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_17_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_17_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_17_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_17_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_17_MUX_inst_Y), .B0_t (KeyExpansionOutput[17]), .Z0_t (RoundKey[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_18_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[18]), .B0_t (key[18]), .Z0_t (KeyReg_Inst_ff_SDE_18_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_18_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_18_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_18_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_18_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_18_MUX_inst_Y), .B0_t (KeyExpansionOutput[18]), .Z0_t (RoundKey[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_19_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[19]), .B0_t (key[19]), .Z0_t (KeyReg_Inst_ff_SDE_19_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_19_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_19_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_19_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_19_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_19_MUX_inst_Y), .B0_t (KeyExpansionOutput[19]), .Z0_t (RoundKey[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_20_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[20]), .B0_t (key[20]), .Z0_t (KeyReg_Inst_ff_SDE_20_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_20_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_20_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_20_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_20_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_20_MUX_inst_Y), .B0_t (KeyExpansionOutput[20]), .Z0_t (RoundKey[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_21_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[21]), .B0_t (key[21]), .Z0_t (KeyReg_Inst_ff_SDE_21_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_21_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_21_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_21_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_21_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_21_MUX_inst_Y), .B0_t (KeyExpansionOutput[21]), .Z0_t (RoundKey[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_22_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[22]), .B0_t (key[22]), .Z0_t (KeyReg_Inst_ff_SDE_22_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_22_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_22_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_22_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_22_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_22_MUX_inst_Y), .B0_t (KeyExpansionOutput[22]), .Z0_t (RoundKey[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_23_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[23]), .B0_t (key[23]), .Z0_t (KeyReg_Inst_ff_SDE_23_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_23_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_23_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_23_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_23_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_23_MUX_inst_Y), .B0_t (KeyExpansionOutput[23]), .Z0_t (RoundKey[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_24_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[24]), .B0_t (key[24]), .Z0_t (KeyReg_Inst_ff_SDE_24_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_24_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_24_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_24_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_24_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_24_MUX_inst_Y), .B0_t (KeyExpansionOutput[24]), .Z0_t (RoundKey[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_25_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[25]), .B0_t (key[25]), .Z0_t (KeyReg_Inst_ff_SDE_25_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_25_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_25_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_25_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_25_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_25_MUX_inst_Y), .B0_t (KeyExpansionOutput[25]), .Z0_t (RoundKey[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_26_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[26]), .B0_t (key[26]), .Z0_t (KeyReg_Inst_ff_SDE_26_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_26_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_26_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_26_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_26_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_26_MUX_inst_Y), .B0_t (KeyExpansionOutput[26]), .Z0_t (RoundKey[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_27_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[27]), .B0_t (key[27]), .Z0_t (KeyReg_Inst_ff_SDE_27_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_27_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_27_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_27_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_27_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_27_MUX_inst_Y), .B0_t (KeyExpansionOutput[27]), .Z0_t (RoundKey[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_28_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[28]), .B0_t (key[28]), .Z0_t (KeyReg_Inst_ff_SDE_28_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_28_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_28_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_28_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_28_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_28_MUX_inst_Y), .B0_t (KeyExpansionOutput[28]), .Z0_t (RoundKey[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_29_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[29]), .B0_t (key[29]), .Z0_t (KeyReg_Inst_ff_SDE_29_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_29_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_29_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_29_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_29_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_29_MUX_inst_Y), .B0_t (KeyExpansionOutput[29]), .Z0_t (RoundKey[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_30_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[30]), .B0_t (key[30]), .Z0_t (KeyReg_Inst_ff_SDE_30_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_30_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_30_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_30_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_30_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_30_MUX_inst_Y), .B0_t (KeyExpansionOutput[30]), .Z0_t (RoundKey[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_31_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[31]), .B0_t (key[31]), .Z0_t (KeyReg_Inst_ff_SDE_31_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_31_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_31_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_31_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_31_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_31_MUX_inst_Y), .B0_t (KeyExpansionOutput[31]), .Z0_t (RoundKey[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_32_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[32]), .B0_t (key[32]), .Z0_t (KeyReg_Inst_ff_SDE_32_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_32_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_32_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_32_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_32_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_32_MUX_inst_Y), .B0_t (KeyExpansionOutput[32]), .Z0_t (RoundKey[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_33_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[33]), .B0_t (key[33]), .Z0_t (KeyReg_Inst_ff_SDE_33_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_33_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_33_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_33_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_33_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_33_MUX_inst_Y), .B0_t (KeyExpansionOutput[33]), .Z0_t (RoundKey[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_34_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[34]), .B0_t (key[34]), .Z0_t (KeyReg_Inst_ff_SDE_34_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_34_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_34_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_34_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_34_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_34_MUX_inst_Y), .B0_t (KeyExpansionOutput[34]), .Z0_t (RoundKey[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_35_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[35]), .B0_t (key[35]), .Z0_t (KeyReg_Inst_ff_SDE_35_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_35_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_35_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_35_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_35_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_35_MUX_inst_Y), .B0_t (KeyExpansionOutput[35]), .Z0_t (RoundKey[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_36_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[36]), .B0_t (key[36]), .Z0_t (KeyReg_Inst_ff_SDE_36_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_36_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_36_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_36_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_36_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_36_MUX_inst_Y), .B0_t (KeyExpansionOutput[36]), .Z0_t (RoundKey[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_37_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[37]), .B0_t (key[37]), .Z0_t (KeyReg_Inst_ff_SDE_37_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_37_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_37_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_37_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_37_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_37_MUX_inst_Y), .B0_t (KeyExpansionOutput[37]), .Z0_t (RoundKey[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_38_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[38]), .B0_t (key[38]), .Z0_t (KeyReg_Inst_ff_SDE_38_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_38_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_38_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_38_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_38_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_38_MUX_inst_Y), .B0_t (KeyExpansionOutput[38]), .Z0_t (RoundKey[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_39_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[39]), .B0_t (key[39]), .Z0_t (KeyReg_Inst_ff_SDE_39_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_39_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_39_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_39_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_39_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_39_MUX_inst_Y), .B0_t (KeyExpansionOutput[39]), .Z0_t (RoundKey[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_40_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[40]), .B0_t (key[40]), .Z0_t (KeyReg_Inst_ff_SDE_40_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_40_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_40_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_40_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_40_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_40_MUX_inst_Y), .B0_t (KeyExpansionOutput[40]), .Z0_t (RoundKey[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_41_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[41]), .B0_t (key[41]), .Z0_t (KeyReg_Inst_ff_SDE_41_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_41_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_41_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_41_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_41_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_41_MUX_inst_Y), .B0_t (KeyExpansionOutput[41]), .Z0_t (RoundKey[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_42_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[42]), .B0_t (key[42]), .Z0_t (KeyReg_Inst_ff_SDE_42_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_42_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_42_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_42_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_42_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_42_MUX_inst_Y), .B0_t (KeyExpansionOutput[42]), .Z0_t (RoundKey[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_43_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[43]), .B0_t (key[43]), .Z0_t (KeyReg_Inst_ff_SDE_43_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_43_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_43_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_43_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_43_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_43_MUX_inst_Y), .B0_t (KeyExpansionOutput[43]), .Z0_t (RoundKey[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_44_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[44]), .B0_t (key[44]), .Z0_t (KeyReg_Inst_ff_SDE_44_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_44_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_44_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_44_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_44_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_44_MUX_inst_Y), .B0_t (KeyExpansionOutput[44]), .Z0_t (RoundKey[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_45_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[45]), .B0_t (key[45]), .Z0_t (KeyReg_Inst_ff_SDE_45_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_45_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_45_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_45_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_45_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_45_MUX_inst_Y), .B0_t (KeyExpansionOutput[45]), .Z0_t (RoundKey[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_46_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[46]), .B0_t (key[46]), .Z0_t (KeyReg_Inst_ff_SDE_46_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_46_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_46_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_46_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_46_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_46_MUX_inst_Y), .B0_t (KeyExpansionOutput[46]), .Z0_t (RoundKey[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_47_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[47]), .B0_t (key[47]), .Z0_t (KeyReg_Inst_ff_SDE_47_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_47_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_47_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_47_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_47_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_47_MUX_inst_Y), .B0_t (KeyExpansionOutput[47]), .Z0_t (RoundKey[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_48_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[48]), .B0_t (key[48]), .Z0_t (KeyReg_Inst_ff_SDE_48_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_48_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_48_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_48_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_48_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_48_MUX_inst_Y), .B0_t (KeyExpansionOutput[48]), .Z0_t (RoundKey[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_49_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[49]), .B0_t (key[49]), .Z0_t (KeyReg_Inst_ff_SDE_49_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_49_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_49_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_49_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_49_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_49_MUX_inst_Y), .B0_t (KeyExpansionOutput[49]), .Z0_t (RoundKey[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_50_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[50]), .B0_t (key[50]), .Z0_t (KeyReg_Inst_ff_SDE_50_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_50_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_50_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_50_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_50_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_50_MUX_inst_Y), .B0_t (KeyExpansionOutput[50]), .Z0_t (RoundKey[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_51_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[51]), .B0_t (key[51]), .Z0_t (KeyReg_Inst_ff_SDE_51_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_51_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_51_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_51_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_51_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_51_MUX_inst_Y), .B0_t (KeyExpansionOutput[51]), .Z0_t (RoundKey[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_52_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[52]), .B0_t (key[52]), .Z0_t (KeyReg_Inst_ff_SDE_52_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_52_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_52_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_52_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_52_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_52_MUX_inst_Y), .B0_t (KeyExpansionOutput[52]), .Z0_t (RoundKey[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_53_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[53]), .B0_t (key[53]), .Z0_t (KeyReg_Inst_ff_SDE_53_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_53_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_53_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_53_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_53_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_53_MUX_inst_Y), .B0_t (KeyExpansionOutput[53]), .Z0_t (RoundKey[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_54_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[54]), .B0_t (key[54]), .Z0_t (KeyReg_Inst_ff_SDE_54_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_54_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_54_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_54_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_54_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_54_MUX_inst_Y), .B0_t (KeyExpansionOutput[54]), .Z0_t (RoundKey[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_55_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[55]), .B0_t (key[55]), .Z0_t (KeyReg_Inst_ff_SDE_55_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_55_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_55_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_55_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_55_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_55_MUX_inst_Y), .B0_t (KeyExpansionOutput[55]), .Z0_t (RoundKey[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_56_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[56]), .B0_t (key[56]), .Z0_t (KeyReg_Inst_ff_SDE_56_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_56_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_56_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_56_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_56_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_56_MUX_inst_Y), .B0_t (KeyExpansionOutput[56]), .Z0_t (RoundKey[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_57_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[57]), .B0_t (key[57]), .Z0_t (KeyReg_Inst_ff_SDE_57_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_57_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_57_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_57_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_57_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_57_MUX_inst_Y), .B0_t (KeyExpansionOutput[57]), .Z0_t (RoundKey[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_58_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[58]), .B0_t (key[58]), .Z0_t (KeyReg_Inst_ff_SDE_58_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_58_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_58_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_58_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_58_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_58_MUX_inst_Y), .B0_t (KeyExpansionOutput[58]), .Z0_t (RoundKey[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_59_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[59]), .B0_t (key[59]), .Z0_t (KeyReg_Inst_ff_SDE_59_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_59_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_59_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_59_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_59_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_59_MUX_inst_Y), .B0_t (KeyExpansionOutput[59]), .Z0_t (RoundKey[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_60_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[60]), .B0_t (key[60]), .Z0_t (KeyReg_Inst_ff_SDE_60_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_60_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_60_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_60_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_60_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_60_MUX_inst_Y), .B0_t (KeyExpansionOutput[60]), .Z0_t (RoundKey[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_61_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[61]), .B0_t (key[61]), .Z0_t (KeyReg_Inst_ff_SDE_61_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_61_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_61_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_61_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_61_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_61_MUX_inst_Y), .B0_t (KeyExpansionOutput[61]), .Z0_t (RoundKey[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_62_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[62]), .B0_t (key[62]), .Z0_t (KeyReg_Inst_ff_SDE_62_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_62_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_62_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_62_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_62_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_62_MUX_inst_Y), .B0_t (KeyExpansionOutput[62]), .Z0_t (RoundKey[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_63_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[63]), .B0_t (key[63]), .Z0_t (KeyReg_Inst_ff_SDE_63_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_63_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_63_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_63_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_63_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_63_MUX_inst_Y), .B0_t (KeyExpansionOutput[63]), .Z0_t (RoundKey[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_64_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[64]), .B0_t (key[64]), .Z0_t (KeyReg_Inst_ff_SDE_64_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_64_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_64_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_64_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_64_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_64_MUX_inst_Y), .B0_t (KeyExpansionOutput[64]), .Z0_t (RoundKey[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_65_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[65]), .B0_t (key[65]), .Z0_t (KeyReg_Inst_ff_SDE_65_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_65_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_65_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_65_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_65_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_65_MUX_inst_Y), .B0_t (KeyExpansionOutput[65]), .Z0_t (RoundKey[65]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_66_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[66]), .B0_t (key[66]), .Z0_t (KeyReg_Inst_ff_SDE_66_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_66_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_66_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_66_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_66_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_66_MUX_inst_Y), .B0_t (KeyExpansionOutput[66]), .Z0_t (RoundKey[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_67_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[67]), .B0_t (key[67]), .Z0_t (KeyReg_Inst_ff_SDE_67_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_67_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_67_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_67_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_67_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_67_MUX_inst_Y), .B0_t (KeyExpansionOutput[67]), .Z0_t (RoundKey[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_68_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[68]), .B0_t (key[68]), .Z0_t (KeyReg_Inst_ff_SDE_68_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_68_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_68_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_68_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_68_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_68_MUX_inst_Y), .B0_t (KeyExpansionOutput[68]), .Z0_t (RoundKey[68]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_69_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[69]), .B0_t (key[69]), .Z0_t (KeyReg_Inst_ff_SDE_69_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_69_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_69_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_69_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_69_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_69_MUX_inst_Y), .B0_t (KeyExpansionOutput[69]), .Z0_t (RoundKey[69]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_70_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[70]), .B0_t (key[70]), .Z0_t (KeyReg_Inst_ff_SDE_70_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_70_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_70_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_70_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_70_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_70_MUX_inst_Y), .B0_t (KeyExpansionOutput[70]), .Z0_t (RoundKey[70]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_71_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[71]), .B0_t (key[71]), .Z0_t (KeyReg_Inst_ff_SDE_71_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_71_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_71_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_71_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_71_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_71_MUX_inst_Y), .B0_t (KeyExpansionOutput[71]), .Z0_t (RoundKey[71]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_72_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[72]), .B0_t (key[72]), .Z0_t (KeyReg_Inst_ff_SDE_72_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_72_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_72_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_72_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_72_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_72_MUX_inst_Y), .B0_t (KeyExpansionOutput[72]), .Z0_t (RoundKey[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_73_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[73]), .B0_t (key[73]), .Z0_t (KeyReg_Inst_ff_SDE_73_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_73_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_73_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_73_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_73_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_73_MUX_inst_Y), .B0_t (KeyExpansionOutput[73]), .Z0_t (RoundKey[73]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_74_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[74]), .B0_t (key[74]), .Z0_t (KeyReg_Inst_ff_SDE_74_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_74_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_74_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_74_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_74_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_74_MUX_inst_Y), .B0_t (KeyExpansionOutput[74]), .Z0_t (RoundKey[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_75_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[75]), .B0_t (key[75]), .Z0_t (KeyReg_Inst_ff_SDE_75_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_75_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_75_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_75_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_75_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_75_MUX_inst_Y), .B0_t (KeyExpansionOutput[75]), .Z0_t (RoundKey[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_76_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[76]), .B0_t (key[76]), .Z0_t (KeyReg_Inst_ff_SDE_76_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_76_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_76_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_76_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_76_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_76_MUX_inst_Y), .B0_t (KeyExpansionOutput[76]), .Z0_t (RoundKey[76]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_77_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[77]), .B0_t (key[77]), .Z0_t (KeyReg_Inst_ff_SDE_77_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_77_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_77_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_77_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_77_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_77_MUX_inst_Y), .B0_t (KeyExpansionOutput[77]), .Z0_t (RoundKey[77]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_78_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[78]), .B0_t (key[78]), .Z0_t (KeyReg_Inst_ff_SDE_78_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_78_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_78_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_78_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_78_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_78_MUX_inst_Y), .B0_t (KeyExpansionOutput[78]), .Z0_t (RoundKey[78]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_79_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[79]), .B0_t (key[79]), .Z0_t (KeyReg_Inst_ff_SDE_79_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_79_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_79_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_79_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_79_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_79_MUX_inst_Y), .B0_t (KeyExpansionOutput[79]), .Z0_t (RoundKey[79]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_80_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[80]), .B0_t (key[80]), .Z0_t (KeyReg_Inst_ff_SDE_80_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_80_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_80_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_80_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_80_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_80_MUX_inst_Y), .B0_t (KeyExpansionOutput[80]), .Z0_t (RoundKey[80]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_81_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[81]), .B0_t (key[81]), .Z0_t (KeyReg_Inst_ff_SDE_81_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_81_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_81_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_81_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_81_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_81_MUX_inst_Y), .B0_t (KeyExpansionOutput[81]), .Z0_t (RoundKey[81]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_82_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[82]), .B0_t (key[82]), .Z0_t (KeyReg_Inst_ff_SDE_82_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_82_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_82_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_82_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_82_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_82_MUX_inst_Y), .B0_t (KeyExpansionOutput[82]), .Z0_t (RoundKey[82]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_83_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[83]), .B0_t (key[83]), .Z0_t (KeyReg_Inst_ff_SDE_83_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_83_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_83_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_83_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_83_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_83_MUX_inst_Y), .B0_t (KeyExpansionOutput[83]), .Z0_t (RoundKey[83]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_84_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[84]), .B0_t (key[84]), .Z0_t (KeyReg_Inst_ff_SDE_84_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_84_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_84_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_84_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_84_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_84_MUX_inst_Y), .B0_t (KeyExpansionOutput[84]), .Z0_t (RoundKey[84]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_85_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[85]), .B0_t (key[85]), .Z0_t (KeyReg_Inst_ff_SDE_85_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_85_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_85_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_85_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_85_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_85_MUX_inst_Y), .B0_t (KeyExpansionOutput[85]), .Z0_t (RoundKey[85]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_86_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[86]), .B0_t (key[86]), .Z0_t (KeyReg_Inst_ff_SDE_86_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_86_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_86_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_86_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_86_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_86_MUX_inst_Y), .B0_t (KeyExpansionOutput[86]), .Z0_t (RoundKey[86]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_87_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[87]), .B0_t (key[87]), .Z0_t (KeyReg_Inst_ff_SDE_87_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_87_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_87_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_87_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_87_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_87_MUX_inst_Y), .B0_t (KeyExpansionOutput[87]), .Z0_t (RoundKey[87]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_88_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[88]), .B0_t (key[88]), .Z0_t (KeyReg_Inst_ff_SDE_88_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_88_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_88_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_88_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_88_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_88_MUX_inst_Y), .B0_t (KeyExpansionOutput[88]), .Z0_t (RoundKey[88]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_89_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[89]), .B0_t (key[89]), .Z0_t (KeyReg_Inst_ff_SDE_89_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_89_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_89_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_89_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_89_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_89_MUX_inst_Y), .B0_t (KeyExpansionOutput[89]), .Z0_t (RoundKey[89]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_90_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[90]), .B0_t (key[90]), .Z0_t (KeyReg_Inst_ff_SDE_90_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_90_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_90_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_90_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_90_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_90_MUX_inst_Y), .B0_t (KeyExpansionOutput[90]), .Z0_t (RoundKey[90]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_91_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[91]), .B0_t (key[91]), .Z0_t (KeyReg_Inst_ff_SDE_91_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_91_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_91_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_91_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_91_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_91_MUX_inst_Y), .B0_t (KeyExpansionOutput[91]), .Z0_t (RoundKey[91]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_92_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[92]), .B0_t (key[92]), .Z0_t (KeyReg_Inst_ff_SDE_92_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_92_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_92_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_92_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_92_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_92_MUX_inst_Y), .B0_t (KeyExpansionOutput[92]), .Z0_t (RoundKey[92]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_93_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[93]), .B0_t (key[93]), .Z0_t (KeyReg_Inst_ff_SDE_93_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_93_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_93_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_93_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_93_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_93_MUX_inst_Y), .B0_t (KeyExpansionOutput[93]), .Z0_t (RoundKey[93]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_94_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[94]), .B0_t (key[94]), .Z0_t (KeyReg_Inst_ff_SDE_94_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_94_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_94_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_94_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_94_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_94_MUX_inst_Y), .B0_t (KeyExpansionOutput[94]), .Z0_t (RoundKey[94]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_95_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[95]), .B0_t (key[95]), .Z0_t (KeyReg_Inst_ff_SDE_95_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_95_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_95_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_95_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_95_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_95_MUX_inst_Y), .B0_t (KeyExpansionOutput[95]), .Z0_t (RoundKey[95]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_96_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[96]), .B0_t (key[96]), .Z0_t (KeyReg_Inst_ff_SDE_96_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_96_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_96_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_96_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_96_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_96_MUX_inst_Y), .B0_t (KeyExpansionOutput[96]), .Z0_t (RoundKey[96]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_97_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[97]), .B0_t (key[97]), .Z0_t (KeyReg_Inst_ff_SDE_97_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_97_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_97_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_97_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_97_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_97_MUX_inst_Y), .B0_t (KeyExpansionOutput[97]), .Z0_t (RoundKey[97]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_98_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[98]), .B0_t (key[98]), .Z0_t (KeyReg_Inst_ff_SDE_98_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_98_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_98_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_98_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_98_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_98_MUX_inst_Y), .B0_t (KeyExpansionOutput[98]), .Z0_t (RoundKey[98]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_99_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[99]), .B0_t (key[99]), .Z0_t (KeyReg_Inst_ff_SDE_99_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_99_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_99_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_99_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_99_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_99_MUX_inst_Y), .B0_t (KeyExpansionOutput[99]), .Z0_t (RoundKey[99]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_100_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[100]), .B0_t (key[100]), .Z0_t (KeyReg_Inst_ff_SDE_100_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_100_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_100_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_100_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_100_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_100_MUX_inst_Y), .B0_t (KeyExpansionOutput[100]), .Z0_t (RoundKey[100]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_101_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[101]), .B0_t (key[101]), .Z0_t (KeyReg_Inst_ff_SDE_101_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_101_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_101_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_101_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_101_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_101_MUX_inst_Y), .B0_t (KeyExpansionOutput[101]), .Z0_t (RoundKey[101]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_102_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[102]), .B0_t (key[102]), .Z0_t (KeyReg_Inst_ff_SDE_102_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_102_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_102_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_102_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_102_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_102_MUX_inst_Y), .B0_t (KeyExpansionOutput[102]), .Z0_t (RoundKey[102]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_103_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[103]), .B0_t (key[103]), .Z0_t (KeyReg_Inst_ff_SDE_103_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_103_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_103_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_103_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_103_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_103_MUX_inst_Y), .B0_t (KeyExpansionOutput[103]), .Z0_t (RoundKey[103]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_104_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[104]), .B0_t (key[104]), .Z0_t (KeyReg_Inst_ff_SDE_104_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_104_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_104_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_104_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_104_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_104_MUX_inst_Y), .B0_t (KeyExpansionOutput[104]), .Z0_t (RoundKey[104]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_105_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[105]), .B0_t (key[105]), .Z0_t (KeyReg_Inst_ff_SDE_105_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_105_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_105_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_105_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_105_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_105_MUX_inst_Y), .B0_t (KeyExpansionOutput[105]), .Z0_t (RoundKey[105]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_106_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[106]), .B0_t (key[106]), .Z0_t (KeyReg_Inst_ff_SDE_106_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_106_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_106_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_106_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_106_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_106_MUX_inst_Y), .B0_t (KeyExpansionOutput[106]), .Z0_t (RoundKey[106]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_107_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[107]), .B0_t (key[107]), .Z0_t (KeyReg_Inst_ff_SDE_107_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_107_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_107_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_107_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_107_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_107_MUX_inst_Y), .B0_t (KeyExpansionOutput[107]), .Z0_t (RoundKey[107]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_108_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[108]), .B0_t (key[108]), .Z0_t (KeyReg_Inst_ff_SDE_108_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_108_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_108_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_108_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_108_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_108_MUX_inst_Y), .B0_t (KeyExpansionOutput[108]), .Z0_t (RoundKey[108]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_109_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[109]), .B0_t (key[109]), .Z0_t (KeyReg_Inst_ff_SDE_109_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_109_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_109_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_109_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_109_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_109_MUX_inst_Y), .B0_t (KeyExpansionOutput[109]), .Z0_t (RoundKey[109]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_110_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[110]), .B0_t (key[110]), .Z0_t (KeyReg_Inst_ff_SDE_110_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_110_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_110_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_110_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_110_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_110_MUX_inst_Y), .B0_t (KeyExpansionOutput[110]), .Z0_t (RoundKey[110]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_111_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[111]), .B0_t (key[111]), .Z0_t (KeyReg_Inst_ff_SDE_111_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_111_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_111_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_111_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_111_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_111_MUX_inst_Y), .B0_t (KeyExpansionOutput[111]), .Z0_t (RoundKey[111]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_112_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[112]), .B0_t (key[112]), .Z0_t (KeyReg_Inst_ff_SDE_112_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_112_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_112_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_112_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_112_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_112_MUX_inst_Y), .B0_t (KeyExpansionOutput[112]), .Z0_t (RoundKey[112]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_113_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[113]), .B0_t (key[113]), .Z0_t (KeyReg_Inst_ff_SDE_113_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_113_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_113_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_113_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_113_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_113_MUX_inst_Y), .B0_t (KeyExpansionOutput[113]), .Z0_t (RoundKey[113]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_114_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[114]), .B0_t (key[114]), .Z0_t (KeyReg_Inst_ff_SDE_114_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_114_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_114_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_114_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_114_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_114_MUX_inst_Y), .B0_t (KeyExpansionOutput[114]), .Z0_t (RoundKey[114]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_115_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[115]), .B0_t (key[115]), .Z0_t (KeyReg_Inst_ff_SDE_115_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_115_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_115_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_115_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_115_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_115_MUX_inst_Y), .B0_t (KeyExpansionOutput[115]), .Z0_t (RoundKey[115]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_116_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[116]), .B0_t (key[116]), .Z0_t (KeyReg_Inst_ff_SDE_116_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_116_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_116_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_116_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_116_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_116_MUX_inst_Y), .B0_t (KeyExpansionOutput[116]), .Z0_t (RoundKey[116]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_117_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[117]), .B0_t (key[117]), .Z0_t (KeyReg_Inst_ff_SDE_117_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_117_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_117_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_117_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_117_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_117_MUX_inst_Y), .B0_t (KeyExpansionOutput[117]), .Z0_t (RoundKey[117]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_118_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[118]), .B0_t (key[118]), .Z0_t (KeyReg_Inst_ff_SDE_118_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_118_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_118_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_118_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_118_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_118_MUX_inst_Y), .B0_t (KeyExpansionOutput[118]), .Z0_t (RoundKey[118]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_119_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[119]), .B0_t (key[119]), .Z0_t (KeyReg_Inst_ff_SDE_119_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_119_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_119_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_119_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_119_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_119_MUX_inst_Y), .B0_t (KeyExpansionOutput[119]), .Z0_t (RoundKey[119]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_120_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[120]), .B0_t (key[120]), .Z0_t (KeyReg_Inst_ff_SDE_120_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_120_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_120_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_120_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_120_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_120_MUX_inst_Y), .B0_t (KeyExpansionOutput[120]), .Z0_t (RoundKey[120]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_121_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[121]), .B0_t (key[121]), .Z0_t (KeyReg_Inst_ff_SDE_121_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_121_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_121_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_121_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_121_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_121_MUX_inst_Y), .B0_t (KeyExpansionOutput[121]), .Z0_t (RoundKey[121]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_122_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[122]), .B0_t (key[122]), .Z0_t (KeyReg_Inst_ff_SDE_122_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_122_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_122_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_122_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_122_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_122_MUX_inst_Y), .B0_t (KeyExpansionOutput[122]), .Z0_t (RoundKey[122]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_123_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[123]), .B0_t (key[123]), .Z0_t (KeyReg_Inst_ff_SDE_123_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_123_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_123_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_123_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_123_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_123_MUX_inst_Y), .B0_t (KeyExpansionOutput[123]), .Z0_t (RoundKey[123]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_124_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[124]), .B0_t (key[124]), .Z0_t (KeyReg_Inst_ff_SDE_124_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_124_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_124_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_124_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_124_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_124_MUX_inst_Y), .B0_t (KeyExpansionOutput[124]), .Z0_t (RoundKey[124]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_125_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[125]), .B0_t (key[125]), .Z0_t (KeyReg_Inst_ff_SDE_125_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_125_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_125_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_125_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_125_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_125_MUX_inst_Y), .B0_t (KeyExpansionOutput[125]), .Z0_t (RoundKey[125]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_126_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[126]), .B0_t (key[126]), .Z0_t (KeyReg_Inst_ff_SDE_126_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_126_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_126_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_126_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_126_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_126_MUX_inst_Y), .B0_t (KeyExpansionOutput[126]), .Z0_t (RoundKey[126]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_127_MUX_inst_XOR1_U1 ( .A0_t (KeyExpansionOutput[127]), .B0_t (key[127]), .Z0_t (KeyReg_Inst_ff_SDE_127_MUX_inst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyReg_Inst_ff_SDE_127_MUX_inst_AND1_U1 ( .A0_t (start), .B0_t (KeyReg_Inst_ff_SDE_127_MUX_inst_X), .Z0_t (KeyReg_Inst_ff_SDE_127_MUX_inst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) KeyReg_Inst_ff_SDE_127_MUX_inst_XOR2_U1 ( .A0_t (KeyReg_Inst_ff_SDE_127_MUX_inst_Y), .B0_t (KeyExpansionOutput[127]), .Z0_t (RoundKey[127]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U128 ( .A0_t (RoundKey[9]), .B0_t (KeyExpansionOutput[41]), .Z0_t (KeyExpansionOutput[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U127 ( .A0_t (RoundKey[8]), .B0_t (KeyExpansionOutput[40]), .Z0_t (KeyExpansionOutput[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U126 ( .A0_t (RoundKey[7]), .B0_t (KeyExpansionOutput[39]), .Z0_t (KeyExpansionOutput[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U125 ( .A0_t (RoundKey[6]), .B0_t (KeyExpansionOutput[38]), .Z0_t (KeyExpansionOutput[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U124 ( .A0_t (RoundKey[5]), .B0_t (KeyExpansionOutput[37]), .Z0_t (KeyExpansionOutput[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U123 ( .A0_t (RoundKey[4]), .B0_t (KeyExpansionOutput[36]), .Z0_t (KeyExpansionOutput[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U122 ( .A0_t (RoundKey[41]), .B0_t (KeyExpansionOutput[73]), .Z0_t (KeyExpansionOutput[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U121 ( .A0_t (RoundKey[73]), .B0_t (KeyExpansionOutput[105]), .Z0_t (KeyExpansionOutput[73]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U120 ( .A0_t (RoundKey[40]), .B0_t (KeyExpansionOutput[72]), .Z0_t (KeyExpansionOutput[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U119 ( .A0_t (RoundKey[72]), .B0_t (KeyExpansionOutput[104]), .Z0_t (KeyExpansionOutput[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U118 ( .A0_t (RoundKey[3]), .B0_t (KeyExpansionOutput[35]), .Z0_t (KeyExpansionOutput[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U117 ( .A0_t (RoundKey[39]), .B0_t (KeyExpansionOutput[71]), .Z0_t (KeyExpansionOutput[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U116 ( .A0_t (RoundKey[71]), .B0_t (KeyExpansionOutput[103]), .Z0_t (KeyExpansionOutput[71]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U115 ( .A0_t (RoundKey[38]), .B0_t (KeyExpansionOutput[70]), .Z0_t (KeyExpansionOutput[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U114 ( .A0_t (RoundKey[70]), .B0_t (KeyExpansionOutput[102]), .Z0_t (KeyExpansionOutput[70]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U113 ( .A0_t (RoundKey[37]), .B0_t (KeyExpansionOutput[69]), .Z0_t (KeyExpansionOutput[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U112 ( .A0_t (RoundKey[69]), .B0_t (KeyExpansionOutput[101]), .Z0_t (KeyExpansionOutput[69]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U111 ( .A0_t (RoundKey[36]), .B0_t (KeyExpansionOutput[68]), .Z0_t (KeyExpansionOutput[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U110 ( .A0_t (RoundKey[68]), .B0_t (KeyExpansionOutput[100]), .Z0_t (KeyExpansionOutput[68]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U109 ( .A0_t (RoundKey[35]), .B0_t (KeyExpansionOutput[67]), .Z0_t (KeyExpansionOutput[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U108 ( .A0_t (RoundKey[67]), .B0_t (KeyExpansionOutput[99]), .Z0_t (KeyExpansionOutput[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U107 ( .A0_t (RoundKey[99]), .B0_t (KeyExpansionIns_tmp[3]), .Z0_t (KeyExpansionOutput[99]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U106 ( .A0_t (RoundKey[31]), .B0_t (KeyExpansionOutput[63]), .Z0_t (KeyExpansionOutput[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U105 ( .A0_t (RoundKey[63]), .B0_t (KeyExpansionOutput[95]), .Z0_t (KeyExpansionOutput[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U104 ( .A0_t (RoundKey[95]), .B0_t (KeyExpansionOutput[127]), .Z0_t (KeyExpansionOutput[95]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U103 ( .A0_t (RoundKey[30]), .B0_t (KeyExpansionOutput[62]), .Z0_t (KeyExpansionOutput[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U102 ( .A0_t (RoundKey[62]), .B0_t (KeyExpansionOutput[94]), .Z0_t (KeyExpansionOutput[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U101 ( .A0_t (RoundKey[94]), .B0_t (KeyExpansionOutput[126]), .Z0_t (KeyExpansionOutput[94]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U100 ( .A0_t (RoundKey[2]), .B0_t (KeyExpansionOutput[34]), .Z0_t (KeyExpansionOutput[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U99 ( .A0_t (RoundKey[34]), .B0_t (KeyExpansionOutput[66]), .Z0_t (KeyExpansionOutput[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U98 ( .A0_t (RoundKey[66]), .B0_t (KeyExpansionOutput[98]), .Z0_t (KeyExpansionOutput[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U97 ( .A0_t (RoundKey[98]), .B0_t (KeyExpansionIns_tmp[2]), .Z0_t (KeyExpansionOutput[98]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U96 ( .A0_t (RoundKey[29]), .B0_t (KeyExpansionOutput[61]), .Z0_t (KeyExpansionOutput[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U95 ( .A0_t (RoundKey[61]), .B0_t (KeyExpansionOutput[93]), .Z0_t (KeyExpansionOutput[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U94 ( .A0_t (RoundKey[93]), .B0_t (KeyExpansionOutput[125]), .Z0_t (KeyExpansionOutput[93]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U93 ( .A0_t (RoundKey[28]), .B0_t (KeyExpansionOutput[60]), .Z0_t (KeyExpansionOutput[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U92 ( .A0_t (RoundKey[60]), .B0_t (KeyExpansionOutput[92]), .Z0_t (KeyExpansionOutput[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U91 ( .A0_t (RoundKey[92]), .B0_t (KeyExpansionOutput[124]), .Z0_t (KeyExpansionOutput[92]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U90 ( .A0_t (RoundKey[27]), .B0_t (KeyExpansionOutput[59]), .Z0_t (KeyExpansionOutput[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U89 ( .A0_t (RoundKey[59]), .B0_t (KeyExpansionOutput[91]), .Z0_t (KeyExpansionOutput[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U88 ( .A0_t (RoundKey[91]), .B0_t (KeyExpansionOutput[123]), .Z0_t (KeyExpansionOutput[91]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U87 ( .A0_t (RoundKey[26]), .B0_t (KeyExpansionOutput[58]), .Z0_t (KeyExpansionOutput[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U86 ( .A0_t (RoundKey[58]), .B0_t (KeyExpansionOutput[90]), .Z0_t (KeyExpansionOutput[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U85 ( .A0_t (RoundKey[90]), .B0_t (KeyExpansionOutput[122]), .Z0_t (KeyExpansionOutput[90]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U84 ( .A0_t (RoundKey[25]), .B0_t (KeyExpansionOutput[57]), .Z0_t (KeyExpansionOutput[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U83 ( .A0_t (RoundKey[57]), .B0_t (KeyExpansionOutput[89]), .Z0_t (KeyExpansionOutput[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U82 ( .A0_t (RoundKey[89]), .B0_t (KeyExpansionOutput[121]), .Z0_t (KeyExpansionOutput[89]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U81 ( .A0_t (RoundKey[24]), .B0_t (KeyExpansionOutput[56]), .Z0_t (KeyExpansionOutput[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U80 ( .A0_t (RoundKey[56]), .B0_t (KeyExpansionOutput[88]), .Z0_t (KeyExpansionOutput[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U79 ( .A0_t (RoundKey[88]), .B0_t (KeyExpansionOutput[120]), .Z0_t (KeyExpansionOutput[88]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U78 ( .A0_t (RoundKey[23]), .B0_t (KeyExpansionOutput[55]), .Z0_t (KeyExpansionOutput[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U77 ( .A0_t (RoundKey[55]), .B0_t (KeyExpansionOutput[87]), .Z0_t (KeyExpansionOutput[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U76 ( .A0_t (RoundKey[87]), .B0_t (KeyExpansionOutput[119]), .Z0_t (KeyExpansionOutput[87]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U75 ( .A0_t (RoundKey[22]), .B0_t (KeyExpansionOutput[54]), .Z0_t (KeyExpansionOutput[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U74 ( .A0_t (RoundKey[54]), .B0_t (KeyExpansionOutput[86]), .Z0_t (KeyExpansionOutput[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U73 ( .A0_t (RoundKey[86]), .B0_t (KeyExpansionOutput[118]), .Z0_t (KeyExpansionOutput[86]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U72 ( .A0_t (RoundKey[21]), .B0_t (KeyExpansionOutput[53]), .Z0_t (KeyExpansionOutput[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U71 ( .A0_t (RoundKey[53]), .B0_t (KeyExpansionOutput[85]), .Z0_t (KeyExpansionOutput[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U70 ( .A0_t (RoundKey[85]), .B0_t (KeyExpansionOutput[117]), .Z0_t (KeyExpansionOutput[85]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U69 ( .A0_t (RoundKey[20]), .B0_t (KeyExpansionOutput[52]), .Z0_t (KeyExpansionOutput[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U68 ( .A0_t (RoundKey[52]), .B0_t (KeyExpansionOutput[84]), .Z0_t (KeyExpansionOutput[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U67 ( .A0_t (RoundKey[84]), .B0_t (KeyExpansionOutput[116]), .Z0_t (KeyExpansionOutput[84]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U66 ( .A0_t (RoundKey[1]), .B0_t (KeyExpansionOutput[33]), .Z0_t (KeyExpansionOutput[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U65 ( .A0_t (RoundKey[33]), .B0_t (KeyExpansionOutput[65]), .Z0_t (KeyExpansionOutput[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U64 ( .A0_t (RoundKey[65]), .B0_t (KeyExpansionOutput[97]), .Z0_t (KeyExpansionOutput[65]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U63 ( .A0_t (RoundKey[97]), .B0_t (KeyExpansionIns_tmp[1]), .Z0_t (KeyExpansionOutput[97]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U62 ( .A0_t (RoundKey[19]), .B0_t (KeyExpansionOutput[51]), .Z0_t (KeyExpansionOutput[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U61 ( .A0_t (RoundKey[51]), .B0_t (KeyExpansionOutput[83]), .Z0_t (KeyExpansionOutput[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U60 ( .A0_t (RoundKey[83]), .B0_t (KeyExpansionOutput[115]), .Z0_t (KeyExpansionOutput[83]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U59 ( .A0_t (RoundKey[18]), .B0_t (KeyExpansionOutput[50]), .Z0_t (KeyExpansionOutput[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U58 ( .A0_t (RoundKey[50]), .B0_t (KeyExpansionOutput[82]), .Z0_t (KeyExpansionOutput[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U57 ( .A0_t (RoundKey[82]), .B0_t (KeyExpansionOutput[114]), .Z0_t (KeyExpansionOutput[82]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U56 ( .A0_t (RoundKey[17]), .B0_t (KeyExpansionOutput[49]), .Z0_t (KeyExpansionOutput[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U55 ( .A0_t (RoundKey[49]), .B0_t (KeyExpansionOutput[81]), .Z0_t (KeyExpansionOutput[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U54 ( .A0_t (RoundKey[81]), .B0_t (KeyExpansionOutput[113]), .Z0_t (KeyExpansionOutput[81]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U53 ( .A0_t (RoundKey[16]), .B0_t (KeyExpansionOutput[48]), .Z0_t (KeyExpansionOutput[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U52 ( .A0_t (RoundKey[48]), .B0_t (KeyExpansionOutput[80]), .Z0_t (KeyExpansionOutput[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U51 ( .A0_t (RoundKey[80]), .B0_t (KeyExpansionOutput[112]), .Z0_t (KeyExpansionOutput[80]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U50 ( .A0_t (RoundKey[15]), .B0_t (KeyExpansionOutput[47]), .Z0_t (KeyExpansionOutput[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U49 ( .A0_t (RoundKey[47]), .B0_t (KeyExpansionOutput[79]), .Z0_t (KeyExpansionOutput[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U48 ( .A0_t (RoundKey[79]), .B0_t (KeyExpansionOutput[111]), .Z0_t (KeyExpansionOutput[79]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U47 ( .A0_t (RoundKey[14]), .B0_t (KeyExpansionOutput[46]), .Z0_t (KeyExpansionOutput[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U46 ( .A0_t (RoundKey[46]), .B0_t (KeyExpansionOutput[78]), .Z0_t (KeyExpansionOutput[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U45 ( .A0_t (RoundKey[78]), .B0_t (KeyExpansionOutput[110]), .Z0_t (KeyExpansionOutput[78]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U44 ( .A0_t (RoundKey[13]), .B0_t (KeyExpansionOutput[45]), .Z0_t (KeyExpansionOutput[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U43 ( .A0_t (RoundKey[45]), .B0_t (KeyExpansionOutput[77]), .Z0_t (KeyExpansionOutput[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U42 ( .A0_t (RoundKey[77]), .B0_t (KeyExpansionOutput[109]), .Z0_t (KeyExpansionOutput[77]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U41 ( .A0_t (RoundKey[12]), .B0_t (KeyExpansionOutput[44]), .Z0_t (KeyExpansionOutput[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U40 ( .A0_t (RoundKey[44]), .B0_t (KeyExpansionOutput[76]), .Z0_t (KeyExpansionOutput[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U39 ( .A0_t (RoundKey[76]), .B0_t (KeyExpansionOutput[108]), .Z0_t (KeyExpansionOutput[76]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U38 ( .A0_t (RoundKey[127]), .B0_t (KeyExpansionIns_tmp[31]), .Z0_t (KeyExpansionOutput[127]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U37 ( .A0_t (RoundKey[126]), .B0_t (KeyExpansionIns_tmp[30]), .Z0_t (KeyExpansionOutput[126]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U36 ( .A0_t (RoundKey[125]), .B0_t (KeyExpansionIns_tmp[29]), .Z0_t (KeyExpansionOutput[125]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U35 ( .A0_t (RoundKey[124]), .B0_t (KeyExpansionIns_tmp[28]), .Z0_t (KeyExpansionOutput[124]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U34 ( .A0_t (RoundKey[123]), .B0_t (KeyExpansionIns_tmp[27]), .Z0_t (KeyExpansionOutput[123]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U33 ( .A0_t (RoundKey[122]), .B0_t (KeyExpansionIns_tmp[26]), .Z0_t (KeyExpansionOutput[122]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U32 ( .A0_t (RoundKey[121]), .B0_t (KeyExpansionIns_tmp[25]), .Z0_t (KeyExpansionOutput[121]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U31 ( .A0_t (RoundKey[120]), .B0_t (KeyExpansionIns_tmp[24]), .Z0_t (KeyExpansionOutput[120]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U30 ( .A0_t (RoundKey[11]), .B0_t (KeyExpansionOutput[43]), .Z0_t (KeyExpansionOutput[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U29 ( .A0_t (RoundKey[43]), .B0_t (KeyExpansionOutput[75]), .Z0_t (KeyExpansionOutput[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U28 ( .A0_t (RoundKey[75]), .B0_t (KeyExpansionOutput[107]), .Z0_t (KeyExpansionOutput[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U27 ( .A0_t (RoundKey[119]), .B0_t (KeyExpansionIns_tmp[23]), .Z0_t (KeyExpansionOutput[119]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U26 ( .A0_t (RoundKey[118]), .B0_t (KeyExpansionIns_tmp[22]), .Z0_t (KeyExpansionOutput[118]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U25 ( .A0_t (RoundKey[117]), .B0_t (KeyExpansionIns_tmp[21]), .Z0_t (KeyExpansionOutput[117]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U24 ( .A0_t (RoundKey[116]), .B0_t (KeyExpansionIns_tmp[20]), .Z0_t (KeyExpansionOutput[116]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U23 ( .A0_t (RoundKey[115]), .B0_t (KeyExpansionIns_tmp[19]), .Z0_t (KeyExpansionOutput[115]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U22 ( .A0_t (RoundKey[114]), .B0_t (KeyExpansionIns_tmp[18]), .Z0_t (KeyExpansionOutput[114]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U21 ( .A0_t (RoundKey[113]), .B0_t (KeyExpansionIns_tmp[17]), .Z0_t (KeyExpansionOutput[113]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U20 ( .A0_t (RoundKey[112]), .B0_t (KeyExpansionIns_tmp[16]), .Z0_t (KeyExpansionOutput[112]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U19 ( .A0_t (RoundKey[111]), .B0_t (KeyExpansionIns_tmp[15]), .Z0_t (KeyExpansionOutput[111]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U18 ( .A0_t (RoundKey[110]), .B0_t (KeyExpansionIns_tmp[14]), .Z0_t (KeyExpansionOutput[110]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U17 ( .A0_t (RoundKey[10]), .B0_t (KeyExpansionOutput[42]), .Z0_t (KeyExpansionOutput[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U16 ( .A0_t (RoundKey[42]), .B0_t (KeyExpansionOutput[74]), .Z0_t (KeyExpansionOutput[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U15 ( .A0_t (RoundKey[74]), .B0_t (KeyExpansionOutput[106]), .Z0_t (KeyExpansionOutput[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U14 ( .A0_t (RoundKey[109]), .B0_t (KeyExpansionIns_tmp[13]), .Z0_t (KeyExpansionOutput[109]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U13 ( .A0_t (RoundKey[108]), .B0_t (KeyExpansionIns_tmp[12]), .Z0_t (KeyExpansionOutput[108]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U12 ( .A0_t (RoundKey[107]), .B0_t (KeyExpansionIns_tmp[11]), .Z0_t (KeyExpansionOutput[107]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U11 ( .A0_t (RoundKey[106]), .B0_t (KeyExpansionIns_tmp[10]), .Z0_t (KeyExpansionOutput[106]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U10 ( .A0_t (RoundKey[105]), .B0_t (KeyExpansionIns_tmp[9]), .Z0_t (KeyExpansionOutput[105]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U9 ( .A0_t (RoundKey[104]), .B0_t (KeyExpansionIns_tmp[8]), .Z0_t (KeyExpansionOutput[104]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U8 ( .A0_t (RoundKey[103]), .B0_t (KeyExpansionIns_tmp[7]), .Z0_t (KeyExpansionOutput[103]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U7 ( .A0_t (RoundKey[102]), .B0_t (KeyExpansionIns_tmp[6]), .Z0_t (KeyExpansionOutput[102]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U6 ( .A0_t (RoundKey[101]), .B0_t (KeyExpansionIns_tmp[5]), .Z0_t (KeyExpansionOutput[101]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U5 ( .A0_t (RoundKey[100]), .B0_t (KeyExpansionIns_tmp[4]), .Z0_t (KeyExpansionOutput[100]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U4 ( .A0_t (RoundKey[0]), .B0_t (KeyExpansionOutput[32]), .Z0_t (KeyExpansionOutput[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U3 ( .A0_t (RoundKey[32]), .B0_t (KeyExpansionOutput[64]), .Z0_t (KeyExpansionOutput[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U2 ( .A0_t (RoundKey[64]), .B0_t (KeyExpansionOutput[96]), .Z0_t (KeyExpansionOutput[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_U1 ( .A0_t (RoundKey[96]), .B0_t (KeyExpansionIns_tmp[0]), .Z0_t (KeyExpansionOutput[96]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U8 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_), .B0_t (n283), .Z0_t (KeyExpansionIns_tmp[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U7 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_), .B0_t (n285), .Z0_t (KeyExpansionIns_tmp[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U6 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_), .B0_t (Rcon[5]), .Z0_t (KeyExpansionIns_tmp[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U5 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_), .B0_t (Rcon[4]), .Z0_t (KeyExpansionIns_tmp[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U4 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_), .B0_t (Rcon[3]), .Z0_t (KeyExpansionIns_tmp[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U3 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_), .B0_t (Rcon[2]), .Z0_t (KeyExpansionIns_tmp[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U2 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_), .B0_t (Rcon[1]), .Z0_t (KeyExpansionIns_tmp[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_), .B0_t (Rcon[0]), .Z0_t (KeyExpansionIns_tmp[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T1_U1 ( .A0_t (RoundKey[23]), .B0_t (RoundKey[20]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T2_U1 ( .A0_t (RoundKey[23]), .B0_t (RoundKey[18]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T3_U1 ( .A0_t (RoundKey[23]), .B0_t (RoundKey[17]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T4_U1 ( .A0_t (RoundKey[20]), .B0_t (RoundKey[18]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T5_U1 ( .A0_t (RoundKey[19]), .B0_t (RoundKey[17]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T7_U1 ( .A0_t (RoundKey[22]), .B0_t (RoundKey[21]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T8_U1 ( .A0_t (RoundKey[16]), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T9_U1 ( .A0_t (RoundKey[16]), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T11_U1 ( .A0_t (RoundKey[22]), .B0_t (RoundKey[18]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T12_U1 ( .A0_t (RoundKey[21]), .B0_t (RoundKey[18]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T18_U1 ( .A0_t (RoundKey[20]), .B0_t (RoundKey[16]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T21_U1 ( .A0_t (RoundKey[17]), .B0_t (RoundKey[16]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .B0_t (RoundKey[16]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M30_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M31_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M32_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M33_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M34_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M35_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M36_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M37_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M38_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M39_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M40_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M41_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M42_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M43_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M44_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M45_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M46_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M47_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M48_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .B0_t (RoundKey[16]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M49_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M50_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M51_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M52_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M53_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M54_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M55_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M56_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M57_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M58_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M59_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M60_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M61_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M62_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M63_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T1_U1 ( .A0_t (RoundKey[15]), .B0_t (RoundKey[12]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T2_U1 ( .A0_t (RoundKey[15]), .B0_t (RoundKey[10]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T3_U1 ( .A0_t (RoundKey[15]), .B0_t (RoundKey[9]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T4_U1 ( .A0_t (RoundKey[12]), .B0_t (RoundKey[10]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T5_U1 ( .A0_t (RoundKey[11]), .B0_t (RoundKey[9]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T7_U1 ( .A0_t (RoundKey[14]), .B0_t (RoundKey[13]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T8_U1 ( .A0_t (RoundKey[8]), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T9_U1 ( .A0_t (RoundKey[8]), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T11_U1 ( .A0_t (RoundKey[14]), .B0_t (RoundKey[10]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T12_U1 ( .A0_t (RoundKey[13]), .B0_t (RoundKey[10]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T18_U1 ( .A0_t (RoundKey[12]), .B0_t (RoundKey[8]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T21_U1 ( .A0_t (RoundKey[9]), .B0_t (RoundKey[8]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .B0_t (RoundKey[8]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M30_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M31_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M32_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M33_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M34_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M35_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M36_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M37_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M38_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M39_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M40_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M41_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M42_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M43_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M44_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M45_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M46_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M47_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M48_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .B0_t (RoundKey[8]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M49_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M50_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M51_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M52_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M53_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M54_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M55_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M56_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M57_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M58_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M59_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M60_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M61_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M62_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M63_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24), .Z0_t (KeyExpansionIns_tmp[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26), .Z0_t (KeyExpansionIns_tmp[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28), .Z0_t (KeyExpansionIns_tmp[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21), .Z0_t (KeyExpansionIns_tmp[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22), .Z0_t (KeyExpansionIns_tmp[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29), .Z0_t (KeyExpansionIns_tmp[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27), .Z0_t (KeyExpansionIns_tmp[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23), .Z0_t (KeyExpansionIns_tmp[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T1_U1 ( .A0_t (RoundKey[7]), .B0_t (RoundKey[4]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T2_U1 ( .A0_t (RoundKey[7]), .B0_t (RoundKey[2]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T3_U1 ( .A0_t (RoundKey[7]), .B0_t (RoundKey[1]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T4_U1 ( .A0_t (RoundKey[4]), .B0_t (RoundKey[2]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T5_U1 ( .A0_t (RoundKey[3]), .B0_t (RoundKey[1]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T7_U1 ( .A0_t (RoundKey[6]), .B0_t (RoundKey[5]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T8_U1 ( .A0_t (RoundKey[0]), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T9_U1 ( .A0_t (RoundKey[0]), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T11_U1 ( .A0_t (RoundKey[6]), .B0_t (RoundKey[2]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T12_U1 ( .A0_t (RoundKey[5]), .B0_t (RoundKey[2]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T18_U1 ( .A0_t (RoundKey[4]), .B0_t (RoundKey[0]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T21_U1 ( .A0_t (RoundKey[1]), .B0_t (RoundKey[0]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .B0_t (RoundKey[0]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M30_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M31_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M32_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M33_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M34_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M35_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M36_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M37_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M38_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M39_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M40_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M41_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M42_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M43_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M44_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M45_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M46_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M47_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M48_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .B0_t (RoundKey[0]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M49_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M50_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M51_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M52_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M53_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M54_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M55_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M56_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M57_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M58_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M59_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M60_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M61_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M62_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M63_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24), .Z0_t (KeyExpansionIns_tmp[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26), .Z0_t (KeyExpansionIns_tmp[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28), .Z0_t (KeyExpansionIns_tmp[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21), .Z0_t (KeyExpansionIns_tmp[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22), .Z0_t (KeyExpansionIns_tmp[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29), .Z0_t (KeyExpansionIns_tmp[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27), .Z0_t (KeyExpansionIns_tmp[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23), .Z0_t (KeyExpansionIns_tmp[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T1_U1 ( .A0_t (RoundKey[31]), .B0_t (RoundKey[28]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T2_U1 ( .A0_t (RoundKey[31]), .B0_t (RoundKey[26]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T3_U1 ( .A0_t (RoundKey[31]), .B0_t (RoundKey[25]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T4_U1 ( .A0_t (RoundKey[28]), .B0_t (RoundKey[26]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T5_U1 ( .A0_t (RoundKey[27]), .B0_t (RoundKey[25]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T7_U1 ( .A0_t (RoundKey[30]), .B0_t (RoundKey[29]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T8_U1 ( .A0_t (RoundKey[24]), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T9_U1 ( .A0_t (RoundKey[24]), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T11_U1 ( .A0_t (RoundKey[30]), .B0_t (RoundKey[26]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T12_U1 ( .A0_t (RoundKey[29]), .B0_t (RoundKey[26]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T18_U1 ( .A0_t (RoundKey[28]), .B0_t (RoundKey[24]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T21_U1 ( .A0_t (RoundKey[25]), .B0_t (RoundKey[24]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .B0_t (RoundKey[24]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M30_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M31_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M32_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M33_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M34_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M35_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M36_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M37_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M38_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M39_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M40_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M41_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M42_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M43_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M44_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M45_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M46_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M47_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M48_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .B0_t (RoundKey[24]), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M49_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M50_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M51_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M52_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M53_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M54_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M55_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M56_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M57_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M58_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M59_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M60_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M61_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M62_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M63_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L8_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L9_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L10_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L11_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L12_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L13_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L14_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L15_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L16_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L17_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L18_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L19_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L20_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L21_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L22_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L23_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L24_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L25_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L26_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L27_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L28_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L29_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17), .Z0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S0_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24), .Z0_t (KeyExpansionIns_tmp[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S1_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26), .Z0_t (KeyExpansionIns_tmp[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S2_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28), .Z0_t (KeyExpansionIns_tmp[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S3_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21), .Z0_t (KeyExpansionIns_tmp[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S4_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22), .Z0_t (KeyExpansionIns_tmp[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S5_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29), .Z0_t (KeyExpansionIns_tmp[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S6_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27), .Z0_t (KeyExpansionIns_tmp[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S7_U1 ( .A0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B0_t (KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23), .Z0_t (KeyExpansionIns_tmp[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) RoundCounterIns_U11 ( .A0_t (start), .B0_t (RoundCounterIns_n5), .Z0_t (RoundCounter[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) RoundCounterIns_U10 ( .A0_t (RoundCounter[2]), .B0_t (RoundCounterIns_n4), .Z0_t (RoundCounterIns_n5) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) RoundCounterIns_U9 ( .A0_t (start), .B0_t (RoundCounterIns_n3), .Z0_t (RoundCounter[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) RoundCounterIns_U8 ( .A0_t (RoundCounter[1]), .B0_t (RoundCounter[0]), .Z0_t (RoundCounterIns_n3) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) RoundCounterIns_U7 ( .A0_t (start), .B0_t (RoundCounterIns_n2), .Z0_t (RoundCounter[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) RoundCounterIns_U6 ( .A0_t (RoundCounter[3]), .B0_t (RoundCounterIns_n1), .Z0_t (RoundCounterIns_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) RoundCounterIns_U5 ( .A0_t (RoundCounterIns_n4), .B0_t (RoundCounter[2]), .Z0_t (RoundCounterIns_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) RoundCounterIns_U4 ( .A0_t (RoundCounter[0]), .B0_t (RoundCounter[1]), .Z0_t (RoundCounterIns_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) RoundCounterIns_U3 ( .A0_t (start), .B0_t (RoundCounter[0]), .Z0_t (RoundCounter[0]) ) ;

    /* register cells */
endmodule
