/* modified netlist. Source: module Cipher in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/10_CRAFT_round_based_encryption_PortParallel/4-AGEMA/Cipher.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module Cipher_SAUBER_Pipeline_d1 (Input_s0_t, Key_s0_t, rst_t, Key_s0_f, Key_s1_t, Key_s1_f, rst_f, Input_s0_f, Input_s1_t, Input_s1_f, Output_s0_t, done_t, Output_s0_f, Output_s1_t, Output_s1_f, done_f);
    input [63:0] Input_s0_t ;
    input [127:0] Key_s0_t ;
    input rst_t ;
    input [127:0] Key_s0_f ;
    input [127:0] Key_s1_t ;
    input [127:0] Key_s1_f ;
    input rst_f ;
    input [63:0] Input_s0_f ;
    input [63:0] Input_s1_t ;
    input [63:0] Input_s1_f ;
    output [63:0] Output_s0_t ;
    output done_t ;
    output [63:0] Output_s0_f ;
    output [63:0] Output_s1_t ;
    output [63:0] Output_s1_f ;
    output done_f ;
    wire RoundConstant_4_ ;
    wire RoundConstant_0 ;
    wire InputMUX_MUXInst_0_U1_Y ;
    wire InputMUX_MUXInst_0_U1_X ;
    wire InputMUX_MUXInst_1_U1_Y ;
    wire InputMUX_MUXInst_1_U1_X ;
    wire InputMUX_MUXInst_2_U1_Y ;
    wire InputMUX_MUXInst_2_U1_X ;
    wire InputMUX_MUXInst_3_U1_Y ;
    wire InputMUX_MUXInst_3_U1_X ;
    wire InputMUX_MUXInst_4_U1_Y ;
    wire InputMUX_MUXInst_4_U1_X ;
    wire InputMUX_MUXInst_5_U1_Y ;
    wire InputMUX_MUXInst_5_U1_X ;
    wire InputMUX_MUXInst_6_U1_Y ;
    wire InputMUX_MUXInst_6_U1_X ;
    wire InputMUX_MUXInst_7_U1_Y ;
    wire InputMUX_MUXInst_7_U1_X ;
    wire InputMUX_MUXInst_8_U1_Y ;
    wire InputMUX_MUXInst_8_U1_X ;
    wire InputMUX_MUXInst_9_U1_Y ;
    wire InputMUX_MUXInst_9_U1_X ;
    wire InputMUX_MUXInst_10_U1_Y ;
    wire InputMUX_MUXInst_10_U1_X ;
    wire InputMUX_MUXInst_11_U1_Y ;
    wire InputMUX_MUXInst_11_U1_X ;
    wire InputMUX_MUXInst_12_U1_Y ;
    wire InputMUX_MUXInst_12_U1_X ;
    wire InputMUX_MUXInst_13_U1_Y ;
    wire InputMUX_MUXInst_13_U1_X ;
    wire InputMUX_MUXInst_14_U1_Y ;
    wire InputMUX_MUXInst_14_U1_X ;
    wire InputMUX_MUXInst_15_U1_Y ;
    wire InputMUX_MUXInst_15_U1_X ;
    wire InputMUX_MUXInst_16_U1_Y ;
    wire InputMUX_MUXInst_16_U1_X ;
    wire InputMUX_MUXInst_17_U1_Y ;
    wire InputMUX_MUXInst_17_U1_X ;
    wire InputMUX_MUXInst_18_U1_Y ;
    wire InputMUX_MUXInst_18_U1_X ;
    wire InputMUX_MUXInst_19_U1_Y ;
    wire InputMUX_MUXInst_19_U1_X ;
    wire InputMUX_MUXInst_20_U1_Y ;
    wire InputMUX_MUXInst_20_U1_X ;
    wire InputMUX_MUXInst_21_U1_Y ;
    wire InputMUX_MUXInst_21_U1_X ;
    wire InputMUX_MUXInst_22_U1_Y ;
    wire InputMUX_MUXInst_22_U1_X ;
    wire InputMUX_MUXInst_23_U1_Y ;
    wire InputMUX_MUXInst_23_U1_X ;
    wire InputMUX_MUXInst_24_U1_Y ;
    wire InputMUX_MUXInst_24_U1_X ;
    wire InputMUX_MUXInst_25_U1_Y ;
    wire InputMUX_MUXInst_25_U1_X ;
    wire InputMUX_MUXInst_26_U1_Y ;
    wire InputMUX_MUXInst_26_U1_X ;
    wire InputMUX_MUXInst_27_U1_Y ;
    wire InputMUX_MUXInst_27_U1_X ;
    wire InputMUX_MUXInst_28_U1_Y ;
    wire InputMUX_MUXInst_28_U1_X ;
    wire InputMUX_MUXInst_29_U1_Y ;
    wire InputMUX_MUXInst_29_U1_X ;
    wire InputMUX_MUXInst_30_U1_Y ;
    wire InputMUX_MUXInst_30_U1_X ;
    wire InputMUX_MUXInst_31_U1_Y ;
    wire InputMUX_MUXInst_31_U1_X ;
    wire InputMUX_MUXInst_32_U1_Y ;
    wire InputMUX_MUXInst_32_U1_X ;
    wire InputMUX_MUXInst_33_U1_Y ;
    wire InputMUX_MUXInst_33_U1_X ;
    wire InputMUX_MUXInst_34_U1_Y ;
    wire InputMUX_MUXInst_34_U1_X ;
    wire InputMUX_MUXInst_35_U1_Y ;
    wire InputMUX_MUXInst_35_U1_X ;
    wire InputMUX_MUXInst_36_U1_Y ;
    wire InputMUX_MUXInst_36_U1_X ;
    wire InputMUX_MUXInst_37_U1_Y ;
    wire InputMUX_MUXInst_37_U1_X ;
    wire InputMUX_MUXInst_38_U1_Y ;
    wire InputMUX_MUXInst_38_U1_X ;
    wire InputMUX_MUXInst_39_U1_Y ;
    wire InputMUX_MUXInst_39_U1_X ;
    wire InputMUX_MUXInst_40_U1_Y ;
    wire InputMUX_MUXInst_40_U1_X ;
    wire InputMUX_MUXInst_41_U1_Y ;
    wire InputMUX_MUXInst_41_U1_X ;
    wire InputMUX_MUXInst_42_U1_Y ;
    wire InputMUX_MUXInst_42_U1_X ;
    wire InputMUX_MUXInst_43_U1_Y ;
    wire InputMUX_MUXInst_43_U1_X ;
    wire InputMUX_MUXInst_44_U1_Y ;
    wire InputMUX_MUXInst_44_U1_X ;
    wire InputMUX_MUXInst_45_U1_Y ;
    wire InputMUX_MUXInst_45_U1_X ;
    wire InputMUX_MUXInst_46_U1_Y ;
    wire InputMUX_MUXInst_46_U1_X ;
    wire InputMUX_MUXInst_47_U1_Y ;
    wire InputMUX_MUXInst_47_U1_X ;
    wire InputMUX_MUXInst_48_U1_Y ;
    wire InputMUX_MUXInst_48_U1_X ;
    wire InputMUX_MUXInst_49_U1_Y ;
    wire InputMUX_MUXInst_49_U1_X ;
    wire InputMUX_MUXInst_50_U1_Y ;
    wire InputMUX_MUXInst_50_U1_X ;
    wire InputMUX_MUXInst_51_U1_Y ;
    wire InputMUX_MUXInst_51_U1_X ;
    wire InputMUX_MUXInst_52_U1_Y ;
    wire InputMUX_MUXInst_52_U1_X ;
    wire InputMUX_MUXInst_53_U1_Y ;
    wire InputMUX_MUXInst_53_U1_X ;
    wire InputMUX_MUXInst_54_U1_Y ;
    wire InputMUX_MUXInst_54_U1_X ;
    wire InputMUX_MUXInst_55_U1_Y ;
    wire InputMUX_MUXInst_55_U1_X ;
    wire InputMUX_MUXInst_56_U1_Y ;
    wire InputMUX_MUXInst_56_U1_X ;
    wire InputMUX_MUXInst_57_U1_Y ;
    wire InputMUX_MUXInst_57_U1_X ;
    wire InputMUX_MUXInst_58_U1_Y ;
    wire InputMUX_MUXInst_58_U1_X ;
    wire InputMUX_MUXInst_59_U1_Y ;
    wire InputMUX_MUXInst_59_U1_X ;
    wire InputMUX_MUXInst_60_U1_Y ;
    wire InputMUX_MUXInst_60_U1_X ;
    wire InputMUX_MUXInst_61_U1_Y ;
    wire InputMUX_MUXInst_61_U1_X ;
    wire InputMUX_MUXInst_62_U1_Y ;
    wire InputMUX_MUXInst_62_U1_X ;
    wire InputMUX_MUXInst_63_U1_Y ;
    wire InputMUX_MUXInst_63_U1_X ;
    wire MCInst_XOR_r0_Inst_0_n1 ;
    wire MCInst_XOR_r0_Inst_1_n1 ;
    wire MCInst_XOR_r0_Inst_2_n1 ;
    wire MCInst_XOR_r0_Inst_3_n1 ;
    wire MCInst_XOR_r0_Inst_4_n1 ;
    wire MCInst_XOR_r0_Inst_5_n1 ;
    wire MCInst_XOR_r0_Inst_6_n1 ;
    wire MCInst_XOR_r0_Inst_7_n1 ;
    wire MCInst_XOR_r0_Inst_8_n1 ;
    wire MCInst_XOR_r0_Inst_9_n1 ;
    wire MCInst_XOR_r0_Inst_10_n1 ;
    wire MCInst_XOR_r0_Inst_11_n1 ;
    wire MCInst_XOR_r0_Inst_12_n1 ;
    wire MCInst_XOR_r0_Inst_13_n1 ;
    wire MCInst_XOR_r0_Inst_14_n1 ;
    wire MCInst_XOR_r0_Inst_15_n1 ;
    wire AddKeyConstXOR_XORInst_0_0_n1 ;
    wire AddKeyConstXOR_XORInst_0_1_n1 ;
    wire AddKeyConstXOR_XORInst_0_2_n1 ;
    wire AddKeyConstXOR_XORInst_1_0_n1 ;
    wire AddKeyConstXOR_XORInst_1_1_n1 ;
    wire AddKeyConstXOR_XORInst_1_2_n1 ;
    wire AddKeyConstXOR_XORInst_1_3_n1 ;
    wire SubCellInst_SboxInst_0_n15 ;
    wire SubCellInst_SboxInst_0_n14 ;
    wire SubCellInst_SboxInst_0_n13 ;
    wire SubCellInst_SboxInst_0_n11 ;
    wire SubCellInst_SboxInst_0_n10 ;
    wire SubCellInst_SboxInst_0_n9 ;
    wire SubCellInst_SboxInst_0_n7 ;
    wire SubCellInst_SboxInst_0_n6 ;
    wire SubCellInst_SboxInst_0_n5 ;
    wire SubCellInst_SboxInst_0_n4 ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_n1 ;
    wire SubCellInst_SboxInst_1_n15 ;
    wire SubCellInst_SboxInst_1_n14 ;
    wire SubCellInst_SboxInst_1_n13 ;
    wire SubCellInst_SboxInst_1_n11 ;
    wire SubCellInst_SboxInst_1_n10 ;
    wire SubCellInst_SboxInst_1_n9 ;
    wire SubCellInst_SboxInst_1_n7 ;
    wire SubCellInst_SboxInst_1_n6 ;
    wire SubCellInst_SboxInst_1_n5 ;
    wire SubCellInst_SboxInst_1_n4 ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_n1 ;
    wire SubCellInst_SboxInst_2_n15 ;
    wire SubCellInst_SboxInst_2_n14 ;
    wire SubCellInst_SboxInst_2_n13 ;
    wire SubCellInst_SboxInst_2_n11 ;
    wire SubCellInst_SboxInst_2_n10 ;
    wire SubCellInst_SboxInst_2_n9 ;
    wire SubCellInst_SboxInst_2_n7 ;
    wire SubCellInst_SboxInst_2_n6 ;
    wire SubCellInst_SboxInst_2_n5 ;
    wire SubCellInst_SboxInst_2_n4 ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_n1 ;
    wire SubCellInst_SboxInst_3_n15 ;
    wire SubCellInst_SboxInst_3_n14 ;
    wire SubCellInst_SboxInst_3_n13 ;
    wire SubCellInst_SboxInst_3_n11 ;
    wire SubCellInst_SboxInst_3_n10 ;
    wire SubCellInst_SboxInst_3_n9 ;
    wire SubCellInst_SboxInst_3_n7 ;
    wire SubCellInst_SboxInst_3_n6 ;
    wire SubCellInst_SboxInst_3_n5 ;
    wire SubCellInst_SboxInst_3_n4 ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_n1 ;
    wire SubCellInst_SboxInst_4_n15 ;
    wire SubCellInst_SboxInst_4_n14 ;
    wire SubCellInst_SboxInst_4_n13 ;
    wire SubCellInst_SboxInst_4_n10 ;
    wire SubCellInst_SboxInst_4_n9 ;
    wire SubCellInst_SboxInst_4_n8 ;
    wire SubCellInst_SboxInst_4_n7 ;
    wire SubCellInst_SboxInst_4_n6 ;
    wire SubCellInst_SboxInst_4_n5 ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_n2 ;
    wire SubCellInst_SboxInst_4_n1 ;
    wire SubCellInst_SboxInst_5_n15 ;
    wire SubCellInst_SboxInst_5_n14 ;
    wire SubCellInst_SboxInst_5_n13 ;
    wire SubCellInst_SboxInst_5_n10 ;
    wire SubCellInst_SboxInst_5_n9 ;
    wire SubCellInst_SboxInst_5_n8 ;
    wire SubCellInst_SboxInst_5_n7 ;
    wire SubCellInst_SboxInst_5_n6 ;
    wire SubCellInst_SboxInst_5_n5 ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_n2 ;
    wire SubCellInst_SboxInst_5_n1 ;
    wire SubCellInst_SboxInst_6_n15 ;
    wire SubCellInst_SboxInst_6_n14 ;
    wire SubCellInst_SboxInst_6_n13 ;
    wire SubCellInst_SboxInst_6_n10 ;
    wire SubCellInst_SboxInst_6_n9 ;
    wire SubCellInst_SboxInst_6_n8 ;
    wire SubCellInst_SboxInst_6_n7 ;
    wire SubCellInst_SboxInst_6_n6 ;
    wire SubCellInst_SboxInst_6_n5 ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_n2 ;
    wire SubCellInst_SboxInst_6_n1 ;
    wire SubCellInst_SboxInst_7_n15 ;
    wire SubCellInst_SboxInst_7_n14 ;
    wire SubCellInst_SboxInst_7_n13 ;
    wire SubCellInst_SboxInst_7_n10 ;
    wire SubCellInst_SboxInst_7_n9 ;
    wire SubCellInst_SboxInst_7_n8 ;
    wire SubCellInst_SboxInst_7_n7 ;
    wire SubCellInst_SboxInst_7_n6 ;
    wire SubCellInst_SboxInst_7_n5 ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_n2 ;
    wire SubCellInst_SboxInst_7_n1 ;
    wire SubCellInst_SboxInst_8_n15 ;
    wire SubCellInst_SboxInst_8_n14 ;
    wire SubCellInst_SboxInst_8_n13 ;
    wire SubCellInst_SboxInst_8_n10 ;
    wire SubCellInst_SboxInst_8_n9 ;
    wire SubCellInst_SboxInst_8_n8 ;
    wire SubCellInst_SboxInst_8_n7 ;
    wire SubCellInst_SboxInst_8_n6 ;
    wire SubCellInst_SboxInst_8_n5 ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_n2 ;
    wire SubCellInst_SboxInst_8_n1 ;
    wire SubCellInst_SboxInst_9_n15 ;
    wire SubCellInst_SboxInst_9_n14 ;
    wire SubCellInst_SboxInst_9_n13 ;
    wire SubCellInst_SboxInst_9_n10 ;
    wire SubCellInst_SboxInst_9_n9 ;
    wire SubCellInst_SboxInst_9_n8 ;
    wire SubCellInst_SboxInst_9_n7 ;
    wire SubCellInst_SboxInst_9_n6 ;
    wire SubCellInst_SboxInst_9_n5 ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_n2 ;
    wire SubCellInst_SboxInst_9_n1 ;
    wire SubCellInst_SboxInst_10_n15 ;
    wire SubCellInst_SboxInst_10_n14 ;
    wire SubCellInst_SboxInst_10_n13 ;
    wire SubCellInst_SboxInst_10_n10 ;
    wire SubCellInst_SboxInst_10_n9 ;
    wire SubCellInst_SboxInst_10_n8 ;
    wire SubCellInst_SboxInst_10_n7 ;
    wire SubCellInst_SboxInst_10_n6 ;
    wire SubCellInst_SboxInst_10_n5 ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_n2 ;
    wire SubCellInst_SboxInst_10_n1 ;
    wire SubCellInst_SboxInst_11_n15 ;
    wire SubCellInst_SboxInst_11_n14 ;
    wire SubCellInst_SboxInst_11_n13 ;
    wire SubCellInst_SboxInst_11_n10 ;
    wire SubCellInst_SboxInst_11_n9 ;
    wire SubCellInst_SboxInst_11_n8 ;
    wire SubCellInst_SboxInst_11_n7 ;
    wire SubCellInst_SboxInst_11_n6 ;
    wire SubCellInst_SboxInst_11_n5 ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_n2 ;
    wire SubCellInst_SboxInst_11_n1 ;
    wire SubCellInst_SboxInst_12_n15 ;
    wire SubCellInst_SboxInst_12_n14 ;
    wire SubCellInst_SboxInst_12_n13 ;
    wire SubCellInst_SboxInst_12_n10 ;
    wire SubCellInst_SboxInst_12_n9 ;
    wire SubCellInst_SboxInst_12_n8 ;
    wire SubCellInst_SboxInst_12_n7 ;
    wire SubCellInst_SboxInst_12_n6 ;
    wire SubCellInst_SboxInst_12_n5 ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_n2 ;
    wire SubCellInst_SboxInst_12_n1 ;
    wire SubCellInst_SboxInst_13_n15 ;
    wire SubCellInst_SboxInst_13_n14 ;
    wire SubCellInst_SboxInst_13_n13 ;
    wire SubCellInst_SboxInst_13_n10 ;
    wire SubCellInst_SboxInst_13_n9 ;
    wire SubCellInst_SboxInst_13_n8 ;
    wire SubCellInst_SboxInst_13_n7 ;
    wire SubCellInst_SboxInst_13_n6 ;
    wire SubCellInst_SboxInst_13_n5 ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_n2 ;
    wire SubCellInst_SboxInst_13_n1 ;
    wire SubCellInst_SboxInst_14_n15 ;
    wire SubCellInst_SboxInst_14_n14 ;
    wire SubCellInst_SboxInst_14_n13 ;
    wire SubCellInst_SboxInst_14_n10 ;
    wire SubCellInst_SboxInst_14_n9 ;
    wire SubCellInst_SboxInst_14_n8 ;
    wire SubCellInst_SboxInst_14_n7 ;
    wire SubCellInst_SboxInst_14_n6 ;
    wire SubCellInst_SboxInst_14_n5 ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_n2 ;
    wire SubCellInst_SboxInst_14_n1 ;
    wire SubCellInst_SboxInst_15_n15 ;
    wire SubCellInst_SboxInst_15_n14 ;
    wire SubCellInst_SboxInst_15_n13 ;
    wire SubCellInst_SboxInst_15_n10 ;
    wire SubCellInst_SboxInst_15_n9 ;
    wire SubCellInst_SboxInst_15_n8 ;
    wire SubCellInst_SboxInst_15_n7 ;
    wire SubCellInst_SboxInst_15_n6 ;
    wire SubCellInst_SboxInst_15_n5 ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_n2 ;
    wire SubCellInst_SboxInst_15_n1 ;
    wire KeyMUX_MUXInst_0_U1_Y ;
    wire KeyMUX_MUXInst_0_U1_X ;
    wire KeyMUX_MUXInst_1_U1_Y ;
    wire KeyMUX_MUXInst_1_U1_X ;
    wire KeyMUX_MUXInst_2_U1_Y ;
    wire KeyMUX_MUXInst_2_U1_X ;
    wire KeyMUX_MUXInst_3_U1_Y ;
    wire KeyMUX_MUXInst_3_U1_X ;
    wire KeyMUX_MUXInst_4_U1_Y ;
    wire KeyMUX_MUXInst_4_U1_X ;
    wire KeyMUX_MUXInst_5_U1_Y ;
    wire KeyMUX_MUXInst_5_U1_X ;
    wire KeyMUX_MUXInst_6_U1_Y ;
    wire KeyMUX_MUXInst_6_U1_X ;
    wire KeyMUX_MUXInst_7_U1_Y ;
    wire KeyMUX_MUXInst_7_U1_X ;
    wire KeyMUX_MUXInst_8_U1_Y ;
    wire KeyMUX_MUXInst_8_U1_X ;
    wire KeyMUX_MUXInst_9_U1_Y ;
    wire KeyMUX_MUXInst_9_U1_X ;
    wire KeyMUX_MUXInst_10_U1_Y ;
    wire KeyMUX_MUXInst_10_U1_X ;
    wire KeyMUX_MUXInst_11_U1_Y ;
    wire KeyMUX_MUXInst_11_U1_X ;
    wire KeyMUX_MUXInst_12_U1_Y ;
    wire KeyMUX_MUXInst_12_U1_X ;
    wire KeyMUX_MUXInst_13_U1_Y ;
    wire KeyMUX_MUXInst_13_U1_X ;
    wire KeyMUX_MUXInst_14_U1_Y ;
    wire KeyMUX_MUXInst_14_U1_X ;
    wire KeyMUX_MUXInst_15_U1_Y ;
    wire KeyMUX_MUXInst_15_U1_X ;
    wire KeyMUX_MUXInst_16_U1_Y ;
    wire KeyMUX_MUXInst_16_U1_X ;
    wire KeyMUX_MUXInst_17_U1_Y ;
    wire KeyMUX_MUXInst_17_U1_X ;
    wire KeyMUX_MUXInst_18_U1_Y ;
    wire KeyMUX_MUXInst_18_U1_X ;
    wire KeyMUX_MUXInst_19_U1_Y ;
    wire KeyMUX_MUXInst_19_U1_X ;
    wire KeyMUX_MUXInst_20_U1_Y ;
    wire KeyMUX_MUXInst_20_U1_X ;
    wire KeyMUX_MUXInst_21_U1_Y ;
    wire KeyMUX_MUXInst_21_U1_X ;
    wire KeyMUX_MUXInst_22_U1_Y ;
    wire KeyMUX_MUXInst_22_U1_X ;
    wire KeyMUX_MUXInst_23_U1_Y ;
    wire KeyMUX_MUXInst_23_U1_X ;
    wire KeyMUX_MUXInst_24_U1_Y ;
    wire KeyMUX_MUXInst_24_U1_X ;
    wire KeyMUX_MUXInst_25_U1_Y ;
    wire KeyMUX_MUXInst_25_U1_X ;
    wire KeyMUX_MUXInst_26_U1_Y ;
    wire KeyMUX_MUXInst_26_U1_X ;
    wire KeyMUX_MUXInst_27_U1_Y ;
    wire KeyMUX_MUXInst_27_U1_X ;
    wire KeyMUX_MUXInst_28_U1_Y ;
    wire KeyMUX_MUXInst_28_U1_X ;
    wire KeyMUX_MUXInst_29_U1_Y ;
    wire KeyMUX_MUXInst_29_U1_X ;
    wire KeyMUX_MUXInst_30_U1_Y ;
    wire KeyMUX_MUXInst_30_U1_X ;
    wire KeyMUX_MUXInst_31_U1_Y ;
    wire KeyMUX_MUXInst_31_U1_X ;
    wire KeyMUX_MUXInst_32_U1_Y ;
    wire KeyMUX_MUXInst_32_U1_X ;
    wire KeyMUX_MUXInst_33_U1_Y ;
    wire KeyMUX_MUXInst_33_U1_X ;
    wire KeyMUX_MUXInst_34_U1_Y ;
    wire KeyMUX_MUXInst_34_U1_X ;
    wire KeyMUX_MUXInst_35_U1_Y ;
    wire KeyMUX_MUXInst_35_U1_X ;
    wire KeyMUX_MUXInst_36_U1_Y ;
    wire KeyMUX_MUXInst_36_U1_X ;
    wire KeyMUX_MUXInst_37_U1_Y ;
    wire KeyMUX_MUXInst_37_U1_X ;
    wire KeyMUX_MUXInst_38_U1_Y ;
    wire KeyMUX_MUXInst_38_U1_X ;
    wire KeyMUX_MUXInst_39_U1_Y ;
    wire KeyMUX_MUXInst_39_U1_X ;
    wire KeyMUX_MUXInst_40_U1_Y ;
    wire KeyMUX_MUXInst_40_U1_X ;
    wire KeyMUX_MUXInst_41_U1_Y ;
    wire KeyMUX_MUXInst_41_U1_X ;
    wire KeyMUX_MUXInst_42_U1_Y ;
    wire KeyMUX_MUXInst_42_U1_X ;
    wire KeyMUX_MUXInst_43_U1_Y ;
    wire KeyMUX_MUXInst_43_U1_X ;
    wire KeyMUX_MUXInst_44_U1_Y ;
    wire KeyMUX_MUXInst_44_U1_X ;
    wire KeyMUX_MUXInst_45_U1_Y ;
    wire KeyMUX_MUXInst_45_U1_X ;
    wire KeyMUX_MUXInst_46_U1_Y ;
    wire KeyMUX_MUXInst_46_U1_X ;
    wire KeyMUX_MUXInst_47_U1_Y ;
    wire KeyMUX_MUXInst_47_U1_X ;
    wire KeyMUX_MUXInst_48_U1_Y ;
    wire KeyMUX_MUXInst_48_U1_X ;
    wire KeyMUX_MUXInst_49_U1_Y ;
    wire KeyMUX_MUXInst_49_U1_X ;
    wire KeyMUX_MUXInst_50_U1_Y ;
    wire KeyMUX_MUXInst_50_U1_X ;
    wire KeyMUX_MUXInst_51_U1_Y ;
    wire KeyMUX_MUXInst_51_U1_X ;
    wire KeyMUX_MUXInst_52_U1_Y ;
    wire KeyMUX_MUXInst_52_U1_X ;
    wire KeyMUX_MUXInst_53_U1_Y ;
    wire KeyMUX_MUXInst_53_U1_X ;
    wire KeyMUX_MUXInst_54_U1_Y ;
    wire KeyMUX_MUXInst_54_U1_X ;
    wire KeyMUX_MUXInst_55_U1_Y ;
    wire KeyMUX_MUXInst_55_U1_X ;
    wire KeyMUX_MUXInst_56_U1_Y ;
    wire KeyMUX_MUXInst_56_U1_X ;
    wire KeyMUX_MUXInst_57_U1_Y ;
    wire KeyMUX_MUXInst_57_U1_X ;
    wire KeyMUX_MUXInst_58_U1_Y ;
    wire KeyMUX_MUXInst_58_U1_X ;
    wire KeyMUX_MUXInst_59_U1_Y ;
    wire KeyMUX_MUXInst_59_U1_X ;
    wire KeyMUX_MUXInst_60_U1_Y ;
    wire KeyMUX_MUXInst_60_U1_X ;
    wire KeyMUX_MUXInst_61_U1_Y ;
    wire KeyMUX_MUXInst_61_U1_X ;
    wire KeyMUX_MUXInst_62_U1_Y ;
    wire KeyMUX_MUXInst_62_U1_X ;
    wire KeyMUX_MUXInst_63_U1_Y ;
    wire KeyMUX_MUXInst_63_U1_X ;
    wire FSMSignalsInst_n5 ;
    wire FSMSignalsInst_n4 ;
    wire FSMSignalsInst_n3 ;
    wire FSMSignalsInst_n2 ;
    wire FSMSignalsInst_n1 ;
    wire [63:0] Feedback ;
    wire [63:32] MCInput ;
    wire [63:0] MCOutput ;
    wire [63:0] SelectedKey ;
    wire [1:0] selects ;
    wire [6:0] FSMReg ;
    wire [5:0] FSMUpdate ;
    wire [1:0] selectsReg ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;

    /* cells in depth 0 */
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_0_U1_XOR1_U1 ( .A0_t (Feedback[0]), .A0_f (new_AGEMA_signal_3223), .A1_t (new_AGEMA_signal_3224), .A1_f (new_AGEMA_signal_3225), .B0_t (Input_s0_t[0]), .B0_f (Input_s0_f[0]), .B1_t (Input_s1_t[0]), .B1_f (Input_s1_f[0]), .Z0_t (InputMUX_MUXInst_0_U1_X), .Z0_f (new_AGEMA_signal_3323), .Z1_t (new_AGEMA_signal_3324), .Z1_f (new_AGEMA_signal_3325) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_0_U1_X), .B0_f (new_AGEMA_signal_3323), .B1_t (new_AGEMA_signal_3324), .B1_f (new_AGEMA_signal_3325), .Z0_t (InputMUX_MUXInst_0_U1_Y), .Z0_f (new_AGEMA_signal_3609), .Z1_t (new_AGEMA_signal_3610), .Z1_f (new_AGEMA_signal_3611) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_0_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_0_U1_Y), .A0_f (new_AGEMA_signal_3609), .A1_t (new_AGEMA_signal_3610), .A1_f (new_AGEMA_signal_3611), .B0_t (Feedback[0]), .B0_f (new_AGEMA_signal_3223), .B1_t (new_AGEMA_signal_3224), .B1_f (new_AGEMA_signal_3225), .Z0_t (MCOutput[0]), .Z0_f (new_AGEMA_signal_3801), .Z1_t (new_AGEMA_signal_3802), .Z1_f (new_AGEMA_signal_3803) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_1_U1_XOR1_U1 ( .A0_t (Feedback[1]), .A0_f (new_AGEMA_signal_2649), .A1_t (new_AGEMA_signal_2650), .A1_f (new_AGEMA_signal_2651), .B0_t (Input_s0_t[1]), .B0_f (Input_s0_f[1]), .B1_t (Input_s1_t[1]), .B1_f (Input_s1_f[1]), .Z0_t (InputMUX_MUXInst_1_U1_X), .Z0_f (new_AGEMA_signal_3034), .Z1_t (new_AGEMA_signal_3035), .Z1_f (new_AGEMA_signal_3036) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_1_U1_X), .B0_f (new_AGEMA_signal_3034), .B1_t (new_AGEMA_signal_3035), .B1_f (new_AGEMA_signal_3036), .Z0_t (InputMUX_MUXInst_1_U1_Y), .Z0_f (new_AGEMA_signal_3326), .Z1_t (new_AGEMA_signal_3327), .Z1_f (new_AGEMA_signal_3328) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_1_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_1_U1_Y), .A0_f (new_AGEMA_signal_3326), .A1_t (new_AGEMA_signal_3327), .A1_f (new_AGEMA_signal_3328), .B0_t (Feedback[1]), .B0_f (new_AGEMA_signal_2649), .B1_t (new_AGEMA_signal_2650), .B1_f (new_AGEMA_signal_2651), .Z0_t (MCOutput[1]), .Z0_f (new_AGEMA_signal_3612), .Z1_t (new_AGEMA_signal_3613), .Z1_f (new_AGEMA_signal_3614) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_2_U1_XOR1_U1 ( .A0_t (Feedback[2]), .A0_f (new_AGEMA_signal_3226), .A1_t (new_AGEMA_signal_3227), .A1_f (new_AGEMA_signal_3228), .B0_t (Input_s0_t[2]), .B0_f (Input_s0_f[2]), .B1_t (Input_s1_t[2]), .B1_f (Input_s1_f[2]), .Z0_t (InputMUX_MUXInst_2_U1_X), .Z0_f (new_AGEMA_signal_3332), .Z1_t (new_AGEMA_signal_3333), .Z1_f (new_AGEMA_signal_3334) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_2_U1_X), .B0_f (new_AGEMA_signal_3332), .B1_t (new_AGEMA_signal_3333), .B1_f (new_AGEMA_signal_3334), .Z0_t (InputMUX_MUXInst_2_U1_Y), .Z0_f (new_AGEMA_signal_3615), .Z1_t (new_AGEMA_signal_3616), .Z1_f (new_AGEMA_signal_3617) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_2_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_2_U1_Y), .A0_f (new_AGEMA_signal_3615), .A1_t (new_AGEMA_signal_3616), .A1_f (new_AGEMA_signal_3617), .B0_t (Feedback[2]), .B0_f (new_AGEMA_signal_3226), .B1_t (new_AGEMA_signal_3227), .B1_f (new_AGEMA_signal_3228), .Z0_t (MCOutput[2]), .Z0_f (new_AGEMA_signal_3804), .Z1_t (new_AGEMA_signal_3805), .Z1_f (new_AGEMA_signal_3806) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_3_U1_XOR1_U1 ( .A0_t (Feedback[3]), .A0_f (new_AGEMA_signal_2655), .A1_t (new_AGEMA_signal_2656), .A1_f (new_AGEMA_signal_2657), .B0_t (Input_s0_t[3]), .B0_f (Input_s0_f[3]), .B1_t (Input_s1_t[3]), .B1_f (Input_s1_f[3]), .Z0_t (InputMUX_MUXInst_3_U1_X), .Z0_f (new_AGEMA_signal_3040), .Z1_t (new_AGEMA_signal_3041), .Z1_f (new_AGEMA_signal_3042) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_3_U1_X), .B0_f (new_AGEMA_signal_3040), .B1_t (new_AGEMA_signal_3041), .B1_f (new_AGEMA_signal_3042), .Z0_t (InputMUX_MUXInst_3_U1_Y), .Z0_f (new_AGEMA_signal_3335), .Z1_t (new_AGEMA_signal_3336), .Z1_f (new_AGEMA_signal_3337) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_3_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_3_U1_Y), .A0_f (new_AGEMA_signal_3335), .A1_t (new_AGEMA_signal_3336), .A1_f (new_AGEMA_signal_3337), .B0_t (Feedback[3]), .B0_f (new_AGEMA_signal_2655), .B1_t (new_AGEMA_signal_2656), .B1_f (new_AGEMA_signal_2657), .Z0_t (MCOutput[3]), .Z0_f (new_AGEMA_signal_3618), .Z1_t (new_AGEMA_signal_3619), .Z1_f (new_AGEMA_signal_3620) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_4_U1_XOR1_U1 ( .A0_t (Feedback[4]), .A0_f (new_AGEMA_signal_3229), .A1_t (new_AGEMA_signal_3230), .A1_f (new_AGEMA_signal_3231), .B0_t (Input_s0_t[4]), .B0_f (Input_s0_f[4]), .B1_t (Input_s1_t[4]), .B1_f (Input_s1_f[4]), .Z0_t (InputMUX_MUXInst_4_U1_X), .Z0_f (new_AGEMA_signal_3341), .Z1_t (new_AGEMA_signal_3342), .Z1_f (new_AGEMA_signal_3343) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_4_U1_X), .B0_f (new_AGEMA_signal_3341), .B1_t (new_AGEMA_signal_3342), .B1_f (new_AGEMA_signal_3343), .Z0_t (InputMUX_MUXInst_4_U1_Y), .Z0_f (new_AGEMA_signal_3621), .Z1_t (new_AGEMA_signal_3622), .Z1_f (new_AGEMA_signal_3623) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_4_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_4_U1_Y), .A0_f (new_AGEMA_signal_3621), .A1_t (new_AGEMA_signal_3622), .A1_f (new_AGEMA_signal_3623), .B0_t (Feedback[4]), .B0_f (new_AGEMA_signal_3229), .B1_t (new_AGEMA_signal_3230), .B1_f (new_AGEMA_signal_3231), .Z0_t (MCOutput[4]), .Z0_f (new_AGEMA_signal_3807), .Z1_t (new_AGEMA_signal_3808), .Z1_f (new_AGEMA_signal_3809) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_5_U1_XOR1_U1 ( .A0_t (Feedback[5]), .A0_f (new_AGEMA_signal_2661), .A1_t (new_AGEMA_signal_2662), .A1_f (new_AGEMA_signal_2663), .B0_t (Input_s0_t[5]), .B0_f (Input_s0_f[5]), .B1_t (Input_s1_t[5]), .B1_f (Input_s1_f[5]), .Z0_t (InputMUX_MUXInst_5_U1_X), .Z0_f (new_AGEMA_signal_3046), .Z1_t (new_AGEMA_signal_3047), .Z1_f (new_AGEMA_signal_3048) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_5_U1_X), .B0_f (new_AGEMA_signal_3046), .B1_t (new_AGEMA_signal_3047), .B1_f (new_AGEMA_signal_3048), .Z0_t (InputMUX_MUXInst_5_U1_Y), .Z0_f (new_AGEMA_signal_3344), .Z1_t (new_AGEMA_signal_3345), .Z1_f (new_AGEMA_signal_3346) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_5_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_5_U1_Y), .A0_f (new_AGEMA_signal_3344), .A1_t (new_AGEMA_signal_3345), .A1_f (new_AGEMA_signal_3346), .B0_t (Feedback[5]), .B0_f (new_AGEMA_signal_2661), .B1_t (new_AGEMA_signal_2662), .B1_f (new_AGEMA_signal_2663), .Z0_t (MCOutput[5]), .Z0_f (new_AGEMA_signal_3624), .Z1_t (new_AGEMA_signal_3625), .Z1_f (new_AGEMA_signal_3626) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_6_U1_XOR1_U1 ( .A0_t (Feedback[6]), .A0_f (new_AGEMA_signal_3232), .A1_t (new_AGEMA_signal_3233), .A1_f (new_AGEMA_signal_3234), .B0_t (Input_s0_t[6]), .B0_f (Input_s0_f[6]), .B1_t (Input_s1_t[6]), .B1_f (Input_s1_f[6]), .Z0_t (InputMUX_MUXInst_6_U1_X), .Z0_f (new_AGEMA_signal_3350), .Z1_t (new_AGEMA_signal_3351), .Z1_f (new_AGEMA_signal_3352) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_6_U1_X), .B0_f (new_AGEMA_signal_3350), .B1_t (new_AGEMA_signal_3351), .B1_f (new_AGEMA_signal_3352), .Z0_t (InputMUX_MUXInst_6_U1_Y), .Z0_f (new_AGEMA_signal_3627), .Z1_t (new_AGEMA_signal_3628), .Z1_f (new_AGEMA_signal_3629) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_6_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_6_U1_Y), .A0_f (new_AGEMA_signal_3627), .A1_t (new_AGEMA_signal_3628), .A1_f (new_AGEMA_signal_3629), .B0_t (Feedback[6]), .B0_f (new_AGEMA_signal_3232), .B1_t (new_AGEMA_signal_3233), .B1_f (new_AGEMA_signal_3234), .Z0_t (MCOutput[6]), .Z0_f (new_AGEMA_signal_3810), .Z1_t (new_AGEMA_signal_3811), .Z1_f (new_AGEMA_signal_3812) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_7_U1_XOR1_U1 ( .A0_t (Feedback[7]), .A0_f (new_AGEMA_signal_2667), .A1_t (new_AGEMA_signal_2668), .A1_f (new_AGEMA_signal_2669), .B0_t (Input_s0_t[7]), .B0_f (Input_s0_f[7]), .B1_t (Input_s1_t[7]), .B1_f (Input_s1_f[7]), .Z0_t (InputMUX_MUXInst_7_U1_X), .Z0_f (new_AGEMA_signal_3052), .Z1_t (new_AGEMA_signal_3053), .Z1_f (new_AGEMA_signal_3054) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_7_U1_X), .B0_f (new_AGEMA_signal_3052), .B1_t (new_AGEMA_signal_3053), .B1_f (new_AGEMA_signal_3054), .Z0_t (InputMUX_MUXInst_7_U1_Y), .Z0_f (new_AGEMA_signal_3353), .Z1_t (new_AGEMA_signal_3354), .Z1_f (new_AGEMA_signal_3355) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_7_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_7_U1_Y), .A0_f (new_AGEMA_signal_3353), .A1_t (new_AGEMA_signal_3354), .A1_f (new_AGEMA_signal_3355), .B0_t (Feedback[7]), .B0_f (new_AGEMA_signal_2667), .B1_t (new_AGEMA_signal_2668), .B1_f (new_AGEMA_signal_2669), .Z0_t (MCOutput[7]), .Z0_f (new_AGEMA_signal_3630), .Z1_t (new_AGEMA_signal_3631), .Z1_f (new_AGEMA_signal_3632) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_8_U1_XOR1_U1 ( .A0_t (Feedback[8]), .A0_f (new_AGEMA_signal_3235), .A1_t (new_AGEMA_signal_3236), .A1_f (new_AGEMA_signal_3237), .B0_t (Input_s0_t[8]), .B0_f (Input_s0_f[8]), .B1_t (Input_s1_t[8]), .B1_f (Input_s1_f[8]), .Z0_t (InputMUX_MUXInst_8_U1_X), .Z0_f (new_AGEMA_signal_3359), .Z1_t (new_AGEMA_signal_3360), .Z1_f (new_AGEMA_signal_3361) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_8_U1_X), .B0_f (new_AGEMA_signal_3359), .B1_t (new_AGEMA_signal_3360), .B1_f (new_AGEMA_signal_3361), .Z0_t (InputMUX_MUXInst_8_U1_Y), .Z0_f (new_AGEMA_signal_3633), .Z1_t (new_AGEMA_signal_3634), .Z1_f (new_AGEMA_signal_3635) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_8_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_8_U1_Y), .A0_f (new_AGEMA_signal_3633), .A1_t (new_AGEMA_signal_3634), .A1_f (new_AGEMA_signal_3635), .B0_t (Feedback[8]), .B0_f (new_AGEMA_signal_3235), .B1_t (new_AGEMA_signal_3236), .B1_f (new_AGEMA_signal_3237), .Z0_t (MCOutput[8]), .Z0_f (new_AGEMA_signal_3813), .Z1_t (new_AGEMA_signal_3814), .Z1_f (new_AGEMA_signal_3815) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_9_U1_XOR1_U1 ( .A0_t (Feedback[9]), .A0_f (new_AGEMA_signal_2673), .A1_t (new_AGEMA_signal_2674), .A1_f (new_AGEMA_signal_2675), .B0_t (Input_s0_t[9]), .B0_f (Input_s0_f[9]), .B1_t (Input_s1_t[9]), .B1_f (Input_s1_f[9]), .Z0_t (InputMUX_MUXInst_9_U1_X), .Z0_f (new_AGEMA_signal_3058), .Z1_t (new_AGEMA_signal_3059), .Z1_f (new_AGEMA_signal_3060) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_9_U1_X), .B0_f (new_AGEMA_signal_3058), .B1_t (new_AGEMA_signal_3059), .B1_f (new_AGEMA_signal_3060), .Z0_t (InputMUX_MUXInst_9_U1_Y), .Z0_f (new_AGEMA_signal_3362), .Z1_t (new_AGEMA_signal_3363), .Z1_f (new_AGEMA_signal_3364) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_9_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_9_U1_Y), .A0_f (new_AGEMA_signal_3362), .A1_t (new_AGEMA_signal_3363), .A1_f (new_AGEMA_signal_3364), .B0_t (Feedback[9]), .B0_f (new_AGEMA_signal_2673), .B1_t (new_AGEMA_signal_2674), .B1_f (new_AGEMA_signal_2675), .Z0_t (MCOutput[9]), .Z0_f (new_AGEMA_signal_3636), .Z1_t (new_AGEMA_signal_3637), .Z1_f (new_AGEMA_signal_3638) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_10_U1_XOR1_U1 ( .A0_t (Feedback[10]), .A0_f (new_AGEMA_signal_3238), .A1_t (new_AGEMA_signal_3239), .A1_f (new_AGEMA_signal_3240), .B0_t (Input_s0_t[10]), .B0_f (Input_s0_f[10]), .B1_t (Input_s1_t[10]), .B1_f (Input_s1_f[10]), .Z0_t (InputMUX_MUXInst_10_U1_X), .Z0_f (new_AGEMA_signal_3368), .Z1_t (new_AGEMA_signal_3369), .Z1_f (new_AGEMA_signal_3370) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_10_U1_X), .B0_f (new_AGEMA_signal_3368), .B1_t (new_AGEMA_signal_3369), .B1_f (new_AGEMA_signal_3370), .Z0_t (InputMUX_MUXInst_10_U1_Y), .Z0_f (new_AGEMA_signal_3639), .Z1_t (new_AGEMA_signal_3640), .Z1_f (new_AGEMA_signal_3641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_10_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_10_U1_Y), .A0_f (new_AGEMA_signal_3639), .A1_t (new_AGEMA_signal_3640), .A1_f (new_AGEMA_signal_3641), .B0_t (Feedback[10]), .B0_f (new_AGEMA_signal_3238), .B1_t (new_AGEMA_signal_3239), .B1_f (new_AGEMA_signal_3240), .Z0_t (MCOutput[10]), .Z0_f (new_AGEMA_signal_3816), .Z1_t (new_AGEMA_signal_3817), .Z1_f (new_AGEMA_signal_3818) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_11_U1_XOR1_U1 ( .A0_t (Feedback[11]), .A0_f (new_AGEMA_signal_2679), .A1_t (new_AGEMA_signal_2680), .A1_f (new_AGEMA_signal_2681), .B0_t (Input_s0_t[11]), .B0_f (Input_s0_f[11]), .B1_t (Input_s1_t[11]), .B1_f (Input_s1_f[11]), .Z0_t (InputMUX_MUXInst_11_U1_X), .Z0_f (new_AGEMA_signal_3064), .Z1_t (new_AGEMA_signal_3065), .Z1_f (new_AGEMA_signal_3066) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_11_U1_X), .B0_f (new_AGEMA_signal_3064), .B1_t (new_AGEMA_signal_3065), .B1_f (new_AGEMA_signal_3066), .Z0_t (InputMUX_MUXInst_11_U1_Y), .Z0_f (new_AGEMA_signal_3371), .Z1_t (new_AGEMA_signal_3372), .Z1_f (new_AGEMA_signal_3373) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_11_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_11_U1_Y), .A0_f (new_AGEMA_signal_3371), .A1_t (new_AGEMA_signal_3372), .A1_f (new_AGEMA_signal_3373), .B0_t (Feedback[11]), .B0_f (new_AGEMA_signal_2679), .B1_t (new_AGEMA_signal_2680), .B1_f (new_AGEMA_signal_2681), .Z0_t (MCOutput[11]), .Z0_f (new_AGEMA_signal_3642), .Z1_t (new_AGEMA_signal_3643), .Z1_f (new_AGEMA_signal_3644) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_12_U1_XOR1_U1 ( .A0_t (Feedback[12]), .A0_f (new_AGEMA_signal_3241), .A1_t (new_AGEMA_signal_3242), .A1_f (new_AGEMA_signal_3243), .B0_t (Input_s0_t[12]), .B0_f (Input_s0_f[12]), .B1_t (Input_s1_t[12]), .B1_f (Input_s1_f[12]), .Z0_t (InputMUX_MUXInst_12_U1_X), .Z0_f (new_AGEMA_signal_3377), .Z1_t (new_AGEMA_signal_3378), .Z1_f (new_AGEMA_signal_3379) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_12_U1_X), .B0_f (new_AGEMA_signal_3377), .B1_t (new_AGEMA_signal_3378), .B1_f (new_AGEMA_signal_3379), .Z0_t (InputMUX_MUXInst_12_U1_Y), .Z0_f (new_AGEMA_signal_3645), .Z1_t (new_AGEMA_signal_3646), .Z1_f (new_AGEMA_signal_3647) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_12_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_12_U1_Y), .A0_f (new_AGEMA_signal_3645), .A1_t (new_AGEMA_signal_3646), .A1_f (new_AGEMA_signal_3647), .B0_t (Feedback[12]), .B0_f (new_AGEMA_signal_3241), .B1_t (new_AGEMA_signal_3242), .B1_f (new_AGEMA_signal_3243), .Z0_t (MCOutput[12]), .Z0_f (new_AGEMA_signal_3819), .Z1_t (new_AGEMA_signal_3820), .Z1_f (new_AGEMA_signal_3821) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_13_U1_XOR1_U1 ( .A0_t (Feedback[13]), .A0_f (new_AGEMA_signal_2685), .A1_t (new_AGEMA_signal_2686), .A1_f (new_AGEMA_signal_2687), .B0_t (Input_s0_t[13]), .B0_f (Input_s0_f[13]), .B1_t (Input_s1_t[13]), .B1_f (Input_s1_f[13]), .Z0_t (InputMUX_MUXInst_13_U1_X), .Z0_f (new_AGEMA_signal_3070), .Z1_t (new_AGEMA_signal_3071), .Z1_f (new_AGEMA_signal_3072) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_13_U1_X), .B0_f (new_AGEMA_signal_3070), .B1_t (new_AGEMA_signal_3071), .B1_f (new_AGEMA_signal_3072), .Z0_t (InputMUX_MUXInst_13_U1_Y), .Z0_f (new_AGEMA_signal_3380), .Z1_t (new_AGEMA_signal_3381), .Z1_f (new_AGEMA_signal_3382) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_13_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_13_U1_Y), .A0_f (new_AGEMA_signal_3380), .A1_t (new_AGEMA_signal_3381), .A1_f (new_AGEMA_signal_3382), .B0_t (Feedback[13]), .B0_f (new_AGEMA_signal_2685), .B1_t (new_AGEMA_signal_2686), .B1_f (new_AGEMA_signal_2687), .Z0_t (MCOutput[13]), .Z0_f (new_AGEMA_signal_3648), .Z1_t (new_AGEMA_signal_3649), .Z1_f (new_AGEMA_signal_3650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_14_U1_XOR1_U1 ( .A0_t (Feedback[14]), .A0_f (new_AGEMA_signal_3244), .A1_t (new_AGEMA_signal_3245), .A1_f (new_AGEMA_signal_3246), .B0_t (Input_s0_t[14]), .B0_f (Input_s0_f[14]), .B1_t (Input_s1_t[14]), .B1_f (Input_s1_f[14]), .Z0_t (InputMUX_MUXInst_14_U1_X), .Z0_f (new_AGEMA_signal_3386), .Z1_t (new_AGEMA_signal_3387), .Z1_f (new_AGEMA_signal_3388) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_14_U1_X), .B0_f (new_AGEMA_signal_3386), .B1_t (new_AGEMA_signal_3387), .B1_f (new_AGEMA_signal_3388), .Z0_t (InputMUX_MUXInst_14_U1_Y), .Z0_f (new_AGEMA_signal_3651), .Z1_t (new_AGEMA_signal_3652), .Z1_f (new_AGEMA_signal_3653) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_14_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_14_U1_Y), .A0_f (new_AGEMA_signal_3651), .A1_t (new_AGEMA_signal_3652), .A1_f (new_AGEMA_signal_3653), .B0_t (Feedback[14]), .B0_f (new_AGEMA_signal_3244), .B1_t (new_AGEMA_signal_3245), .B1_f (new_AGEMA_signal_3246), .Z0_t (MCOutput[14]), .Z0_f (new_AGEMA_signal_3822), .Z1_t (new_AGEMA_signal_3823), .Z1_f (new_AGEMA_signal_3824) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_15_U1_XOR1_U1 ( .A0_t (Feedback[15]), .A0_f (new_AGEMA_signal_2691), .A1_t (new_AGEMA_signal_2692), .A1_f (new_AGEMA_signal_2693), .B0_t (Input_s0_t[15]), .B0_f (Input_s0_f[15]), .B1_t (Input_s1_t[15]), .B1_f (Input_s1_f[15]), .Z0_t (InputMUX_MUXInst_15_U1_X), .Z0_f (new_AGEMA_signal_3076), .Z1_t (new_AGEMA_signal_3077), .Z1_f (new_AGEMA_signal_3078) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_15_U1_X), .B0_f (new_AGEMA_signal_3076), .B1_t (new_AGEMA_signal_3077), .B1_f (new_AGEMA_signal_3078), .Z0_t (InputMUX_MUXInst_15_U1_Y), .Z0_f (new_AGEMA_signal_3389), .Z1_t (new_AGEMA_signal_3390), .Z1_f (new_AGEMA_signal_3391) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_15_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_15_U1_Y), .A0_f (new_AGEMA_signal_3389), .A1_t (new_AGEMA_signal_3390), .A1_f (new_AGEMA_signal_3391), .B0_t (Feedback[15]), .B0_f (new_AGEMA_signal_2691), .B1_t (new_AGEMA_signal_2692), .B1_f (new_AGEMA_signal_2693), .Z0_t (MCOutput[15]), .Z0_f (new_AGEMA_signal_3654), .Z1_t (new_AGEMA_signal_3655), .Z1_f (new_AGEMA_signal_3656) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_16_U1_XOR1_U1 ( .A0_t (Feedback[16]), .A0_f (new_AGEMA_signal_3247), .A1_t (new_AGEMA_signal_3248), .A1_f (new_AGEMA_signal_3249), .B0_t (Input_s0_t[16]), .B0_f (Input_s0_f[16]), .B1_t (Input_s1_t[16]), .B1_f (Input_s1_f[16]), .Z0_t (InputMUX_MUXInst_16_U1_X), .Z0_f (new_AGEMA_signal_3395), .Z1_t (new_AGEMA_signal_3396), .Z1_f (new_AGEMA_signal_3397) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_16_U1_X), .B0_f (new_AGEMA_signal_3395), .B1_t (new_AGEMA_signal_3396), .B1_f (new_AGEMA_signal_3397), .Z0_t (InputMUX_MUXInst_16_U1_Y), .Z0_f (new_AGEMA_signal_3657), .Z1_t (new_AGEMA_signal_3658), .Z1_f (new_AGEMA_signal_3659) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_16_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_16_U1_Y), .A0_f (new_AGEMA_signal_3657), .A1_t (new_AGEMA_signal_3658), .A1_f (new_AGEMA_signal_3659), .B0_t (Feedback[16]), .B0_f (new_AGEMA_signal_3247), .B1_t (new_AGEMA_signal_3248), .B1_f (new_AGEMA_signal_3249), .Z0_t (MCOutput[16]), .Z0_f (new_AGEMA_signal_3825), .Z1_t (new_AGEMA_signal_3826), .Z1_f (new_AGEMA_signal_3827) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_17_U1_XOR1_U1 ( .A0_t (Feedback[17]), .A0_f (new_AGEMA_signal_2694), .A1_t (new_AGEMA_signal_2695), .A1_f (new_AGEMA_signal_2696), .B0_t (Input_s0_t[17]), .B0_f (Input_s0_f[17]), .B1_t (Input_s1_t[17]), .B1_f (Input_s1_f[17]), .Z0_t (InputMUX_MUXInst_17_U1_X), .Z0_f (new_AGEMA_signal_3082), .Z1_t (new_AGEMA_signal_3083), .Z1_f (new_AGEMA_signal_3084) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_17_U1_X), .B0_f (new_AGEMA_signal_3082), .B1_t (new_AGEMA_signal_3083), .B1_f (new_AGEMA_signal_3084), .Z0_t (InputMUX_MUXInst_17_U1_Y), .Z0_f (new_AGEMA_signal_3398), .Z1_t (new_AGEMA_signal_3399), .Z1_f (new_AGEMA_signal_3400) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_17_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_17_U1_Y), .A0_f (new_AGEMA_signal_3398), .A1_t (new_AGEMA_signal_3399), .A1_f (new_AGEMA_signal_3400), .B0_t (Feedback[17]), .B0_f (new_AGEMA_signal_2694), .B1_t (new_AGEMA_signal_2695), .B1_f (new_AGEMA_signal_2696), .Z0_t (MCOutput[17]), .Z0_f (new_AGEMA_signal_3660), .Z1_t (new_AGEMA_signal_3661), .Z1_f (new_AGEMA_signal_3662) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_18_U1_XOR1_U1 ( .A0_t (Feedback[18]), .A0_f (new_AGEMA_signal_3250), .A1_t (new_AGEMA_signal_3251), .A1_f (new_AGEMA_signal_3252), .B0_t (Input_s0_t[18]), .B0_f (Input_s0_f[18]), .B1_t (Input_s1_t[18]), .B1_f (Input_s1_f[18]), .Z0_t (InputMUX_MUXInst_18_U1_X), .Z0_f (new_AGEMA_signal_3404), .Z1_t (new_AGEMA_signal_3405), .Z1_f (new_AGEMA_signal_3406) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_18_U1_X), .B0_f (new_AGEMA_signal_3404), .B1_t (new_AGEMA_signal_3405), .B1_f (new_AGEMA_signal_3406), .Z0_t (InputMUX_MUXInst_18_U1_Y), .Z0_f (new_AGEMA_signal_3663), .Z1_t (new_AGEMA_signal_3664), .Z1_f (new_AGEMA_signal_3665) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_18_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_18_U1_Y), .A0_f (new_AGEMA_signal_3663), .A1_t (new_AGEMA_signal_3664), .A1_f (new_AGEMA_signal_3665), .B0_t (Feedback[18]), .B0_f (new_AGEMA_signal_3250), .B1_t (new_AGEMA_signal_3251), .B1_f (new_AGEMA_signal_3252), .Z0_t (MCOutput[18]), .Z0_f (new_AGEMA_signal_3828), .Z1_t (new_AGEMA_signal_3829), .Z1_f (new_AGEMA_signal_3830) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_19_U1_XOR1_U1 ( .A0_t (Feedback[19]), .A0_f (new_AGEMA_signal_2697), .A1_t (new_AGEMA_signal_2698), .A1_f (new_AGEMA_signal_2699), .B0_t (Input_s0_t[19]), .B0_f (Input_s0_f[19]), .B1_t (Input_s1_t[19]), .B1_f (Input_s1_f[19]), .Z0_t (InputMUX_MUXInst_19_U1_X), .Z0_f (new_AGEMA_signal_3088), .Z1_t (new_AGEMA_signal_3089), .Z1_f (new_AGEMA_signal_3090) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_19_U1_X), .B0_f (new_AGEMA_signal_3088), .B1_t (new_AGEMA_signal_3089), .B1_f (new_AGEMA_signal_3090), .Z0_t (InputMUX_MUXInst_19_U1_Y), .Z0_f (new_AGEMA_signal_3407), .Z1_t (new_AGEMA_signal_3408), .Z1_f (new_AGEMA_signal_3409) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_19_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_19_U1_Y), .A0_f (new_AGEMA_signal_3407), .A1_t (new_AGEMA_signal_3408), .A1_f (new_AGEMA_signal_3409), .B0_t (Feedback[19]), .B0_f (new_AGEMA_signal_2697), .B1_t (new_AGEMA_signal_2698), .B1_f (new_AGEMA_signal_2699), .Z0_t (MCOutput[19]), .Z0_f (new_AGEMA_signal_3666), .Z1_t (new_AGEMA_signal_3667), .Z1_f (new_AGEMA_signal_3668) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_20_U1_XOR1_U1 ( .A0_t (Feedback[20]), .A0_f (new_AGEMA_signal_3253), .A1_t (new_AGEMA_signal_3254), .A1_f (new_AGEMA_signal_3255), .B0_t (Input_s0_t[20]), .B0_f (Input_s0_f[20]), .B1_t (Input_s1_t[20]), .B1_f (Input_s1_f[20]), .Z0_t (InputMUX_MUXInst_20_U1_X), .Z0_f (new_AGEMA_signal_3413), .Z1_t (new_AGEMA_signal_3414), .Z1_f (new_AGEMA_signal_3415) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_20_U1_X), .B0_f (new_AGEMA_signal_3413), .B1_t (new_AGEMA_signal_3414), .B1_f (new_AGEMA_signal_3415), .Z0_t (InputMUX_MUXInst_20_U1_Y), .Z0_f (new_AGEMA_signal_3669), .Z1_t (new_AGEMA_signal_3670), .Z1_f (new_AGEMA_signal_3671) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_20_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_20_U1_Y), .A0_f (new_AGEMA_signal_3669), .A1_t (new_AGEMA_signal_3670), .A1_f (new_AGEMA_signal_3671), .B0_t (Feedback[20]), .B0_f (new_AGEMA_signal_3253), .B1_t (new_AGEMA_signal_3254), .B1_f (new_AGEMA_signal_3255), .Z0_t (MCOutput[20]), .Z0_f (new_AGEMA_signal_3831), .Z1_t (new_AGEMA_signal_3832), .Z1_f (new_AGEMA_signal_3833) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_21_U1_XOR1_U1 ( .A0_t (Feedback[21]), .A0_f (new_AGEMA_signal_2706), .A1_t (new_AGEMA_signal_2707), .A1_f (new_AGEMA_signal_2708), .B0_t (Input_s0_t[21]), .B0_f (Input_s0_f[21]), .B1_t (Input_s1_t[21]), .B1_f (Input_s1_f[21]), .Z0_t (InputMUX_MUXInst_21_U1_X), .Z0_f (new_AGEMA_signal_3094), .Z1_t (new_AGEMA_signal_3095), .Z1_f (new_AGEMA_signal_3096) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_21_U1_X), .B0_f (new_AGEMA_signal_3094), .B1_t (new_AGEMA_signal_3095), .B1_f (new_AGEMA_signal_3096), .Z0_t (InputMUX_MUXInst_21_U1_Y), .Z0_f (new_AGEMA_signal_3416), .Z1_t (new_AGEMA_signal_3417), .Z1_f (new_AGEMA_signal_3418) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_21_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_21_U1_Y), .A0_f (new_AGEMA_signal_3416), .A1_t (new_AGEMA_signal_3417), .A1_f (new_AGEMA_signal_3418), .B0_t (Feedback[21]), .B0_f (new_AGEMA_signal_2706), .B1_t (new_AGEMA_signal_2707), .B1_f (new_AGEMA_signal_2708), .Z0_t (MCOutput[21]), .Z0_f (new_AGEMA_signal_3672), .Z1_t (new_AGEMA_signal_3673), .Z1_f (new_AGEMA_signal_3674) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_22_U1_XOR1_U1 ( .A0_t (Feedback[22]), .A0_f (new_AGEMA_signal_3256), .A1_t (new_AGEMA_signal_3257), .A1_f (new_AGEMA_signal_3258), .B0_t (Input_s0_t[22]), .B0_f (Input_s0_f[22]), .B1_t (Input_s1_t[22]), .B1_f (Input_s1_f[22]), .Z0_t (InputMUX_MUXInst_22_U1_X), .Z0_f (new_AGEMA_signal_3422), .Z1_t (new_AGEMA_signal_3423), .Z1_f (new_AGEMA_signal_3424) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_22_U1_X), .B0_f (new_AGEMA_signal_3422), .B1_t (new_AGEMA_signal_3423), .B1_f (new_AGEMA_signal_3424), .Z0_t (InputMUX_MUXInst_22_U1_Y), .Z0_f (new_AGEMA_signal_3675), .Z1_t (new_AGEMA_signal_3676), .Z1_f (new_AGEMA_signal_3677) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_22_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_22_U1_Y), .A0_f (new_AGEMA_signal_3675), .A1_t (new_AGEMA_signal_3676), .A1_f (new_AGEMA_signal_3677), .B0_t (Feedback[22]), .B0_f (new_AGEMA_signal_3256), .B1_t (new_AGEMA_signal_3257), .B1_f (new_AGEMA_signal_3258), .Z0_t (MCOutput[22]), .Z0_f (new_AGEMA_signal_3834), .Z1_t (new_AGEMA_signal_3835), .Z1_f (new_AGEMA_signal_3836) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_23_U1_XOR1_U1 ( .A0_t (Feedback[23]), .A0_f (new_AGEMA_signal_2709), .A1_t (new_AGEMA_signal_2710), .A1_f (new_AGEMA_signal_2711), .B0_t (Input_s0_t[23]), .B0_f (Input_s0_f[23]), .B1_t (Input_s1_t[23]), .B1_f (Input_s1_f[23]), .Z0_t (InputMUX_MUXInst_23_U1_X), .Z0_f (new_AGEMA_signal_3100), .Z1_t (new_AGEMA_signal_3101), .Z1_f (new_AGEMA_signal_3102) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_23_U1_X), .B0_f (new_AGEMA_signal_3100), .B1_t (new_AGEMA_signal_3101), .B1_f (new_AGEMA_signal_3102), .Z0_t (InputMUX_MUXInst_23_U1_Y), .Z0_f (new_AGEMA_signal_3425), .Z1_t (new_AGEMA_signal_3426), .Z1_f (new_AGEMA_signal_3427) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_23_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_23_U1_Y), .A0_f (new_AGEMA_signal_3425), .A1_t (new_AGEMA_signal_3426), .A1_f (new_AGEMA_signal_3427), .B0_t (Feedback[23]), .B0_f (new_AGEMA_signal_2709), .B1_t (new_AGEMA_signal_2710), .B1_f (new_AGEMA_signal_2711), .Z0_t (MCOutput[23]), .Z0_f (new_AGEMA_signal_3678), .Z1_t (new_AGEMA_signal_3679), .Z1_f (new_AGEMA_signal_3680) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_24_U1_XOR1_U1 ( .A0_t (Feedback[24]), .A0_f (new_AGEMA_signal_3259), .A1_t (new_AGEMA_signal_3260), .A1_f (new_AGEMA_signal_3261), .B0_t (Input_s0_t[24]), .B0_f (Input_s0_f[24]), .B1_t (Input_s1_t[24]), .B1_f (Input_s1_f[24]), .Z0_t (InputMUX_MUXInst_24_U1_X), .Z0_f (new_AGEMA_signal_3431), .Z1_t (new_AGEMA_signal_3432), .Z1_f (new_AGEMA_signal_3433) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_24_U1_X), .B0_f (new_AGEMA_signal_3431), .B1_t (new_AGEMA_signal_3432), .B1_f (new_AGEMA_signal_3433), .Z0_t (InputMUX_MUXInst_24_U1_Y), .Z0_f (new_AGEMA_signal_3681), .Z1_t (new_AGEMA_signal_3682), .Z1_f (new_AGEMA_signal_3683) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_24_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_24_U1_Y), .A0_f (new_AGEMA_signal_3681), .A1_t (new_AGEMA_signal_3682), .A1_f (new_AGEMA_signal_3683), .B0_t (Feedback[24]), .B0_f (new_AGEMA_signal_3259), .B1_t (new_AGEMA_signal_3260), .B1_f (new_AGEMA_signal_3261), .Z0_t (MCOutput[24]), .Z0_f (new_AGEMA_signal_3837), .Z1_t (new_AGEMA_signal_3838), .Z1_f (new_AGEMA_signal_3839) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_25_U1_XOR1_U1 ( .A0_t (Feedback[25]), .A0_f (new_AGEMA_signal_2718), .A1_t (new_AGEMA_signal_2719), .A1_f (new_AGEMA_signal_2720), .B0_t (Input_s0_t[25]), .B0_f (Input_s0_f[25]), .B1_t (Input_s1_t[25]), .B1_f (Input_s1_f[25]), .Z0_t (InputMUX_MUXInst_25_U1_X), .Z0_f (new_AGEMA_signal_3106), .Z1_t (new_AGEMA_signal_3107), .Z1_f (new_AGEMA_signal_3108) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_25_U1_X), .B0_f (new_AGEMA_signal_3106), .B1_t (new_AGEMA_signal_3107), .B1_f (new_AGEMA_signal_3108), .Z0_t (InputMUX_MUXInst_25_U1_Y), .Z0_f (new_AGEMA_signal_3434), .Z1_t (new_AGEMA_signal_3435), .Z1_f (new_AGEMA_signal_3436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_25_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_25_U1_Y), .A0_f (new_AGEMA_signal_3434), .A1_t (new_AGEMA_signal_3435), .A1_f (new_AGEMA_signal_3436), .B0_t (Feedback[25]), .B0_f (new_AGEMA_signal_2718), .B1_t (new_AGEMA_signal_2719), .B1_f (new_AGEMA_signal_2720), .Z0_t (MCOutput[25]), .Z0_f (new_AGEMA_signal_3684), .Z1_t (new_AGEMA_signal_3685), .Z1_f (new_AGEMA_signal_3686) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_26_U1_XOR1_U1 ( .A0_t (Feedback[26]), .A0_f (new_AGEMA_signal_3262), .A1_t (new_AGEMA_signal_3263), .A1_f (new_AGEMA_signal_3264), .B0_t (Input_s0_t[26]), .B0_f (Input_s0_f[26]), .B1_t (Input_s1_t[26]), .B1_f (Input_s1_f[26]), .Z0_t (InputMUX_MUXInst_26_U1_X), .Z0_f (new_AGEMA_signal_3440), .Z1_t (new_AGEMA_signal_3441), .Z1_f (new_AGEMA_signal_3442) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_26_U1_X), .B0_f (new_AGEMA_signal_3440), .B1_t (new_AGEMA_signal_3441), .B1_f (new_AGEMA_signal_3442), .Z0_t (InputMUX_MUXInst_26_U1_Y), .Z0_f (new_AGEMA_signal_3687), .Z1_t (new_AGEMA_signal_3688), .Z1_f (new_AGEMA_signal_3689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_26_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_26_U1_Y), .A0_f (new_AGEMA_signal_3687), .A1_t (new_AGEMA_signal_3688), .A1_f (new_AGEMA_signal_3689), .B0_t (Feedback[26]), .B0_f (new_AGEMA_signal_3262), .B1_t (new_AGEMA_signal_3263), .B1_f (new_AGEMA_signal_3264), .Z0_t (MCOutput[26]), .Z0_f (new_AGEMA_signal_3840), .Z1_t (new_AGEMA_signal_3841), .Z1_f (new_AGEMA_signal_3842) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_27_U1_XOR1_U1 ( .A0_t (Feedback[27]), .A0_f (new_AGEMA_signal_2721), .A1_t (new_AGEMA_signal_2722), .A1_f (new_AGEMA_signal_2723), .B0_t (Input_s0_t[27]), .B0_f (Input_s0_f[27]), .B1_t (Input_s1_t[27]), .B1_f (Input_s1_f[27]), .Z0_t (InputMUX_MUXInst_27_U1_X), .Z0_f (new_AGEMA_signal_3112), .Z1_t (new_AGEMA_signal_3113), .Z1_f (new_AGEMA_signal_3114) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_27_U1_X), .B0_f (new_AGEMA_signal_3112), .B1_t (new_AGEMA_signal_3113), .B1_f (new_AGEMA_signal_3114), .Z0_t (InputMUX_MUXInst_27_U1_Y), .Z0_f (new_AGEMA_signal_3443), .Z1_t (new_AGEMA_signal_3444), .Z1_f (new_AGEMA_signal_3445) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_27_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_27_U1_Y), .A0_f (new_AGEMA_signal_3443), .A1_t (new_AGEMA_signal_3444), .A1_f (new_AGEMA_signal_3445), .B0_t (Feedback[27]), .B0_f (new_AGEMA_signal_2721), .B1_t (new_AGEMA_signal_2722), .B1_f (new_AGEMA_signal_2723), .Z0_t (MCOutput[27]), .Z0_f (new_AGEMA_signal_3690), .Z1_t (new_AGEMA_signal_3691), .Z1_f (new_AGEMA_signal_3692) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_28_U1_XOR1_U1 ( .A0_t (Feedback[28]), .A0_f (new_AGEMA_signal_3265), .A1_t (new_AGEMA_signal_3266), .A1_f (new_AGEMA_signal_3267), .B0_t (Input_s0_t[28]), .B0_f (Input_s0_f[28]), .B1_t (Input_s1_t[28]), .B1_f (Input_s1_f[28]), .Z0_t (InputMUX_MUXInst_28_U1_X), .Z0_f (new_AGEMA_signal_3449), .Z1_t (new_AGEMA_signal_3450), .Z1_f (new_AGEMA_signal_3451) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_28_U1_X), .B0_f (new_AGEMA_signal_3449), .B1_t (new_AGEMA_signal_3450), .B1_f (new_AGEMA_signal_3451), .Z0_t (InputMUX_MUXInst_28_U1_Y), .Z0_f (new_AGEMA_signal_3693), .Z1_t (new_AGEMA_signal_3694), .Z1_f (new_AGEMA_signal_3695) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_28_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_28_U1_Y), .A0_f (new_AGEMA_signal_3693), .A1_t (new_AGEMA_signal_3694), .A1_f (new_AGEMA_signal_3695), .B0_t (Feedback[28]), .B0_f (new_AGEMA_signal_3265), .B1_t (new_AGEMA_signal_3266), .B1_f (new_AGEMA_signal_3267), .Z0_t (MCOutput[28]), .Z0_f (new_AGEMA_signal_3843), .Z1_t (new_AGEMA_signal_3844), .Z1_f (new_AGEMA_signal_3845) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_29_U1_XOR1_U1 ( .A0_t (Feedback[29]), .A0_f (new_AGEMA_signal_2730), .A1_t (new_AGEMA_signal_2731), .A1_f (new_AGEMA_signal_2732), .B0_t (Input_s0_t[29]), .B0_f (Input_s0_f[29]), .B1_t (Input_s1_t[29]), .B1_f (Input_s1_f[29]), .Z0_t (InputMUX_MUXInst_29_U1_X), .Z0_f (new_AGEMA_signal_3118), .Z1_t (new_AGEMA_signal_3119), .Z1_f (new_AGEMA_signal_3120) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_29_U1_X), .B0_f (new_AGEMA_signal_3118), .B1_t (new_AGEMA_signal_3119), .B1_f (new_AGEMA_signal_3120), .Z0_t (InputMUX_MUXInst_29_U1_Y), .Z0_f (new_AGEMA_signal_3452), .Z1_t (new_AGEMA_signal_3453), .Z1_f (new_AGEMA_signal_3454) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_29_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_29_U1_Y), .A0_f (new_AGEMA_signal_3452), .A1_t (new_AGEMA_signal_3453), .A1_f (new_AGEMA_signal_3454), .B0_t (Feedback[29]), .B0_f (new_AGEMA_signal_2730), .B1_t (new_AGEMA_signal_2731), .B1_f (new_AGEMA_signal_2732), .Z0_t (MCOutput[29]), .Z0_f (new_AGEMA_signal_3696), .Z1_t (new_AGEMA_signal_3697), .Z1_f (new_AGEMA_signal_3698) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_30_U1_XOR1_U1 ( .A0_t (Feedback[30]), .A0_f (new_AGEMA_signal_3268), .A1_t (new_AGEMA_signal_3269), .A1_f (new_AGEMA_signal_3270), .B0_t (Input_s0_t[30]), .B0_f (Input_s0_f[30]), .B1_t (Input_s1_t[30]), .B1_f (Input_s1_f[30]), .Z0_t (InputMUX_MUXInst_30_U1_X), .Z0_f (new_AGEMA_signal_3458), .Z1_t (new_AGEMA_signal_3459), .Z1_f (new_AGEMA_signal_3460) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_30_U1_X), .B0_f (new_AGEMA_signal_3458), .B1_t (new_AGEMA_signal_3459), .B1_f (new_AGEMA_signal_3460), .Z0_t (InputMUX_MUXInst_30_U1_Y), .Z0_f (new_AGEMA_signal_3699), .Z1_t (new_AGEMA_signal_3700), .Z1_f (new_AGEMA_signal_3701) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_30_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_30_U1_Y), .A0_f (new_AGEMA_signal_3699), .A1_t (new_AGEMA_signal_3700), .A1_f (new_AGEMA_signal_3701), .B0_t (Feedback[30]), .B0_f (new_AGEMA_signal_3268), .B1_t (new_AGEMA_signal_3269), .B1_f (new_AGEMA_signal_3270), .Z0_t (MCOutput[30]), .Z0_f (new_AGEMA_signal_3846), .Z1_t (new_AGEMA_signal_3847), .Z1_f (new_AGEMA_signal_3848) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_31_U1_XOR1_U1 ( .A0_t (Feedback[31]), .A0_f (new_AGEMA_signal_2733), .A1_t (new_AGEMA_signal_2734), .A1_f (new_AGEMA_signal_2735), .B0_t (Input_s0_t[31]), .B0_f (Input_s0_f[31]), .B1_t (Input_s1_t[31]), .B1_f (Input_s1_f[31]), .Z0_t (InputMUX_MUXInst_31_U1_X), .Z0_f (new_AGEMA_signal_3124), .Z1_t (new_AGEMA_signal_3125), .Z1_f (new_AGEMA_signal_3126) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_31_U1_X), .B0_f (new_AGEMA_signal_3124), .B1_t (new_AGEMA_signal_3125), .B1_f (new_AGEMA_signal_3126), .Z0_t (InputMUX_MUXInst_31_U1_Y), .Z0_f (new_AGEMA_signal_3461), .Z1_t (new_AGEMA_signal_3462), .Z1_f (new_AGEMA_signal_3463) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_31_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_31_U1_Y), .A0_f (new_AGEMA_signal_3461), .A1_t (new_AGEMA_signal_3462), .A1_f (new_AGEMA_signal_3463), .B0_t (Feedback[31]), .B0_f (new_AGEMA_signal_2733), .B1_t (new_AGEMA_signal_2734), .B1_f (new_AGEMA_signal_2735), .Z0_t (MCOutput[31]), .Z0_f (new_AGEMA_signal_3702), .Z1_t (new_AGEMA_signal_3703), .Z1_f (new_AGEMA_signal_3704) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_32_U1_XOR1_U1 ( .A0_t (Feedback[32]), .A0_f (new_AGEMA_signal_3274), .A1_t (new_AGEMA_signal_3275), .A1_f (new_AGEMA_signal_3276), .B0_t (Input_s0_t[32]), .B0_f (Input_s0_f[32]), .B1_t (Input_s1_t[32]), .B1_f (Input_s1_f[32]), .Z0_t (InputMUX_MUXInst_32_U1_X), .Z0_f (new_AGEMA_signal_3467), .Z1_t (new_AGEMA_signal_3468), .Z1_f (new_AGEMA_signal_3469) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_32_U1_X), .B0_f (new_AGEMA_signal_3467), .B1_t (new_AGEMA_signal_3468), .B1_f (new_AGEMA_signal_3469), .Z0_t (InputMUX_MUXInst_32_U1_Y), .Z0_f (new_AGEMA_signal_3705), .Z1_t (new_AGEMA_signal_3706), .Z1_f (new_AGEMA_signal_3707) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_32_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_32_U1_Y), .A0_f (new_AGEMA_signal_3705), .A1_t (new_AGEMA_signal_3706), .A1_f (new_AGEMA_signal_3707), .B0_t (Feedback[32]), .B0_f (new_AGEMA_signal_3274), .B1_t (new_AGEMA_signal_3275), .B1_f (new_AGEMA_signal_3276), .Z0_t (MCInput[32]), .Z0_f (new_AGEMA_signal_3849), .Z1_t (new_AGEMA_signal_3850), .Z1_f (new_AGEMA_signal_3851) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_33_U1_XOR1_U1 ( .A0_t (Feedback[33]), .A0_f (new_AGEMA_signal_2742), .A1_t (new_AGEMA_signal_2743), .A1_f (new_AGEMA_signal_2744), .B0_t (Input_s0_t[33]), .B0_f (Input_s0_f[33]), .B1_t (Input_s1_t[33]), .B1_f (Input_s1_f[33]), .Z0_t (InputMUX_MUXInst_33_U1_X), .Z0_f (new_AGEMA_signal_3130), .Z1_t (new_AGEMA_signal_3131), .Z1_f (new_AGEMA_signal_3132) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_33_U1_X), .B0_f (new_AGEMA_signal_3130), .B1_t (new_AGEMA_signal_3131), .B1_f (new_AGEMA_signal_3132), .Z0_t (InputMUX_MUXInst_33_U1_Y), .Z0_f (new_AGEMA_signal_3470), .Z1_t (new_AGEMA_signal_3471), .Z1_f (new_AGEMA_signal_3472) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_33_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_33_U1_Y), .A0_f (new_AGEMA_signal_3470), .A1_t (new_AGEMA_signal_3471), .A1_f (new_AGEMA_signal_3472), .B0_t (Feedback[33]), .B0_f (new_AGEMA_signal_2742), .B1_t (new_AGEMA_signal_2743), .B1_f (new_AGEMA_signal_2744), .Z0_t (MCInput[33]), .Z0_f (new_AGEMA_signal_3708), .Z1_t (new_AGEMA_signal_3709), .Z1_f (new_AGEMA_signal_3710) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_34_U1_XOR1_U1 ( .A0_t (Feedback[34]), .A0_f (new_AGEMA_signal_3271), .A1_t (new_AGEMA_signal_3272), .A1_f (new_AGEMA_signal_3273), .B0_t (Input_s0_t[34]), .B0_f (Input_s0_f[34]), .B1_t (Input_s1_t[34]), .B1_f (Input_s1_f[34]), .Z0_t (InputMUX_MUXInst_34_U1_X), .Z0_f (new_AGEMA_signal_3476), .Z1_t (new_AGEMA_signal_3477), .Z1_f (new_AGEMA_signal_3478) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_34_U1_X), .B0_f (new_AGEMA_signal_3476), .B1_t (new_AGEMA_signal_3477), .B1_f (new_AGEMA_signal_3478), .Z0_t (InputMUX_MUXInst_34_U1_Y), .Z0_f (new_AGEMA_signal_3711), .Z1_t (new_AGEMA_signal_3712), .Z1_f (new_AGEMA_signal_3713) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_34_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_34_U1_Y), .A0_f (new_AGEMA_signal_3711), .A1_t (new_AGEMA_signal_3712), .A1_f (new_AGEMA_signal_3713), .B0_t (Feedback[34]), .B0_f (new_AGEMA_signal_3271), .B1_t (new_AGEMA_signal_3272), .B1_f (new_AGEMA_signal_3273), .Z0_t (MCInput[34]), .Z0_f (new_AGEMA_signal_3852), .Z1_t (new_AGEMA_signal_3853), .Z1_f (new_AGEMA_signal_3854) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_35_U1_XOR1_U1 ( .A0_t (Feedback[35]), .A0_f (new_AGEMA_signal_2745), .A1_t (new_AGEMA_signal_2746), .A1_f (new_AGEMA_signal_2747), .B0_t (Input_s0_t[35]), .B0_f (Input_s0_f[35]), .B1_t (Input_s1_t[35]), .B1_f (Input_s1_f[35]), .Z0_t (InputMUX_MUXInst_35_U1_X), .Z0_f (new_AGEMA_signal_3136), .Z1_t (new_AGEMA_signal_3137), .Z1_f (new_AGEMA_signal_3138) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_35_U1_X), .B0_f (new_AGEMA_signal_3136), .B1_t (new_AGEMA_signal_3137), .B1_f (new_AGEMA_signal_3138), .Z0_t (InputMUX_MUXInst_35_U1_Y), .Z0_f (new_AGEMA_signal_3479), .Z1_t (new_AGEMA_signal_3480), .Z1_f (new_AGEMA_signal_3481) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_35_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_35_U1_Y), .A0_f (new_AGEMA_signal_3479), .A1_t (new_AGEMA_signal_3480), .A1_f (new_AGEMA_signal_3481), .B0_t (Feedback[35]), .B0_f (new_AGEMA_signal_2745), .B1_t (new_AGEMA_signal_2746), .B1_f (new_AGEMA_signal_2747), .Z0_t (MCInput[35]), .Z0_f (new_AGEMA_signal_3714), .Z1_t (new_AGEMA_signal_3715), .Z1_f (new_AGEMA_signal_3716) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_36_U1_XOR1_U1 ( .A0_t (Feedback[36]), .A0_f (new_AGEMA_signal_3280), .A1_t (new_AGEMA_signal_3281), .A1_f (new_AGEMA_signal_3282), .B0_t (Input_s0_t[36]), .B0_f (Input_s0_f[36]), .B1_t (Input_s1_t[36]), .B1_f (Input_s1_f[36]), .Z0_t (InputMUX_MUXInst_36_U1_X), .Z0_f (new_AGEMA_signal_3485), .Z1_t (new_AGEMA_signal_3486), .Z1_f (new_AGEMA_signal_3487) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_36_U1_X), .B0_f (new_AGEMA_signal_3485), .B1_t (new_AGEMA_signal_3486), .B1_f (new_AGEMA_signal_3487), .Z0_t (InputMUX_MUXInst_36_U1_Y), .Z0_f (new_AGEMA_signal_3717), .Z1_t (new_AGEMA_signal_3718), .Z1_f (new_AGEMA_signal_3719) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_36_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_36_U1_Y), .A0_f (new_AGEMA_signal_3717), .A1_t (new_AGEMA_signal_3718), .A1_f (new_AGEMA_signal_3719), .B0_t (Feedback[36]), .B0_f (new_AGEMA_signal_3280), .B1_t (new_AGEMA_signal_3281), .B1_f (new_AGEMA_signal_3282), .Z0_t (MCInput[36]), .Z0_f (new_AGEMA_signal_3855), .Z1_t (new_AGEMA_signal_3856), .Z1_f (new_AGEMA_signal_3857) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_37_U1_XOR1_U1 ( .A0_t (Feedback[37]), .A0_f (new_AGEMA_signal_2754), .A1_t (new_AGEMA_signal_2755), .A1_f (new_AGEMA_signal_2756), .B0_t (Input_s0_t[37]), .B0_f (Input_s0_f[37]), .B1_t (Input_s1_t[37]), .B1_f (Input_s1_f[37]), .Z0_t (InputMUX_MUXInst_37_U1_X), .Z0_f (new_AGEMA_signal_3142), .Z1_t (new_AGEMA_signal_3143), .Z1_f (new_AGEMA_signal_3144) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_37_U1_X), .B0_f (new_AGEMA_signal_3142), .B1_t (new_AGEMA_signal_3143), .B1_f (new_AGEMA_signal_3144), .Z0_t (InputMUX_MUXInst_37_U1_Y), .Z0_f (new_AGEMA_signal_3488), .Z1_t (new_AGEMA_signal_3489), .Z1_f (new_AGEMA_signal_3490) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_37_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_37_U1_Y), .A0_f (new_AGEMA_signal_3488), .A1_t (new_AGEMA_signal_3489), .A1_f (new_AGEMA_signal_3490), .B0_t (Feedback[37]), .B0_f (new_AGEMA_signal_2754), .B1_t (new_AGEMA_signal_2755), .B1_f (new_AGEMA_signal_2756), .Z0_t (MCInput[37]), .Z0_f (new_AGEMA_signal_3720), .Z1_t (new_AGEMA_signal_3721), .Z1_f (new_AGEMA_signal_3722) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_38_U1_XOR1_U1 ( .A0_t (Feedback[38]), .A0_f (new_AGEMA_signal_3277), .A1_t (new_AGEMA_signal_3278), .A1_f (new_AGEMA_signal_3279), .B0_t (Input_s0_t[38]), .B0_f (Input_s0_f[38]), .B1_t (Input_s1_t[38]), .B1_f (Input_s1_f[38]), .Z0_t (InputMUX_MUXInst_38_U1_X), .Z0_f (new_AGEMA_signal_3494), .Z1_t (new_AGEMA_signal_3495), .Z1_f (new_AGEMA_signal_3496) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_38_U1_X), .B0_f (new_AGEMA_signal_3494), .B1_t (new_AGEMA_signal_3495), .B1_f (new_AGEMA_signal_3496), .Z0_t (InputMUX_MUXInst_38_U1_Y), .Z0_f (new_AGEMA_signal_3723), .Z1_t (new_AGEMA_signal_3724), .Z1_f (new_AGEMA_signal_3725) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_38_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_38_U1_Y), .A0_f (new_AGEMA_signal_3723), .A1_t (new_AGEMA_signal_3724), .A1_f (new_AGEMA_signal_3725), .B0_t (Feedback[38]), .B0_f (new_AGEMA_signal_3277), .B1_t (new_AGEMA_signal_3278), .B1_f (new_AGEMA_signal_3279), .Z0_t (MCInput[38]), .Z0_f (new_AGEMA_signal_3858), .Z1_t (new_AGEMA_signal_3859), .Z1_f (new_AGEMA_signal_3860) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_39_U1_XOR1_U1 ( .A0_t (Feedback[39]), .A0_f (new_AGEMA_signal_2757), .A1_t (new_AGEMA_signal_2758), .A1_f (new_AGEMA_signal_2759), .B0_t (Input_s0_t[39]), .B0_f (Input_s0_f[39]), .B1_t (Input_s1_t[39]), .B1_f (Input_s1_f[39]), .Z0_t (InputMUX_MUXInst_39_U1_X), .Z0_f (new_AGEMA_signal_3148), .Z1_t (new_AGEMA_signal_3149), .Z1_f (new_AGEMA_signal_3150) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_39_U1_X), .B0_f (new_AGEMA_signal_3148), .B1_t (new_AGEMA_signal_3149), .B1_f (new_AGEMA_signal_3150), .Z0_t (InputMUX_MUXInst_39_U1_Y), .Z0_f (new_AGEMA_signal_3497), .Z1_t (new_AGEMA_signal_3498), .Z1_f (new_AGEMA_signal_3499) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_39_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_39_U1_Y), .A0_f (new_AGEMA_signal_3497), .A1_t (new_AGEMA_signal_3498), .A1_f (new_AGEMA_signal_3499), .B0_t (Feedback[39]), .B0_f (new_AGEMA_signal_2757), .B1_t (new_AGEMA_signal_2758), .B1_f (new_AGEMA_signal_2759), .Z0_t (MCInput[39]), .Z0_f (new_AGEMA_signal_3726), .Z1_t (new_AGEMA_signal_3727), .Z1_f (new_AGEMA_signal_3728) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_40_U1_XOR1_U1 ( .A0_t (Feedback[40]), .A0_f (new_AGEMA_signal_3286), .A1_t (new_AGEMA_signal_3287), .A1_f (new_AGEMA_signal_3288), .B0_t (Input_s0_t[40]), .B0_f (Input_s0_f[40]), .B1_t (Input_s1_t[40]), .B1_f (Input_s1_f[40]), .Z0_t (InputMUX_MUXInst_40_U1_X), .Z0_f (new_AGEMA_signal_3503), .Z1_t (new_AGEMA_signal_3504), .Z1_f (new_AGEMA_signal_3505) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_40_U1_X), .B0_f (new_AGEMA_signal_3503), .B1_t (new_AGEMA_signal_3504), .B1_f (new_AGEMA_signal_3505), .Z0_t (InputMUX_MUXInst_40_U1_Y), .Z0_f (new_AGEMA_signal_3729), .Z1_t (new_AGEMA_signal_3730), .Z1_f (new_AGEMA_signal_3731) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_40_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_40_U1_Y), .A0_f (new_AGEMA_signal_3729), .A1_t (new_AGEMA_signal_3730), .A1_f (new_AGEMA_signal_3731), .B0_t (Feedback[40]), .B0_f (new_AGEMA_signal_3286), .B1_t (new_AGEMA_signal_3287), .B1_f (new_AGEMA_signal_3288), .Z0_t (MCInput[40]), .Z0_f (new_AGEMA_signal_3861), .Z1_t (new_AGEMA_signal_3862), .Z1_f (new_AGEMA_signal_3863) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_41_U1_XOR1_U1 ( .A0_t (Feedback[41]), .A0_f (new_AGEMA_signal_2766), .A1_t (new_AGEMA_signal_2767), .A1_f (new_AGEMA_signal_2768), .B0_t (Input_s0_t[41]), .B0_f (Input_s0_f[41]), .B1_t (Input_s1_t[41]), .B1_f (Input_s1_f[41]), .Z0_t (InputMUX_MUXInst_41_U1_X), .Z0_f (new_AGEMA_signal_3154), .Z1_t (new_AGEMA_signal_3155), .Z1_f (new_AGEMA_signal_3156) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_41_U1_X), .B0_f (new_AGEMA_signal_3154), .B1_t (new_AGEMA_signal_3155), .B1_f (new_AGEMA_signal_3156), .Z0_t (InputMUX_MUXInst_41_U1_Y), .Z0_f (new_AGEMA_signal_3506), .Z1_t (new_AGEMA_signal_3507), .Z1_f (new_AGEMA_signal_3508) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_41_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_41_U1_Y), .A0_f (new_AGEMA_signal_3506), .A1_t (new_AGEMA_signal_3507), .A1_f (new_AGEMA_signal_3508), .B0_t (Feedback[41]), .B0_f (new_AGEMA_signal_2766), .B1_t (new_AGEMA_signal_2767), .B1_f (new_AGEMA_signal_2768), .Z0_t (MCInput[41]), .Z0_f (new_AGEMA_signal_3732), .Z1_t (new_AGEMA_signal_3733), .Z1_f (new_AGEMA_signal_3734) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_42_U1_XOR1_U1 ( .A0_t (Feedback[42]), .A0_f (new_AGEMA_signal_3283), .A1_t (new_AGEMA_signal_3284), .A1_f (new_AGEMA_signal_3285), .B0_t (Input_s0_t[42]), .B0_f (Input_s0_f[42]), .B1_t (Input_s1_t[42]), .B1_f (Input_s1_f[42]), .Z0_t (InputMUX_MUXInst_42_U1_X), .Z0_f (new_AGEMA_signal_3512), .Z1_t (new_AGEMA_signal_3513), .Z1_f (new_AGEMA_signal_3514) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_42_U1_X), .B0_f (new_AGEMA_signal_3512), .B1_t (new_AGEMA_signal_3513), .B1_f (new_AGEMA_signal_3514), .Z0_t (InputMUX_MUXInst_42_U1_Y), .Z0_f (new_AGEMA_signal_3735), .Z1_t (new_AGEMA_signal_3736), .Z1_f (new_AGEMA_signal_3737) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_42_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_42_U1_Y), .A0_f (new_AGEMA_signal_3735), .A1_t (new_AGEMA_signal_3736), .A1_f (new_AGEMA_signal_3737), .B0_t (Feedback[42]), .B0_f (new_AGEMA_signal_3283), .B1_t (new_AGEMA_signal_3284), .B1_f (new_AGEMA_signal_3285), .Z0_t (MCInput[42]), .Z0_f (new_AGEMA_signal_3864), .Z1_t (new_AGEMA_signal_3865), .Z1_f (new_AGEMA_signal_3866) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_43_U1_XOR1_U1 ( .A0_t (Feedback[43]), .A0_f (new_AGEMA_signal_2769), .A1_t (new_AGEMA_signal_2770), .A1_f (new_AGEMA_signal_2771), .B0_t (Input_s0_t[43]), .B0_f (Input_s0_f[43]), .B1_t (Input_s1_t[43]), .B1_f (Input_s1_f[43]), .Z0_t (InputMUX_MUXInst_43_U1_X), .Z0_f (new_AGEMA_signal_3160), .Z1_t (new_AGEMA_signal_3161), .Z1_f (new_AGEMA_signal_3162) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_43_U1_X), .B0_f (new_AGEMA_signal_3160), .B1_t (new_AGEMA_signal_3161), .B1_f (new_AGEMA_signal_3162), .Z0_t (InputMUX_MUXInst_43_U1_Y), .Z0_f (new_AGEMA_signal_3515), .Z1_t (new_AGEMA_signal_3516), .Z1_f (new_AGEMA_signal_3517) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_43_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_43_U1_Y), .A0_f (new_AGEMA_signal_3515), .A1_t (new_AGEMA_signal_3516), .A1_f (new_AGEMA_signal_3517), .B0_t (Feedback[43]), .B0_f (new_AGEMA_signal_2769), .B1_t (new_AGEMA_signal_2770), .B1_f (new_AGEMA_signal_2771), .Z0_t (MCInput[43]), .Z0_f (new_AGEMA_signal_3738), .Z1_t (new_AGEMA_signal_3739), .Z1_f (new_AGEMA_signal_3740) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_44_U1_XOR1_U1 ( .A0_t (Feedback[44]), .A0_f (new_AGEMA_signal_3292), .A1_t (new_AGEMA_signal_3293), .A1_f (new_AGEMA_signal_3294), .B0_t (Input_s0_t[44]), .B0_f (Input_s0_f[44]), .B1_t (Input_s1_t[44]), .B1_f (Input_s1_f[44]), .Z0_t (InputMUX_MUXInst_44_U1_X), .Z0_f (new_AGEMA_signal_3521), .Z1_t (new_AGEMA_signal_3522), .Z1_f (new_AGEMA_signal_3523) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_44_U1_X), .B0_f (new_AGEMA_signal_3521), .B1_t (new_AGEMA_signal_3522), .B1_f (new_AGEMA_signal_3523), .Z0_t (InputMUX_MUXInst_44_U1_Y), .Z0_f (new_AGEMA_signal_3741), .Z1_t (new_AGEMA_signal_3742), .Z1_f (new_AGEMA_signal_3743) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_44_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_44_U1_Y), .A0_f (new_AGEMA_signal_3741), .A1_t (new_AGEMA_signal_3742), .A1_f (new_AGEMA_signal_3743), .B0_t (Feedback[44]), .B0_f (new_AGEMA_signal_3292), .B1_t (new_AGEMA_signal_3293), .B1_f (new_AGEMA_signal_3294), .Z0_t (MCInput[44]), .Z0_f (new_AGEMA_signal_3867), .Z1_t (new_AGEMA_signal_3868), .Z1_f (new_AGEMA_signal_3869) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_45_U1_XOR1_U1 ( .A0_t (Feedback[45]), .A0_f (new_AGEMA_signal_2778), .A1_t (new_AGEMA_signal_2779), .A1_f (new_AGEMA_signal_2780), .B0_t (Input_s0_t[45]), .B0_f (Input_s0_f[45]), .B1_t (Input_s1_t[45]), .B1_f (Input_s1_f[45]), .Z0_t (InputMUX_MUXInst_45_U1_X), .Z0_f (new_AGEMA_signal_3166), .Z1_t (new_AGEMA_signal_3167), .Z1_f (new_AGEMA_signal_3168) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_45_U1_X), .B0_f (new_AGEMA_signal_3166), .B1_t (new_AGEMA_signal_3167), .B1_f (new_AGEMA_signal_3168), .Z0_t (InputMUX_MUXInst_45_U1_Y), .Z0_f (new_AGEMA_signal_3524), .Z1_t (new_AGEMA_signal_3525), .Z1_f (new_AGEMA_signal_3526) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_45_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_45_U1_Y), .A0_f (new_AGEMA_signal_3524), .A1_t (new_AGEMA_signal_3525), .A1_f (new_AGEMA_signal_3526), .B0_t (Feedback[45]), .B0_f (new_AGEMA_signal_2778), .B1_t (new_AGEMA_signal_2779), .B1_f (new_AGEMA_signal_2780), .Z0_t (MCInput[45]), .Z0_f (new_AGEMA_signal_3744), .Z1_t (new_AGEMA_signal_3745), .Z1_f (new_AGEMA_signal_3746) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_46_U1_XOR1_U1 ( .A0_t (Feedback[46]), .A0_f (new_AGEMA_signal_3289), .A1_t (new_AGEMA_signal_3290), .A1_f (new_AGEMA_signal_3291), .B0_t (Input_s0_t[46]), .B0_f (Input_s0_f[46]), .B1_t (Input_s1_t[46]), .B1_f (Input_s1_f[46]), .Z0_t (InputMUX_MUXInst_46_U1_X), .Z0_f (new_AGEMA_signal_3530), .Z1_t (new_AGEMA_signal_3531), .Z1_f (new_AGEMA_signal_3532) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_46_U1_X), .B0_f (new_AGEMA_signal_3530), .B1_t (new_AGEMA_signal_3531), .B1_f (new_AGEMA_signal_3532), .Z0_t (InputMUX_MUXInst_46_U1_Y), .Z0_f (new_AGEMA_signal_3747), .Z1_t (new_AGEMA_signal_3748), .Z1_f (new_AGEMA_signal_3749) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_46_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_46_U1_Y), .A0_f (new_AGEMA_signal_3747), .A1_t (new_AGEMA_signal_3748), .A1_f (new_AGEMA_signal_3749), .B0_t (Feedback[46]), .B0_f (new_AGEMA_signal_3289), .B1_t (new_AGEMA_signal_3290), .B1_f (new_AGEMA_signal_3291), .Z0_t (MCInput[46]), .Z0_f (new_AGEMA_signal_3870), .Z1_t (new_AGEMA_signal_3871), .Z1_f (new_AGEMA_signal_3872) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_47_U1_XOR1_U1 ( .A0_t (Feedback[47]), .A0_f (new_AGEMA_signal_2781), .A1_t (new_AGEMA_signal_2782), .A1_f (new_AGEMA_signal_2783), .B0_t (Input_s0_t[47]), .B0_f (Input_s0_f[47]), .B1_t (Input_s1_t[47]), .B1_f (Input_s1_f[47]), .Z0_t (InputMUX_MUXInst_47_U1_X), .Z0_f (new_AGEMA_signal_3172), .Z1_t (new_AGEMA_signal_3173), .Z1_f (new_AGEMA_signal_3174) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_47_U1_X), .B0_f (new_AGEMA_signal_3172), .B1_t (new_AGEMA_signal_3173), .B1_f (new_AGEMA_signal_3174), .Z0_t (InputMUX_MUXInst_47_U1_Y), .Z0_f (new_AGEMA_signal_3533), .Z1_t (new_AGEMA_signal_3534), .Z1_f (new_AGEMA_signal_3535) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_47_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_47_U1_Y), .A0_f (new_AGEMA_signal_3533), .A1_t (new_AGEMA_signal_3534), .A1_f (new_AGEMA_signal_3535), .B0_t (Feedback[47]), .B0_f (new_AGEMA_signal_2781), .B1_t (new_AGEMA_signal_2782), .B1_f (new_AGEMA_signal_2783), .Z0_t (MCInput[47]), .Z0_f (new_AGEMA_signal_3750), .Z1_t (new_AGEMA_signal_3751), .Z1_f (new_AGEMA_signal_3752) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_48_U1_XOR1_U1 ( .A0_t (Feedback[48]), .A0_f (new_AGEMA_signal_3298), .A1_t (new_AGEMA_signal_3299), .A1_f (new_AGEMA_signal_3300), .B0_t (Input_s0_t[48]), .B0_f (Input_s0_f[48]), .B1_t (Input_s1_t[48]), .B1_f (Input_s1_f[48]), .Z0_t (InputMUX_MUXInst_48_U1_X), .Z0_f (new_AGEMA_signal_3539), .Z1_t (new_AGEMA_signal_3540), .Z1_f (new_AGEMA_signal_3541) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_48_U1_X), .B0_f (new_AGEMA_signal_3539), .B1_t (new_AGEMA_signal_3540), .B1_f (new_AGEMA_signal_3541), .Z0_t (InputMUX_MUXInst_48_U1_Y), .Z0_f (new_AGEMA_signal_3753), .Z1_t (new_AGEMA_signal_3754), .Z1_f (new_AGEMA_signal_3755) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_48_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_48_U1_Y), .A0_f (new_AGEMA_signal_3753), .A1_t (new_AGEMA_signal_3754), .A1_f (new_AGEMA_signal_3755), .B0_t (Feedback[48]), .B0_f (new_AGEMA_signal_3298), .B1_t (new_AGEMA_signal_3299), .B1_f (new_AGEMA_signal_3300), .Z0_t (MCInput[48]), .Z0_f (new_AGEMA_signal_3873), .Z1_t (new_AGEMA_signal_3874), .Z1_f (new_AGEMA_signal_3875) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_49_U1_XOR1_U1 ( .A0_t (Feedback[49]), .A0_f (new_AGEMA_signal_2790), .A1_t (new_AGEMA_signal_2791), .A1_f (new_AGEMA_signal_2792), .B0_t (Input_s0_t[49]), .B0_f (Input_s0_f[49]), .B1_t (Input_s1_t[49]), .B1_f (Input_s1_f[49]), .Z0_t (InputMUX_MUXInst_49_U1_X), .Z0_f (new_AGEMA_signal_3178), .Z1_t (new_AGEMA_signal_3179), .Z1_f (new_AGEMA_signal_3180) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_49_U1_X), .B0_f (new_AGEMA_signal_3178), .B1_t (new_AGEMA_signal_3179), .B1_f (new_AGEMA_signal_3180), .Z0_t (InputMUX_MUXInst_49_U1_Y), .Z0_f (new_AGEMA_signal_3542), .Z1_t (new_AGEMA_signal_3543), .Z1_f (new_AGEMA_signal_3544) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_49_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_49_U1_Y), .A0_f (new_AGEMA_signal_3542), .A1_t (new_AGEMA_signal_3543), .A1_f (new_AGEMA_signal_3544), .B0_t (Feedback[49]), .B0_f (new_AGEMA_signal_2790), .B1_t (new_AGEMA_signal_2791), .B1_f (new_AGEMA_signal_2792), .Z0_t (MCInput[49]), .Z0_f (new_AGEMA_signal_3756), .Z1_t (new_AGEMA_signal_3757), .Z1_f (new_AGEMA_signal_3758) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_50_U1_XOR1_U1 ( .A0_t (Feedback[50]), .A0_f (new_AGEMA_signal_3295), .A1_t (new_AGEMA_signal_3296), .A1_f (new_AGEMA_signal_3297), .B0_t (Input_s0_t[50]), .B0_f (Input_s0_f[50]), .B1_t (Input_s1_t[50]), .B1_f (Input_s1_f[50]), .Z0_t (InputMUX_MUXInst_50_U1_X), .Z0_f (new_AGEMA_signal_3548), .Z1_t (new_AGEMA_signal_3549), .Z1_f (new_AGEMA_signal_3550) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_50_U1_X), .B0_f (new_AGEMA_signal_3548), .B1_t (new_AGEMA_signal_3549), .B1_f (new_AGEMA_signal_3550), .Z0_t (InputMUX_MUXInst_50_U1_Y), .Z0_f (new_AGEMA_signal_3759), .Z1_t (new_AGEMA_signal_3760), .Z1_f (new_AGEMA_signal_3761) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_50_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_50_U1_Y), .A0_f (new_AGEMA_signal_3759), .A1_t (new_AGEMA_signal_3760), .A1_f (new_AGEMA_signal_3761), .B0_t (Feedback[50]), .B0_f (new_AGEMA_signal_3295), .B1_t (new_AGEMA_signal_3296), .B1_f (new_AGEMA_signal_3297), .Z0_t (MCInput[50]), .Z0_f (new_AGEMA_signal_3876), .Z1_t (new_AGEMA_signal_3877), .Z1_f (new_AGEMA_signal_3878) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_51_U1_XOR1_U1 ( .A0_t (Feedback[51]), .A0_f (new_AGEMA_signal_2793), .A1_t (new_AGEMA_signal_2794), .A1_f (new_AGEMA_signal_2795), .B0_t (Input_s0_t[51]), .B0_f (Input_s0_f[51]), .B1_t (Input_s1_t[51]), .B1_f (Input_s1_f[51]), .Z0_t (InputMUX_MUXInst_51_U1_X), .Z0_f (new_AGEMA_signal_3184), .Z1_t (new_AGEMA_signal_3185), .Z1_f (new_AGEMA_signal_3186) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_51_U1_X), .B0_f (new_AGEMA_signal_3184), .B1_t (new_AGEMA_signal_3185), .B1_f (new_AGEMA_signal_3186), .Z0_t (InputMUX_MUXInst_51_U1_Y), .Z0_f (new_AGEMA_signal_3551), .Z1_t (new_AGEMA_signal_3552), .Z1_f (new_AGEMA_signal_3553) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_51_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_51_U1_Y), .A0_f (new_AGEMA_signal_3551), .A1_t (new_AGEMA_signal_3552), .A1_f (new_AGEMA_signal_3553), .B0_t (Feedback[51]), .B0_f (new_AGEMA_signal_2793), .B1_t (new_AGEMA_signal_2794), .B1_f (new_AGEMA_signal_2795), .Z0_t (MCInput[51]), .Z0_f (new_AGEMA_signal_3762), .Z1_t (new_AGEMA_signal_3763), .Z1_f (new_AGEMA_signal_3764) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_52_U1_XOR1_U1 ( .A0_t (Feedback[52]), .A0_f (new_AGEMA_signal_3304), .A1_t (new_AGEMA_signal_3305), .A1_f (new_AGEMA_signal_3306), .B0_t (Input_s0_t[52]), .B0_f (Input_s0_f[52]), .B1_t (Input_s1_t[52]), .B1_f (Input_s1_f[52]), .Z0_t (InputMUX_MUXInst_52_U1_X), .Z0_f (new_AGEMA_signal_3557), .Z1_t (new_AGEMA_signal_3558), .Z1_f (new_AGEMA_signal_3559) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_52_U1_X), .B0_f (new_AGEMA_signal_3557), .B1_t (new_AGEMA_signal_3558), .B1_f (new_AGEMA_signal_3559), .Z0_t (InputMUX_MUXInst_52_U1_Y), .Z0_f (new_AGEMA_signal_3765), .Z1_t (new_AGEMA_signal_3766), .Z1_f (new_AGEMA_signal_3767) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_52_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_52_U1_Y), .A0_f (new_AGEMA_signal_3765), .A1_t (new_AGEMA_signal_3766), .A1_f (new_AGEMA_signal_3767), .B0_t (Feedback[52]), .B0_f (new_AGEMA_signal_3304), .B1_t (new_AGEMA_signal_3305), .B1_f (new_AGEMA_signal_3306), .Z0_t (MCInput[52]), .Z0_f (new_AGEMA_signal_3879), .Z1_t (new_AGEMA_signal_3880), .Z1_f (new_AGEMA_signal_3881) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_53_U1_XOR1_U1 ( .A0_t (Feedback[53]), .A0_f (new_AGEMA_signal_2802), .A1_t (new_AGEMA_signal_2803), .A1_f (new_AGEMA_signal_2804), .B0_t (Input_s0_t[53]), .B0_f (Input_s0_f[53]), .B1_t (Input_s1_t[53]), .B1_f (Input_s1_f[53]), .Z0_t (InputMUX_MUXInst_53_U1_X), .Z0_f (new_AGEMA_signal_3190), .Z1_t (new_AGEMA_signal_3191), .Z1_f (new_AGEMA_signal_3192) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_53_U1_X), .B0_f (new_AGEMA_signal_3190), .B1_t (new_AGEMA_signal_3191), .B1_f (new_AGEMA_signal_3192), .Z0_t (InputMUX_MUXInst_53_U1_Y), .Z0_f (new_AGEMA_signal_3560), .Z1_t (new_AGEMA_signal_3561), .Z1_f (new_AGEMA_signal_3562) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_53_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_53_U1_Y), .A0_f (new_AGEMA_signal_3560), .A1_t (new_AGEMA_signal_3561), .A1_f (new_AGEMA_signal_3562), .B0_t (Feedback[53]), .B0_f (new_AGEMA_signal_2802), .B1_t (new_AGEMA_signal_2803), .B1_f (new_AGEMA_signal_2804), .Z0_t (MCInput[53]), .Z0_f (new_AGEMA_signal_3768), .Z1_t (new_AGEMA_signal_3769), .Z1_f (new_AGEMA_signal_3770) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_54_U1_XOR1_U1 ( .A0_t (Feedback[54]), .A0_f (new_AGEMA_signal_3301), .A1_t (new_AGEMA_signal_3302), .A1_f (new_AGEMA_signal_3303), .B0_t (Input_s0_t[54]), .B0_f (Input_s0_f[54]), .B1_t (Input_s1_t[54]), .B1_f (Input_s1_f[54]), .Z0_t (InputMUX_MUXInst_54_U1_X), .Z0_f (new_AGEMA_signal_3566), .Z1_t (new_AGEMA_signal_3567), .Z1_f (new_AGEMA_signal_3568) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_54_U1_X), .B0_f (new_AGEMA_signal_3566), .B1_t (new_AGEMA_signal_3567), .B1_f (new_AGEMA_signal_3568), .Z0_t (InputMUX_MUXInst_54_U1_Y), .Z0_f (new_AGEMA_signal_3771), .Z1_t (new_AGEMA_signal_3772), .Z1_f (new_AGEMA_signal_3773) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_54_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_54_U1_Y), .A0_f (new_AGEMA_signal_3771), .A1_t (new_AGEMA_signal_3772), .A1_f (new_AGEMA_signal_3773), .B0_t (Feedback[54]), .B0_f (new_AGEMA_signal_3301), .B1_t (new_AGEMA_signal_3302), .B1_f (new_AGEMA_signal_3303), .Z0_t (MCInput[54]), .Z0_f (new_AGEMA_signal_3882), .Z1_t (new_AGEMA_signal_3883), .Z1_f (new_AGEMA_signal_3884) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_55_U1_XOR1_U1 ( .A0_t (Feedback[55]), .A0_f (new_AGEMA_signal_2805), .A1_t (new_AGEMA_signal_2806), .A1_f (new_AGEMA_signal_2807), .B0_t (Input_s0_t[55]), .B0_f (Input_s0_f[55]), .B1_t (Input_s1_t[55]), .B1_f (Input_s1_f[55]), .Z0_t (InputMUX_MUXInst_55_U1_X), .Z0_f (new_AGEMA_signal_3196), .Z1_t (new_AGEMA_signal_3197), .Z1_f (new_AGEMA_signal_3198) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_55_U1_X), .B0_f (new_AGEMA_signal_3196), .B1_t (new_AGEMA_signal_3197), .B1_f (new_AGEMA_signal_3198), .Z0_t (InputMUX_MUXInst_55_U1_Y), .Z0_f (new_AGEMA_signal_3569), .Z1_t (new_AGEMA_signal_3570), .Z1_f (new_AGEMA_signal_3571) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_55_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_55_U1_Y), .A0_f (new_AGEMA_signal_3569), .A1_t (new_AGEMA_signal_3570), .A1_f (new_AGEMA_signal_3571), .B0_t (Feedback[55]), .B0_f (new_AGEMA_signal_2805), .B1_t (new_AGEMA_signal_2806), .B1_f (new_AGEMA_signal_2807), .Z0_t (MCInput[55]), .Z0_f (new_AGEMA_signal_3774), .Z1_t (new_AGEMA_signal_3775), .Z1_f (new_AGEMA_signal_3776) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_56_U1_XOR1_U1 ( .A0_t (Feedback[56]), .A0_f (new_AGEMA_signal_3310), .A1_t (new_AGEMA_signal_3311), .A1_f (new_AGEMA_signal_3312), .B0_t (Input_s0_t[56]), .B0_f (Input_s0_f[56]), .B1_t (Input_s1_t[56]), .B1_f (Input_s1_f[56]), .Z0_t (InputMUX_MUXInst_56_U1_X), .Z0_f (new_AGEMA_signal_3575), .Z1_t (new_AGEMA_signal_3576), .Z1_f (new_AGEMA_signal_3577) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_56_U1_X), .B0_f (new_AGEMA_signal_3575), .B1_t (new_AGEMA_signal_3576), .B1_f (new_AGEMA_signal_3577), .Z0_t (InputMUX_MUXInst_56_U1_Y), .Z0_f (new_AGEMA_signal_3777), .Z1_t (new_AGEMA_signal_3778), .Z1_f (new_AGEMA_signal_3779) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_56_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_56_U1_Y), .A0_f (new_AGEMA_signal_3777), .A1_t (new_AGEMA_signal_3778), .A1_f (new_AGEMA_signal_3779), .B0_t (Feedback[56]), .B0_f (new_AGEMA_signal_3310), .B1_t (new_AGEMA_signal_3311), .B1_f (new_AGEMA_signal_3312), .Z0_t (MCInput[56]), .Z0_f (new_AGEMA_signal_3885), .Z1_t (new_AGEMA_signal_3886), .Z1_f (new_AGEMA_signal_3887) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_57_U1_XOR1_U1 ( .A0_t (Feedback[57]), .A0_f (new_AGEMA_signal_2814), .A1_t (new_AGEMA_signal_2815), .A1_f (new_AGEMA_signal_2816), .B0_t (Input_s0_t[57]), .B0_f (Input_s0_f[57]), .B1_t (Input_s1_t[57]), .B1_f (Input_s1_f[57]), .Z0_t (InputMUX_MUXInst_57_U1_X), .Z0_f (new_AGEMA_signal_3202), .Z1_t (new_AGEMA_signal_3203), .Z1_f (new_AGEMA_signal_3204) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_57_U1_X), .B0_f (new_AGEMA_signal_3202), .B1_t (new_AGEMA_signal_3203), .B1_f (new_AGEMA_signal_3204), .Z0_t (InputMUX_MUXInst_57_U1_Y), .Z0_f (new_AGEMA_signal_3578), .Z1_t (new_AGEMA_signal_3579), .Z1_f (new_AGEMA_signal_3580) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_57_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_57_U1_Y), .A0_f (new_AGEMA_signal_3578), .A1_t (new_AGEMA_signal_3579), .A1_f (new_AGEMA_signal_3580), .B0_t (Feedback[57]), .B0_f (new_AGEMA_signal_2814), .B1_t (new_AGEMA_signal_2815), .B1_f (new_AGEMA_signal_2816), .Z0_t (MCInput[57]), .Z0_f (new_AGEMA_signal_3780), .Z1_t (new_AGEMA_signal_3781), .Z1_f (new_AGEMA_signal_3782) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_58_U1_XOR1_U1 ( .A0_t (Feedback[58]), .A0_f (new_AGEMA_signal_3307), .A1_t (new_AGEMA_signal_3308), .A1_f (new_AGEMA_signal_3309), .B0_t (Input_s0_t[58]), .B0_f (Input_s0_f[58]), .B1_t (Input_s1_t[58]), .B1_f (Input_s1_f[58]), .Z0_t (InputMUX_MUXInst_58_U1_X), .Z0_f (new_AGEMA_signal_3584), .Z1_t (new_AGEMA_signal_3585), .Z1_f (new_AGEMA_signal_3586) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_58_U1_X), .B0_f (new_AGEMA_signal_3584), .B1_t (new_AGEMA_signal_3585), .B1_f (new_AGEMA_signal_3586), .Z0_t (InputMUX_MUXInst_58_U1_Y), .Z0_f (new_AGEMA_signal_3783), .Z1_t (new_AGEMA_signal_3784), .Z1_f (new_AGEMA_signal_3785) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_58_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_58_U1_Y), .A0_f (new_AGEMA_signal_3783), .A1_t (new_AGEMA_signal_3784), .A1_f (new_AGEMA_signal_3785), .B0_t (Feedback[58]), .B0_f (new_AGEMA_signal_3307), .B1_t (new_AGEMA_signal_3308), .B1_f (new_AGEMA_signal_3309), .Z0_t (MCInput[58]), .Z0_f (new_AGEMA_signal_3888), .Z1_t (new_AGEMA_signal_3889), .Z1_f (new_AGEMA_signal_3890) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_59_U1_XOR1_U1 ( .A0_t (Feedback[59]), .A0_f (new_AGEMA_signal_2817), .A1_t (new_AGEMA_signal_2818), .A1_f (new_AGEMA_signal_2819), .B0_t (Input_s0_t[59]), .B0_f (Input_s0_f[59]), .B1_t (Input_s1_t[59]), .B1_f (Input_s1_f[59]), .Z0_t (InputMUX_MUXInst_59_U1_X), .Z0_f (new_AGEMA_signal_3208), .Z1_t (new_AGEMA_signal_3209), .Z1_f (new_AGEMA_signal_3210) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_59_U1_X), .B0_f (new_AGEMA_signal_3208), .B1_t (new_AGEMA_signal_3209), .B1_f (new_AGEMA_signal_3210), .Z0_t (InputMUX_MUXInst_59_U1_Y), .Z0_f (new_AGEMA_signal_3587), .Z1_t (new_AGEMA_signal_3588), .Z1_f (new_AGEMA_signal_3589) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_59_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_59_U1_Y), .A0_f (new_AGEMA_signal_3587), .A1_t (new_AGEMA_signal_3588), .A1_f (new_AGEMA_signal_3589), .B0_t (Feedback[59]), .B0_f (new_AGEMA_signal_2817), .B1_t (new_AGEMA_signal_2818), .B1_f (new_AGEMA_signal_2819), .Z0_t (MCInput[59]), .Z0_f (new_AGEMA_signal_3786), .Z1_t (new_AGEMA_signal_3787), .Z1_f (new_AGEMA_signal_3788) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_60_U1_XOR1_U1 ( .A0_t (Feedback[60]), .A0_f (new_AGEMA_signal_3316), .A1_t (new_AGEMA_signal_3317), .A1_f (new_AGEMA_signal_3318), .B0_t (Input_s0_t[60]), .B0_f (Input_s0_f[60]), .B1_t (Input_s1_t[60]), .B1_f (Input_s1_f[60]), .Z0_t (InputMUX_MUXInst_60_U1_X), .Z0_f (new_AGEMA_signal_3593), .Z1_t (new_AGEMA_signal_3594), .Z1_f (new_AGEMA_signal_3595) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_60_U1_X), .B0_f (new_AGEMA_signal_3593), .B1_t (new_AGEMA_signal_3594), .B1_f (new_AGEMA_signal_3595), .Z0_t (InputMUX_MUXInst_60_U1_Y), .Z0_f (new_AGEMA_signal_3789), .Z1_t (new_AGEMA_signal_3790), .Z1_f (new_AGEMA_signal_3791) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_60_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_60_U1_Y), .A0_f (new_AGEMA_signal_3789), .A1_t (new_AGEMA_signal_3790), .A1_f (new_AGEMA_signal_3791), .B0_t (Feedback[60]), .B0_f (new_AGEMA_signal_3316), .B1_t (new_AGEMA_signal_3317), .B1_f (new_AGEMA_signal_3318), .Z0_t (MCInput[60]), .Z0_f (new_AGEMA_signal_3891), .Z1_t (new_AGEMA_signal_3892), .Z1_f (new_AGEMA_signal_3893) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_61_U1_XOR1_U1 ( .A0_t (Feedback[61]), .A0_f (new_AGEMA_signal_2826), .A1_t (new_AGEMA_signal_2827), .A1_f (new_AGEMA_signal_2828), .B0_t (Input_s0_t[61]), .B0_f (Input_s0_f[61]), .B1_t (Input_s1_t[61]), .B1_f (Input_s1_f[61]), .Z0_t (InputMUX_MUXInst_61_U1_X), .Z0_f (new_AGEMA_signal_3214), .Z1_t (new_AGEMA_signal_3215), .Z1_f (new_AGEMA_signal_3216) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_61_U1_X), .B0_f (new_AGEMA_signal_3214), .B1_t (new_AGEMA_signal_3215), .B1_f (new_AGEMA_signal_3216), .Z0_t (InputMUX_MUXInst_61_U1_Y), .Z0_f (new_AGEMA_signal_3596), .Z1_t (new_AGEMA_signal_3597), .Z1_f (new_AGEMA_signal_3598) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_61_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_61_U1_Y), .A0_f (new_AGEMA_signal_3596), .A1_t (new_AGEMA_signal_3597), .A1_f (new_AGEMA_signal_3598), .B0_t (Feedback[61]), .B0_f (new_AGEMA_signal_2826), .B1_t (new_AGEMA_signal_2827), .B1_f (new_AGEMA_signal_2828), .Z0_t (MCInput[61]), .Z0_f (new_AGEMA_signal_3792), .Z1_t (new_AGEMA_signal_3793), .Z1_f (new_AGEMA_signal_3794) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_62_U1_XOR1_U1 ( .A0_t (Feedback[62]), .A0_f (new_AGEMA_signal_3313), .A1_t (new_AGEMA_signal_3314), .A1_f (new_AGEMA_signal_3315), .B0_t (Input_s0_t[62]), .B0_f (Input_s0_f[62]), .B1_t (Input_s1_t[62]), .B1_f (Input_s1_f[62]), .Z0_t (InputMUX_MUXInst_62_U1_X), .Z0_f (new_AGEMA_signal_3602), .Z1_t (new_AGEMA_signal_3603), .Z1_f (new_AGEMA_signal_3604) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_62_U1_X), .B0_f (new_AGEMA_signal_3602), .B1_t (new_AGEMA_signal_3603), .B1_f (new_AGEMA_signal_3604), .Z0_t (InputMUX_MUXInst_62_U1_Y), .Z0_f (new_AGEMA_signal_3795), .Z1_t (new_AGEMA_signal_3796), .Z1_f (new_AGEMA_signal_3797) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_62_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_62_U1_Y), .A0_f (new_AGEMA_signal_3795), .A1_t (new_AGEMA_signal_3796), .A1_f (new_AGEMA_signal_3797), .B0_t (Feedback[62]), .B0_f (new_AGEMA_signal_3313), .B1_t (new_AGEMA_signal_3314), .B1_f (new_AGEMA_signal_3315), .Z0_t (MCInput[62]), .Z0_f (new_AGEMA_signal_3894), .Z1_t (new_AGEMA_signal_3895), .Z1_f (new_AGEMA_signal_3896) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_63_U1_XOR1_U1 ( .A0_t (Feedback[63]), .A0_f (new_AGEMA_signal_2829), .A1_t (new_AGEMA_signal_2830), .A1_f (new_AGEMA_signal_2831), .B0_t (Input_s0_t[63]), .B0_f (Input_s0_f[63]), .B1_t (Input_s1_t[63]), .B1_f (Input_s1_f[63]), .Z0_t (InputMUX_MUXInst_63_U1_X), .Z0_f (new_AGEMA_signal_3220), .Z1_t (new_AGEMA_signal_3221), .Z1_f (new_AGEMA_signal_3222) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (rst_t), .A1_f (rst_f), .B0_t (InputMUX_MUXInst_63_U1_X), .B0_f (new_AGEMA_signal_3220), .B1_t (new_AGEMA_signal_3221), .B1_f (new_AGEMA_signal_3222), .Z0_t (InputMUX_MUXInst_63_U1_Y), .Z0_f (new_AGEMA_signal_3605), .Z1_t (new_AGEMA_signal_3606), .Z1_f (new_AGEMA_signal_3607) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) InputMUX_MUXInst_63_U1_XOR2_U1 ( .A0_t (InputMUX_MUXInst_63_U1_Y), .A0_f (new_AGEMA_signal_3605), .A1_t (new_AGEMA_signal_3606), .A1_f (new_AGEMA_signal_3607), .B0_t (Feedback[63]), .B0_f (new_AGEMA_signal_2829), .B1_t (new_AGEMA_signal_2830), .B1_f (new_AGEMA_signal_2831), .Z0_t (MCInput[63]), .Z0_f (new_AGEMA_signal_3798), .Z1_t (new_AGEMA_signal_3799), .Z1_f (new_AGEMA_signal_3800) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_0_U2 ( .A0_t (MCInst_XOR_r0_Inst_0_n1), .A0_f (new_AGEMA_signal_3945), .A1_t (new_AGEMA_signal_3946), .A1_f (new_AGEMA_signal_3947), .B0_t (MCOutput[0]), .B0_f (new_AGEMA_signal_3801), .B1_t (new_AGEMA_signal_3802), .B1_f (new_AGEMA_signal_3803), .Z0_t (MCOutput[48]), .Z0_f (new_AGEMA_signal_4026), .Z1_t (new_AGEMA_signal_4027), .Z1_f (new_AGEMA_signal_4028) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_0_U1 ( .A0_t (MCInput[48]), .A0_f (new_AGEMA_signal_3873), .A1_t (new_AGEMA_signal_3874), .A1_f (new_AGEMA_signal_3875), .B0_t (MCOutput[16]), .B0_f (new_AGEMA_signal_3825), .B1_t (new_AGEMA_signal_3826), .B1_f (new_AGEMA_signal_3827), .Z0_t (MCInst_XOR_r0_Inst_0_n1), .Z0_f (new_AGEMA_signal_3945), .Z1_t (new_AGEMA_signal_3946), .Z1_f (new_AGEMA_signal_3947) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_0_U1 ( .A0_t (MCInput[32]), .A0_f (new_AGEMA_signal_3849), .A1_t (new_AGEMA_signal_3850), .A1_f (new_AGEMA_signal_3851), .B0_t (MCOutput[0]), .B0_f (new_AGEMA_signal_3801), .B1_t (new_AGEMA_signal_3802), .B1_f (new_AGEMA_signal_3803), .Z0_t (MCOutput[32]), .Z0_f (new_AGEMA_signal_3948), .Z1_t (new_AGEMA_signal_3949), .Z1_f (new_AGEMA_signal_3950) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_1_U2 ( .A0_t (MCInst_XOR_r0_Inst_1_n1), .A0_f (new_AGEMA_signal_3897), .A1_t (new_AGEMA_signal_3898), .A1_f (new_AGEMA_signal_3899), .B0_t (MCOutput[1]), .B0_f (new_AGEMA_signal_3612), .B1_t (new_AGEMA_signal_3613), .B1_f (new_AGEMA_signal_3614), .Z0_t (MCOutput[49]), .Z0_f (new_AGEMA_signal_3951), .Z1_t (new_AGEMA_signal_3952), .Z1_f (new_AGEMA_signal_3953) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_1_U1 ( .A0_t (MCInput[49]), .A0_f (new_AGEMA_signal_3756), .A1_t (new_AGEMA_signal_3757), .A1_f (new_AGEMA_signal_3758), .B0_t (MCOutput[17]), .B0_f (new_AGEMA_signal_3660), .B1_t (new_AGEMA_signal_3661), .B1_f (new_AGEMA_signal_3662), .Z0_t (MCInst_XOR_r0_Inst_1_n1), .Z0_f (new_AGEMA_signal_3897), .Z1_t (new_AGEMA_signal_3898), .Z1_f (new_AGEMA_signal_3899) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_1_U1 ( .A0_t (MCInput[33]), .A0_f (new_AGEMA_signal_3708), .A1_t (new_AGEMA_signal_3709), .A1_f (new_AGEMA_signal_3710), .B0_t (MCOutput[1]), .B0_f (new_AGEMA_signal_3612), .B1_t (new_AGEMA_signal_3613), .B1_f (new_AGEMA_signal_3614), .Z0_t (MCOutput[33]), .Z0_f (new_AGEMA_signal_3900), .Z1_t (new_AGEMA_signal_3901), .Z1_f (new_AGEMA_signal_3902) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_2_U2 ( .A0_t (MCInst_XOR_r0_Inst_2_n1), .A0_f (new_AGEMA_signal_3954), .A1_t (new_AGEMA_signal_3955), .A1_f (new_AGEMA_signal_3956), .B0_t (MCOutput[2]), .B0_f (new_AGEMA_signal_3804), .B1_t (new_AGEMA_signal_3805), .B1_f (new_AGEMA_signal_3806), .Z0_t (MCOutput[50]), .Z0_f (new_AGEMA_signal_4029), .Z1_t (new_AGEMA_signal_4030), .Z1_f (new_AGEMA_signal_4031) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_2_U1 ( .A0_t (MCInput[50]), .A0_f (new_AGEMA_signal_3876), .A1_t (new_AGEMA_signal_3877), .A1_f (new_AGEMA_signal_3878), .B0_t (MCOutput[18]), .B0_f (new_AGEMA_signal_3828), .B1_t (new_AGEMA_signal_3829), .B1_f (new_AGEMA_signal_3830), .Z0_t (MCInst_XOR_r0_Inst_2_n1), .Z0_f (new_AGEMA_signal_3954), .Z1_t (new_AGEMA_signal_3955), .Z1_f (new_AGEMA_signal_3956) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_2_U1 ( .A0_t (MCInput[34]), .A0_f (new_AGEMA_signal_3852), .A1_t (new_AGEMA_signal_3853), .A1_f (new_AGEMA_signal_3854), .B0_t (MCOutput[2]), .B0_f (new_AGEMA_signal_3804), .B1_t (new_AGEMA_signal_3805), .B1_f (new_AGEMA_signal_3806), .Z0_t (MCOutput[34]), .Z0_f (new_AGEMA_signal_3957), .Z1_t (new_AGEMA_signal_3958), .Z1_f (new_AGEMA_signal_3959) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_3_U2 ( .A0_t (MCInst_XOR_r0_Inst_3_n1), .A0_f (new_AGEMA_signal_3903), .A1_t (new_AGEMA_signal_3904), .A1_f (new_AGEMA_signal_3905), .B0_t (MCOutput[3]), .B0_f (new_AGEMA_signal_3618), .B1_t (new_AGEMA_signal_3619), .B1_f (new_AGEMA_signal_3620), .Z0_t (MCOutput[51]), .Z0_f (new_AGEMA_signal_3960), .Z1_t (new_AGEMA_signal_3961), .Z1_f (new_AGEMA_signal_3962) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_3_U1 ( .A0_t (MCInput[51]), .A0_f (new_AGEMA_signal_3762), .A1_t (new_AGEMA_signal_3763), .A1_f (new_AGEMA_signal_3764), .B0_t (MCOutput[19]), .B0_f (new_AGEMA_signal_3666), .B1_t (new_AGEMA_signal_3667), .B1_f (new_AGEMA_signal_3668), .Z0_t (MCInst_XOR_r0_Inst_3_n1), .Z0_f (new_AGEMA_signal_3903), .Z1_t (new_AGEMA_signal_3904), .Z1_f (new_AGEMA_signal_3905) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_3_U1 ( .A0_t (MCInput[35]), .A0_f (new_AGEMA_signal_3714), .A1_t (new_AGEMA_signal_3715), .A1_f (new_AGEMA_signal_3716), .B0_t (MCOutput[3]), .B0_f (new_AGEMA_signal_3618), .B1_t (new_AGEMA_signal_3619), .B1_f (new_AGEMA_signal_3620), .Z0_t (MCOutput[35]), .Z0_f (new_AGEMA_signal_3906), .Z1_t (new_AGEMA_signal_3907), .Z1_f (new_AGEMA_signal_3908) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_4_U2 ( .A0_t (MCInst_XOR_r0_Inst_4_n1), .A0_f (new_AGEMA_signal_3963), .A1_t (new_AGEMA_signal_3964), .A1_f (new_AGEMA_signal_3965), .B0_t (MCOutput[4]), .B0_f (new_AGEMA_signal_3807), .B1_t (new_AGEMA_signal_3808), .B1_f (new_AGEMA_signal_3809), .Z0_t (MCOutput[52]), .Z0_f (new_AGEMA_signal_4032), .Z1_t (new_AGEMA_signal_4033), .Z1_f (new_AGEMA_signal_4034) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_4_U1 ( .A0_t (MCInput[52]), .A0_f (new_AGEMA_signal_3879), .A1_t (new_AGEMA_signal_3880), .A1_f (new_AGEMA_signal_3881), .B0_t (MCOutput[20]), .B0_f (new_AGEMA_signal_3831), .B1_t (new_AGEMA_signal_3832), .B1_f (new_AGEMA_signal_3833), .Z0_t (MCInst_XOR_r0_Inst_4_n1), .Z0_f (new_AGEMA_signal_3963), .Z1_t (new_AGEMA_signal_3964), .Z1_f (new_AGEMA_signal_3965) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_4_U1 ( .A0_t (MCInput[36]), .A0_f (new_AGEMA_signal_3855), .A1_t (new_AGEMA_signal_3856), .A1_f (new_AGEMA_signal_3857), .B0_t (MCOutput[4]), .B0_f (new_AGEMA_signal_3807), .B1_t (new_AGEMA_signal_3808), .B1_f (new_AGEMA_signal_3809), .Z0_t (MCOutput[36]), .Z0_f (new_AGEMA_signal_3966), .Z1_t (new_AGEMA_signal_3967), .Z1_f (new_AGEMA_signal_3968) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_5_U2 ( .A0_t (MCInst_XOR_r0_Inst_5_n1), .A0_f (new_AGEMA_signal_3909), .A1_t (new_AGEMA_signal_3910), .A1_f (new_AGEMA_signal_3911), .B0_t (MCOutput[5]), .B0_f (new_AGEMA_signal_3624), .B1_t (new_AGEMA_signal_3625), .B1_f (new_AGEMA_signal_3626), .Z0_t (MCOutput[53]), .Z0_f (new_AGEMA_signal_3969), .Z1_t (new_AGEMA_signal_3970), .Z1_f (new_AGEMA_signal_3971) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_5_U1 ( .A0_t (MCInput[53]), .A0_f (new_AGEMA_signal_3768), .A1_t (new_AGEMA_signal_3769), .A1_f (new_AGEMA_signal_3770), .B0_t (MCOutput[21]), .B0_f (new_AGEMA_signal_3672), .B1_t (new_AGEMA_signal_3673), .B1_f (new_AGEMA_signal_3674), .Z0_t (MCInst_XOR_r0_Inst_5_n1), .Z0_f (new_AGEMA_signal_3909), .Z1_t (new_AGEMA_signal_3910), .Z1_f (new_AGEMA_signal_3911) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_5_U1 ( .A0_t (MCInput[37]), .A0_f (new_AGEMA_signal_3720), .A1_t (new_AGEMA_signal_3721), .A1_f (new_AGEMA_signal_3722), .B0_t (MCOutput[5]), .B0_f (new_AGEMA_signal_3624), .B1_t (new_AGEMA_signal_3625), .B1_f (new_AGEMA_signal_3626), .Z0_t (MCOutput[37]), .Z0_f (new_AGEMA_signal_3912), .Z1_t (new_AGEMA_signal_3913), .Z1_f (new_AGEMA_signal_3914) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_6_U2 ( .A0_t (MCInst_XOR_r0_Inst_6_n1), .A0_f (new_AGEMA_signal_3972), .A1_t (new_AGEMA_signal_3973), .A1_f (new_AGEMA_signal_3974), .B0_t (MCOutput[6]), .B0_f (new_AGEMA_signal_3810), .B1_t (new_AGEMA_signal_3811), .B1_f (new_AGEMA_signal_3812), .Z0_t (MCOutput[54]), .Z0_f (new_AGEMA_signal_4035), .Z1_t (new_AGEMA_signal_4036), .Z1_f (new_AGEMA_signal_4037) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_6_U1 ( .A0_t (MCInput[54]), .A0_f (new_AGEMA_signal_3882), .A1_t (new_AGEMA_signal_3883), .A1_f (new_AGEMA_signal_3884), .B0_t (MCOutput[22]), .B0_f (new_AGEMA_signal_3834), .B1_t (new_AGEMA_signal_3835), .B1_f (new_AGEMA_signal_3836), .Z0_t (MCInst_XOR_r0_Inst_6_n1), .Z0_f (new_AGEMA_signal_3972), .Z1_t (new_AGEMA_signal_3973), .Z1_f (new_AGEMA_signal_3974) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_6_U1 ( .A0_t (MCInput[38]), .A0_f (new_AGEMA_signal_3858), .A1_t (new_AGEMA_signal_3859), .A1_f (new_AGEMA_signal_3860), .B0_t (MCOutput[6]), .B0_f (new_AGEMA_signal_3810), .B1_t (new_AGEMA_signal_3811), .B1_f (new_AGEMA_signal_3812), .Z0_t (MCOutput[38]), .Z0_f (new_AGEMA_signal_3975), .Z1_t (new_AGEMA_signal_3976), .Z1_f (new_AGEMA_signal_3977) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_7_U2 ( .A0_t (MCInst_XOR_r0_Inst_7_n1), .A0_f (new_AGEMA_signal_3915), .A1_t (new_AGEMA_signal_3916), .A1_f (new_AGEMA_signal_3917), .B0_t (MCOutput[7]), .B0_f (new_AGEMA_signal_3630), .B1_t (new_AGEMA_signal_3631), .B1_f (new_AGEMA_signal_3632), .Z0_t (MCOutput[55]), .Z0_f (new_AGEMA_signal_3978), .Z1_t (new_AGEMA_signal_3979), .Z1_f (new_AGEMA_signal_3980) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_7_U1 ( .A0_t (MCInput[55]), .A0_f (new_AGEMA_signal_3774), .A1_t (new_AGEMA_signal_3775), .A1_f (new_AGEMA_signal_3776), .B0_t (MCOutput[23]), .B0_f (new_AGEMA_signal_3678), .B1_t (new_AGEMA_signal_3679), .B1_f (new_AGEMA_signal_3680), .Z0_t (MCInst_XOR_r0_Inst_7_n1), .Z0_f (new_AGEMA_signal_3915), .Z1_t (new_AGEMA_signal_3916), .Z1_f (new_AGEMA_signal_3917) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_7_U1 ( .A0_t (MCInput[39]), .A0_f (new_AGEMA_signal_3726), .A1_t (new_AGEMA_signal_3727), .A1_f (new_AGEMA_signal_3728), .B0_t (MCOutput[7]), .B0_f (new_AGEMA_signal_3630), .B1_t (new_AGEMA_signal_3631), .B1_f (new_AGEMA_signal_3632), .Z0_t (MCOutput[39]), .Z0_f (new_AGEMA_signal_3918), .Z1_t (new_AGEMA_signal_3919), .Z1_f (new_AGEMA_signal_3920) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_8_U2 ( .A0_t (MCInst_XOR_r0_Inst_8_n1), .A0_f (new_AGEMA_signal_3981), .A1_t (new_AGEMA_signal_3982), .A1_f (new_AGEMA_signal_3983), .B0_t (MCOutput[8]), .B0_f (new_AGEMA_signal_3813), .B1_t (new_AGEMA_signal_3814), .B1_f (new_AGEMA_signal_3815), .Z0_t (MCOutput[56]), .Z0_f (new_AGEMA_signal_4038), .Z1_t (new_AGEMA_signal_4039), .Z1_f (new_AGEMA_signal_4040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_8_U1 ( .A0_t (MCInput[56]), .A0_f (new_AGEMA_signal_3885), .A1_t (new_AGEMA_signal_3886), .A1_f (new_AGEMA_signal_3887), .B0_t (MCOutput[24]), .B0_f (new_AGEMA_signal_3837), .B1_t (new_AGEMA_signal_3838), .B1_f (new_AGEMA_signal_3839), .Z0_t (MCInst_XOR_r0_Inst_8_n1), .Z0_f (new_AGEMA_signal_3981), .Z1_t (new_AGEMA_signal_3982), .Z1_f (new_AGEMA_signal_3983) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_8_U1 ( .A0_t (MCInput[40]), .A0_f (new_AGEMA_signal_3861), .A1_t (new_AGEMA_signal_3862), .A1_f (new_AGEMA_signal_3863), .B0_t (MCOutput[8]), .B0_f (new_AGEMA_signal_3813), .B1_t (new_AGEMA_signal_3814), .B1_f (new_AGEMA_signal_3815), .Z0_t (MCOutput[40]), .Z0_f (new_AGEMA_signal_3984), .Z1_t (new_AGEMA_signal_3985), .Z1_f (new_AGEMA_signal_3986) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_9_U2 ( .A0_t (MCInst_XOR_r0_Inst_9_n1), .A0_f (new_AGEMA_signal_3921), .A1_t (new_AGEMA_signal_3922), .A1_f (new_AGEMA_signal_3923), .B0_t (MCOutput[9]), .B0_f (new_AGEMA_signal_3636), .B1_t (new_AGEMA_signal_3637), .B1_f (new_AGEMA_signal_3638), .Z0_t (MCOutput[57]), .Z0_f (new_AGEMA_signal_3987), .Z1_t (new_AGEMA_signal_3988), .Z1_f (new_AGEMA_signal_3989) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_9_U1 ( .A0_t (MCInput[57]), .A0_f (new_AGEMA_signal_3780), .A1_t (new_AGEMA_signal_3781), .A1_f (new_AGEMA_signal_3782), .B0_t (MCOutput[25]), .B0_f (new_AGEMA_signal_3684), .B1_t (new_AGEMA_signal_3685), .B1_f (new_AGEMA_signal_3686), .Z0_t (MCInst_XOR_r0_Inst_9_n1), .Z0_f (new_AGEMA_signal_3921), .Z1_t (new_AGEMA_signal_3922), .Z1_f (new_AGEMA_signal_3923) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_9_U1 ( .A0_t (MCInput[41]), .A0_f (new_AGEMA_signal_3732), .A1_t (new_AGEMA_signal_3733), .A1_f (new_AGEMA_signal_3734), .B0_t (MCOutput[9]), .B0_f (new_AGEMA_signal_3636), .B1_t (new_AGEMA_signal_3637), .B1_f (new_AGEMA_signal_3638), .Z0_t (MCOutput[41]), .Z0_f (new_AGEMA_signal_3924), .Z1_t (new_AGEMA_signal_3925), .Z1_f (new_AGEMA_signal_3926) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_10_U2 ( .A0_t (MCInst_XOR_r0_Inst_10_n1), .A0_f (new_AGEMA_signal_3990), .A1_t (new_AGEMA_signal_3991), .A1_f (new_AGEMA_signal_3992), .B0_t (MCOutput[10]), .B0_f (new_AGEMA_signal_3816), .B1_t (new_AGEMA_signal_3817), .B1_f (new_AGEMA_signal_3818), .Z0_t (MCOutput[58]), .Z0_f (new_AGEMA_signal_4041), .Z1_t (new_AGEMA_signal_4042), .Z1_f (new_AGEMA_signal_4043) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_10_U1 ( .A0_t (MCInput[58]), .A0_f (new_AGEMA_signal_3888), .A1_t (new_AGEMA_signal_3889), .A1_f (new_AGEMA_signal_3890), .B0_t (MCOutput[26]), .B0_f (new_AGEMA_signal_3840), .B1_t (new_AGEMA_signal_3841), .B1_f (new_AGEMA_signal_3842), .Z0_t (MCInst_XOR_r0_Inst_10_n1), .Z0_f (new_AGEMA_signal_3990), .Z1_t (new_AGEMA_signal_3991), .Z1_f (new_AGEMA_signal_3992) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_10_U1 ( .A0_t (MCInput[42]), .A0_f (new_AGEMA_signal_3864), .A1_t (new_AGEMA_signal_3865), .A1_f (new_AGEMA_signal_3866), .B0_t (MCOutput[10]), .B0_f (new_AGEMA_signal_3816), .B1_t (new_AGEMA_signal_3817), .B1_f (new_AGEMA_signal_3818), .Z0_t (MCOutput[42]), .Z0_f (new_AGEMA_signal_3993), .Z1_t (new_AGEMA_signal_3994), .Z1_f (new_AGEMA_signal_3995) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_11_U2 ( .A0_t (MCInst_XOR_r0_Inst_11_n1), .A0_f (new_AGEMA_signal_3927), .A1_t (new_AGEMA_signal_3928), .A1_f (new_AGEMA_signal_3929), .B0_t (MCOutput[11]), .B0_f (new_AGEMA_signal_3642), .B1_t (new_AGEMA_signal_3643), .B1_f (new_AGEMA_signal_3644), .Z0_t (MCOutput[59]), .Z0_f (new_AGEMA_signal_3996), .Z1_t (new_AGEMA_signal_3997), .Z1_f (new_AGEMA_signal_3998) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_11_U1 ( .A0_t (MCInput[59]), .A0_f (new_AGEMA_signal_3786), .A1_t (new_AGEMA_signal_3787), .A1_f (new_AGEMA_signal_3788), .B0_t (MCOutput[27]), .B0_f (new_AGEMA_signal_3690), .B1_t (new_AGEMA_signal_3691), .B1_f (new_AGEMA_signal_3692), .Z0_t (MCInst_XOR_r0_Inst_11_n1), .Z0_f (new_AGEMA_signal_3927), .Z1_t (new_AGEMA_signal_3928), .Z1_f (new_AGEMA_signal_3929) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_11_U1 ( .A0_t (MCInput[43]), .A0_f (new_AGEMA_signal_3738), .A1_t (new_AGEMA_signal_3739), .A1_f (new_AGEMA_signal_3740), .B0_t (MCOutput[11]), .B0_f (new_AGEMA_signal_3642), .B1_t (new_AGEMA_signal_3643), .B1_f (new_AGEMA_signal_3644), .Z0_t (MCOutput[43]), .Z0_f (new_AGEMA_signal_3930), .Z1_t (new_AGEMA_signal_3931), .Z1_f (new_AGEMA_signal_3932) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_12_U2 ( .A0_t (MCInst_XOR_r0_Inst_12_n1), .A0_f (new_AGEMA_signal_3999), .A1_t (new_AGEMA_signal_4000), .A1_f (new_AGEMA_signal_4001), .B0_t (MCOutput[12]), .B0_f (new_AGEMA_signal_3819), .B1_t (new_AGEMA_signal_3820), .B1_f (new_AGEMA_signal_3821), .Z0_t (MCOutput[60]), .Z0_f (new_AGEMA_signal_4044), .Z1_t (new_AGEMA_signal_4045), .Z1_f (new_AGEMA_signal_4046) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_12_U1 ( .A0_t (MCInput[60]), .A0_f (new_AGEMA_signal_3891), .A1_t (new_AGEMA_signal_3892), .A1_f (new_AGEMA_signal_3893), .B0_t (MCOutput[28]), .B0_f (new_AGEMA_signal_3843), .B1_t (new_AGEMA_signal_3844), .B1_f (new_AGEMA_signal_3845), .Z0_t (MCInst_XOR_r0_Inst_12_n1), .Z0_f (new_AGEMA_signal_3999), .Z1_t (new_AGEMA_signal_4000), .Z1_f (new_AGEMA_signal_4001) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_12_U1 ( .A0_t (MCInput[44]), .A0_f (new_AGEMA_signal_3867), .A1_t (new_AGEMA_signal_3868), .A1_f (new_AGEMA_signal_3869), .B0_t (MCOutput[12]), .B0_f (new_AGEMA_signal_3819), .B1_t (new_AGEMA_signal_3820), .B1_f (new_AGEMA_signal_3821), .Z0_t (MCOutput[44]), .Z0_f (new_AGEMA_signal_4002), .Z1_t (new_AGEMA_signal_4003), .Z1_f (new_AGEMA_signal_4004) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_13_U2 ( .A0_t (MCInst_XOR_r0_Inst_13_n1), .A0_f (new_AGEMA_signal_3933), .A1_t (new_AGEMA_signal_3934), .A1_f (new_AGEMA_signal_3935), .B0_t (MCOutput[13]), .B0_f (new_AGEMA_signal_3648), .B1_t (new_AGEMA_signal_3649), .B1_f (new_AGEMA_signal_3650), .Z0_t (MCOutput[61]), .Z0_f (new_AGEMA_signal_4005), .Z1_t (new_AGEMA_signal_4006), .Z1_f (new_AGEMA_signal_4007) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_13_U1 ( .A0_t (MCInput[61]), .A0_f (new_AGEMA_signal_3792), .A1_t (new_AGEMA_signal_3793), .A1_f (new_AGEMA_signal_3794), .B0_t (MCOutput[29]), .B0_f (new_AGEMA_signal_3696), .B1_t (new_AGEMA_signal_3697), .B1_f (new_AGEMA_signal_3698), .Z0_t (MCInst_XOR_r0_Inst_13_n1), .Z0_f (new_AGEMA_signal_3933), .Z1_t (new_AGEMA_signal_3934), .Z1_f (new_AGEMA_signal_3935) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_13_U1 ( .A0_t (MCInput[45]), .A0_f (new_AGEMA_signal_3744), .A1_t (new_AGEMA_signal_3745), .A1_f (new_AGEMA_signal_3746), .B0_t (MCOutput[13]), .B0_f (new_AGEMA_signal_3648), .B1_t (new_AGEMA_signal_3649), .B1_f (new_AGEMA_signal_3650), .Z0_t (MCOutput[45]), .Z0_f (new_AGEMA_signal_3936), .Z1_t (new_AGEMA_signal_3937), .Z1_f (new_AGEMA_signal_3938) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_14_U2 ( .A0_t (MCInst_XOR_r0_Inst_14_n1), .A0_f (new_AGEMA_signal_4008), .A1_t (new_AGEMA_signal_4009), .A1_f (new_AGEMA_signal_4010), .B0_t (MCOutput[14]), .B0_f (new_AGEMA_signal_3822), .B1_t (new_AGEMA_signal_3823), .B1_f (new_AGEMA_signal_3824), .Z0_t (MCOutput[62]), .Z0_f (new_AGEMA_signal_4047), .Z1_t (new_AGEMA_signal_4048), .Z1_f (new_AGEMA_signal_4049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_14_U1 ( .A0_t (MCInput[62]), .A0_f (new_AGEMA_signal_3894), .A1_t (new_AGEMA_signal_3895), .A1_f (new_AGEMA_signal_3896), .B0_t (MCOutput[30]), .B0_f (new_AGEMA_signal_3846), .B1_t (new_AGEMA_signal_3847), .B1_f (new_AGEMA_signal_3848), .Z0_t (MCInst_XOR_r0_Inst_14_n1), .Z0_f (new_AGEMA_signal_4008), .Z1_t (new_AGEMA_signal_4009), .Z1_f (new_AGEMA_signal_4010) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_14_U1 ( .A0_t (MCInput[46]), .A0_f (new_AGEMA_signal_3870), .A1_t (new_AGEMA_signal_3871), .A1_f (new_AGEMA_signal_3872), .B0_t (MCOutput[14]), .B0_f (new_AGEMA_signal_3822), .B1_t (new_AGEMA_signal_3823), .B1_f (new_AGEMA_signal_3824), .Z0_t (MCOutput[46]), .Z0_f (new_AGEMA_signal_4011), .Z1_t (new_AGEMA_signal_4012), .Z1_f (new_AGEMA_signal_4013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_15_U2 ( .A0_t (MCInst_XOR_r0_Inst_15_n1), .A0_f (new_AGEMA_signal_3939), .A1_t (new_AGEMA_signal_3940), .A1_f (new_AGEMA_signal_3941), .B0_t (MCOutput[15]), .B0_f (new_AGEMA_signal_3654), .B1_t (new_AGEMA_signal_3655), .B1_f (new_AGEMA_signal_3656), .Z0_t (MCOutput[63]), .Z0_f (new_AGEMA_signal_4014), .Z1_t (new_AGEMA_signal_4015), .Z1_f (new_AGEMA_signal_4016) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_XOR_r0_Inst_15_U1 ( .A0_t (MCInput[63]), .A0_f (new_AGEMA_signal_3798), .A1_t (new_AGEMA_signal_3799), .A1_f (new_AGEMA_signal_3800), .B0_t (MCOutput[31]), .B0_f (new_AGEMA_signal_3702), .B1_t (new_AGEMA_signal_3703), .B1_f (new_AGEMA_signal_3704), .Z0_t (MCInst_XOR_r0_Inst_15_n1), .Z0_f (new_AGEMA_signal_3939), .Z1_t (new_AGEMA_signal_3940), .Z1_f (new_AGEMA_signal_3941) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_XOR_r1_Inst_15_U1 ( .A0_t (MCInput[47]), .A0_f (new_AGEMA_signal_3750), .A1_t (new_AGEMA_signal_3751), .A1_f (new_AGEMA_signal_3752), .B0_t (MCOutput[15]), .B0_f (new_AGEMA_signal_3654), .B1_t (new_AGEMA_signal_3655), .B1_f (new_AGEMA_signal_3656), .Z0_t (MCOutput[47]), .Z0_f (new_AGEMA_signal_3942), .Z1_t (new_AGEMA_signal_3943), .Z1_f (new_AGEMA_signal_3944) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_0_0_U1 ( .A0_t (MCOutput[48]), .A0_f (new_AGEMA_signal_4026), .A1_t (new_AGEMA_signal_4027), .A1_f (new_AGEMA_signal_4028), .B0_t (SelectedKey[48]), .B0_f (new_AGEMA_signal_2982), .B1_t (new_AGEMA_signal_2983), .B1_f (new_AGEMA_signal_2984), .Z0_t (Output_s0_t[48]), .Z0_f (Output_s0_f[48]), .Z1_t (Output_s1_t[48]), .Z1_f (Output_s1_f[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_0_1_U1 ( .A0_t (MCOutput[49]), .A0_f (new_AGEMA_signal_3951), .A1_t (new_AGEMA_signal_3952), .A1_f (new_AGEMA_signal_3953), .B0_t (SelectedKey[49]), .B0_f (new_AGEMA_signal_2985), .B1_t (new_AGEMA_signal_2986), .B1_f (new_AGEMA_signal_2987), .Z0_t (Output_s0_t[49]), .Z0_f (Output_s0_f[49]), .Z1_t (Output_s1_t[49]), .Z1_f (Output_s1_f[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_0_2_U1 ( .A0_t (MCOutput[50]), .A0_f (new_AGEMA_signal_4029), .A1_t (new_AGEMA_signal_4030), .A1_f (new_AGEMA_signal_4031), .B0_t (SelectedKey[50]), .B0_f (new_AGEMA_signal_2988), .B1_t (new_AGEMA_signal_2989), .B1_f (new_AGEMA_signal_2990), .Z0_t (Output_s0_t[50]), .Z0_f (Output_s0_f[50]), .Z1_t (Output_s1_t[50]), .Z1_f (Output_s1_f[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_0_3_U1 ( .A0_t (MCOutput[51]), .A0_f (new_AGEMA_signal_3960), .A1_t (new_AGEMA_signal_3961), .A1_f (new_AGEMA_signal_3962), .B0_t (SelectedKey[51]), .B0_f (new_AGEMA_signal_2991), .B1_t (new_AGEMA_signal_2992), .B1_f (new_AGEMA_signal_2993), .Z0_t (Output_s0_t[51]), .Z0_f (Output_s0_f[51]), .Z1_t (Output_s1_t[51]), .Z1_f (Output_s1_f[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_1_0_U1 ( .A0_t (MCOutput[52]), .A0_f (new_AGEMA_signal_4032), .A1_t (new_AGEMA_signal_4033), .A1_f (new_AGEMA_signal_4034), .B0_t (SelectedKey[52]), .B0_f (new_AGEMA_signal_2994), .B1_t (new_AGEMA_signal_2995), .B1_f (new_AGEMA_signal_2996), .Z0_t (Output_s0_t[52]), .Z0_f (Output_s0_f[52]), .Z1_t (Output_s1_t[52]), .Z1_f (Output_s1_f[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_1_1_U1 ( .A0_t (MCOutput[53]), .A0_f (new_AGEMA_signal_3969), .A1_t (new_AGEMA_signal_3970), .A1_f (new_AGEMA_signal_3971), .B0_t (SelectedKey[53]), .B0_f (new_AGEMA_signal_2997), .B1_t (new_AGEMA_signal_2998), .B1_f (new_AGEMA_signal_2999), .Z0_t (Output_s0_t[53]), .Z0_f (Output_s0_f[53]), .Z1_t (Output_s1_t[53]), .Z1_f (Output_s1_f[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_1_2_U1 ( .A0_t (MCOutput[54]), .A0_f (new_AGEMA_signal_4035), .A1_t (new_AGEMA_signal_4036), .A1_f (new_AGEMA_signal_4037), .B0_t (SelectedKey[54]), .B0_f (new_AGEMA_signal_3000), .B1_t (new_AGEMA_signal_3001), .B1_f (new_AGEMA_signal_3002), .Z0_t (Output_s0_t[54]), .Z0_f (Output_s0_f[54]), .Z1_t (Output_s1_t[54]), .Z1_f (Output_s1_f[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_1_3_U1 ( .A0_t (MCOutput[55]), .A0_f (new_AGEMA_signal_3978), .A1_t (new_AGEMA_signal_3979), .A1_f (new_AGEMA_signal_3980), .B0_t (SelectedKey[55]), .B0_f (new_AGEMA_signal_3003), .B1_t (new_AGEMA_signal_3004), .B1_f (new_AGEMA_signal_3005), .Z0_t (Output_s0_t[55]), .Z0_f (Output_s0_f[55]), .Z1_t (Output_s1_t[55]), .Z1_f (Output_s1_f[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_2_0_U1 ( .A0_t (MCOutput[56]), .A0_f (new_AGEMA_signal_4038), .A1_t (new_AGEMA_signal_4039), .A1_f (new_AGEMA_signal_4040), .B0_t (SelectedKey[56]), .B0_f (new_AGEMA_signal_3006), .B1_t (new_AGEMA_signal_3007), .B1_f (new_AGEMA_signal_3008), .Z0_t (Output_s0_t[56]), .Z0_f (Output_s0_f[56]), .Z1_t (Output_s1_t[56]), .Z1_f (Output_s1_f[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_2_1_U1 ( .A0_t (MCOutput[57]), .A0_f (new_AGEMA_signal_3987), .A1_t (new_AGEMA_signal_3988), .A1_f (new_AGEMA_signal_3989), .B0_t (SelectedKey[57]), .B0_f (new_AGEMA_signal_3009), .B1_t (new_AGEMA_signal_3010), .B1_f (new_AGEMA_signal_3011), .Z0_t (Output_s0_t[57]), .Z0_f (Output_s0_f[57]), .Z1_t (Output_s1_t[57]), .Z1_f (Output_s1_f[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_2_2_U1 ( .A0_t (MCOutput[58]), .A0_f (new_AGEMA_signal_4041), .A1_t (new_AGEMA_signal_4042), .A1_f (new_AGEMA_signal_4043), .B0_t (SelectedKey[58]), .B0_f (new_AGEMA_signal_3012), .B1_t (new_AGEMA_signal_3013), .B1_f (new_AGEMA_signal_3014), .Z0_t (Output_s0_t[58]), .Z0_f (Output_s0_f[58]), .Z1_t (Output_s1_t[58]), .Z1_f (Output_s1_f[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_2_3_U1 ( .A0_t (MCOutput[59]), .A0_f (new_AGEMA_signal_3996), .A1_t (new_AGEMA_signal_3997), .A1_f (new_AGEMA_signal_3998), .B0_t (SelectedKey[59]), .B0_f (new_AGEMA_signal_3015), .B1_t (new_AGEMA_signal_3016), .B1_f (new_AGEMA_signal_3017), .Z0_t (Output_s0_t[59]), .Z0_f (Output_s0_f[59]), .Z1_t (Output_s1_t[59]), .Z1_f (Output_s1_f[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_3_0_U1 ( .A0_t (MCOutput[60]), .A0_f (new_AGEMA_signal_4044), .A1_t (new_AGEMA_signal_4045), .A1_f (new_AGEMA_signal_4046), .B0_t (SelectedKey[60]), .B0_f (new_AGEMA_signal_3018), .B1_t (new_AGEMA_signal_3019), .B1_f (new_AGEMA_signal_3020), .Z0_t (Output_s0_t[60]), .Z0_f (Output_s0_f[60]), .Z1_t (Output_s1_t[60]), .Z1_f (Output_s1_f[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_3_1_U1 ( .A0_t (MCOutput[61]), .A0_f (new_AGEMA_signal_4005), .A1_t (new_AGEMA_signal_4006), .A1_f (new_AGEMA_signal_4007), .B0_t (SelectedKey[61]), .B0_f (new_AGEMA_signal_3021), .B1_t (new_AGEMA_signal_3022), .B1_f (new_AGEMA_signal_3023), .Z0_t (Output_s0_t[61]), .Z0_f (Output_s0_f[61]), .Z1_t (Output_s1_t[61]), .Z1_f (Output_s1_f[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_3_2_U1 ( .A0_t (MCOutput[62]), .A0_f (new_AGEMA_signal_4047), .A1_t (new_AGEMA_signal_4048), .A1_f (new_AGEMA_signal_4049), .B0_t (SelectedKey[62]), .B0_f (new_AGEMA_signal_3024), .B1_t (new_AGEMA_signal_3025), .B1_f (new_AGEMA_signal_3026), .Z0_t (Output_s0_t[62]), .Z0_f (Output_s0_f[62]), .Z1_t (Output_s1_t[62]), .Z1_f (Output_s1_f[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR1_XORInst_3_3_U1 ( .A0_t (MCOutput[63]), .A0_f (new_AGEMA_signal_4014), .A1_t (new_AGEMA_signal_4015), .A1_f (new_AGEMA_signal_4016), .B0_t (SelectedKey[63]), .B0_f (new_AGEMA_signal_3027), .B1_t (new_AGEMA_signal_3028), .B1_f (new_AGEMA_signal_3029), .Z0_t (Output_s0_t[63]), .Z0_f (Output_s0_f[63]), .Z1_t (Output_s1_t[63]), .Z1_f (Output_s1_f[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_0_0_U2 ( .A0_t (AddKeyConstXOR_XORInst_0_0_n1), .A0_f (new_AGEMA_signal_4050), .A1_t (new_AGEMA_signal_4051), .A1_f (new_AGEMA_signal_4052), .B0_t (SelectedKey[40]), .B0_f (new_AGEMA_signal_2958), .B1_t (new_AGEMA_signal_2959), .B1_f (new_AGEMA_signal_2960), .Z0_t (Output_s0_t[40]), .Z0_f (Output_s0_f[40]), .Z1_t (Output_s1_t[40]), .Z1_f (Output_s1_f[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_0_0_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (RoundConstant_0), .A1_f (new_AGEMA_signal_2194), .B0_t (MCOutput[40]), .B0_f (new_AGEMA_signal_3984), .B1_t (new_AGEMA_signal_3985), .B1_f (new_AGEMA_signal_3986), .Z0_t (AddKeyConstXOR_XORInst_0_0_n1), .Z0_f (new_AGEMA_signal_4050), .Z1_t (new_AGEMA_signal_4051), .Z1_f (new_AGEMA_signal_4052) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_0_1_U2 ( .A0_t (AddKeyConstXOR_XORInst_0_1_n1), .A0_f (new_AGEMA_signal_4017), .A1_t (new_AGEMA_signal_4018), .A1_f (new_AGEMA_signal_4019), .B0_t (SelectedKey[41]), .B0_f (new_AGEMA_signal_2961), .B1_t (new_AGEMA_signal_2962), .B1_f (new_AGEMA_signal_2963), .Z0_t (Output_s0_t[41]), .Z0_f (Output_s0_f[41]), .Z1_t (Output_s1_t[41]), .Z1_f (Output_s1_f[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_0_1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (FSMUpdate[0]), .A1_f (new_AGEMA_signal_2196), .B0_t (MCOutput[41]), .B0_f (new_AGEMA_signal_3924), .B1_t (new_AGEMA_signal_3925), .B1_f (new_AGEMA_signal_3926), .Z0_t (AddKeyConstXOR_XORInst_0_1_n1), .Z0_f (new_AGEMA_signal_4017), .Z1_t (new_AGEMA_signal_4018), .Z1_f (new_AGEMA_signal_4019) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_0_2_U2 ( .A0_t (AddKeyConstXOR_XORInst_0_2_n1), .A0_f (new_AGEMA_signal_4053), .A1_t (new_AGEMA_signal_4054), .A1_f (new_AGEMA_signal_4055), .B0_t (SelectedKey[42]), .B0_f (new_AGEMA_signal_2964), .B1_t (new_AGEMA_signal_2965), .B1_f (new_AGEMA_signal_2966), .Z0_t (Output_s0_t[42]), .Z0_f (Output_s0_f[42]), .Z1_t (Output_s1_t[42]), .Z1_f (Output_s1_f[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_0_2_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (FSMUpdate[1]), .A1_f (new_AGEMA_signal_2198), .B0_t (MCOutput[42]), .B0_f (new_AGEMA_signal_3993), .B1_t (new_AGEMA_signal_3994), .B1_f (new_AGEMA_signal_3995), .Z0_t (AddKeyConstXOR_XORInst_0_2_n1), .Z0_f (new_AGEMA_signal_4053), .Z1_t (new_AGEMA_signal_4054), .Z1_f (new_AGEMA_signal_4055) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyConstXOR_XORInst_0_3_U1 ( .A0_t (MCOutput[43]), .A0_f (new_AGEMA_signal_3930), .A1_t (new_AGEMA_signal_3931), .A1_f (new_AGEMA_signal_3932), .B0_t (SelectedKey[43]), .B0_f (new_AGEMA_signal_2967), .B1_t (new_AGEMA_signal_2968), .B1_f (new_AGEMA_signal_2969), .Z0_t (Output_s0_t[43]), .Z0_f (Output_s0_f[43]), .Z1_t (Output_s1_t[43]), .Z1_f (Output_s1_f[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_1_0_U2 ( .A0_t (AddKeyConstXOR_XORInst_1_0_n1), .A0_f (new_AGEMA_signal_4056), .A1_t (new_AGEMA_signal_4057), .A1_f (new_AGEMA_signal_4058), .B0_t (SelectedKey[44]), .B0_f (new_AGEMA_signal_2970), .B1_t (new_AGEMA_signal_2971), .B1_f (new_AGEMA_signal_2972), .Z0_t (Output_s0_t[44]), .Z0_f (Output_s0_f[44]), .Z1_t (Output_s1_t[44]), .Z1_f (Output_s1_f[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_1_0_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (RoundConstant_4_), .A1_f (new_AGEMA_signal_2200), .B0_t (MCOutput[44]), .B0_f (new_AGEMA_signal_4002), .B1_t (new_AGEMA_signal_4003), .B1_f (new_AGEMA_signal_4004), .Z0_t (AddKeyConstXOR_XORInst_1_0_n1), .Z0_f (new_AGEMA_signal_4056), .Z1_t (new_AGEMA_signal_4057), .Z1_f (new_AGEMA_signal_4058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_1_1_U2 ( .A0_t (AddKeyConstXOR_XORInst_1_1_n1), .A0_f (new_AGEMA_signal_4020), .A1_t (new_AGEMA_signal_4021), .A1_f (new_AGEMA_signal_4022), .B0_t (SelectedKey[45]), .B0_f (new_AGEMA_signal_2973), .B1_t (new_AGEMA_signal_2974), .B1_f (new_AGEMA_signal_2975), .Z0_t (Output_s0_t[45]), .Z0_f (Output_s0_f[45]), .Z1_t (Output_s1_t[45]), .Z1_f (Output_s1_f[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_1_1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (FSMUpdate[3]), .A1_f (new_AGEMA_signal_2202), .B0_t (MCOutput[45]), .B0_f (new_AGEMA_signal_3936), .B1_t (new_AGEMA_signal_3937), .B1_f (new_AGEMA_signal_3938), .Z0_t (AddKeyConstXOR_XORInst_1_1_n1), .Z0_f (new_AGEMA_signal_4020), .Z1_t (new_AGEMA_signal_4021), .Z1_f (new_AGEMA_signal_4022) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_1_2_U2 ( .A0_t (AddKeyConstXOR_XORInst_1_2_n1), .A0_f (new_AGEMA_signal_4059), .A1_t (new_AGEMA_signal_4060), .A1_f (new_AGEMA_signal_4061), .B0_t (SelectedKey[46]), .B0_f (new_AGEMA_signal_2976), .B1_t (new_AGEMA_signal_2977), .B1_f (new_AGEMA_signal_2978), .Z0_t (Output_s0_t[46]), .Z0_f (Output_s0_f[46]), .Z1_t (Output_s1_t[46]), .Z1_f (Output_s1_f[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_1_2_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (FSMUpdate[4]), .A1_f (new_AGEMA_signal_2204), .B0_t (MCOutput[46]), .B0_f (new_AGEMA_signal_4011), .B1_t (new_AGEMA_signal_4012), .B1_f (new_AGEMA_signal_4013), .Z0_t (AddKeyConstXOR_XORInst_1_2_n1), .Z0_f (new_AGEMA_signal_4059), .Z1_t (new_AGEMA_signal_4060), .Z1_f (new_AGEMA_signal_4061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) AddKeyConstXOR_XORInst_1_3_U2 ( .A0_t (AddKeyConstXOR_XORInst_1_3_n1), .A0_f (new_AGEMA_signal_4023), .A1_t (new_AGEMA_signal_4024), .A1_f (new_AGEMA_signal_4025), .B0_t (SelectedKey[47]), .B0_f (new_AGEMA_signal_2979), .B1_t (new_AGEMA_signal_2980), .B1_f (new_AGEMA_signal_2981), .Z0_t (Output_s0_t[47]), .Z0_f (Output_s0_f[47]), .Z1_t (Output_s1_t[47]), .Z1_f (Output_s1_f[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) AddKeyConstXOR_XORInst_1_3_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (FSMUpdate[5]), .A1_f (new_AGEMA_signal_2206), .B0_t (MCOutput[47]), .B0_f (new_AGEMA_signal_3942), .B1_t (new_AGEMA_signal_3943), .B1_f (new_AGEMA_signal_3944), .Z0_t (AddKeyConstXOR_XORInst_1_3_n1), .Z0_f (new_AGEMA_signal_4023), .Z1_t (new_AGEMA_signal_4024), .Z1_f (new_AGEMA_signal_4025) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_0_0_U1 ( .A0_t (MCOutput[0]), .A0_f (new_AGEMA_signal_3801), .A1_t (new_AGEMA_signal_3802), .A1_f (new_AGEMA_signal_3803), .B0_t (SelectedKey[0]), .B0_f (new_AGEMA_signal_2838), .B1_t (new_AGEMA_signal_2839), .B1_f (new_AGEMA_signal_2840), .Z0_t (Output_s0_t[0]), .Z0_f (Output_s0_f[0]), .Z1_t (Output_s1_t[0]), .Z1_f (Output_s1_f[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_0_1_U1 ( .A0_t (MCOutput[1]), .A0_f (new_AGEMA_signal_3612), .A1_t (new_AGEMA_signal_3613), .A1_f (new_AGEMA_signal_3614), .B0_t (SelectedKey[1]), .B0_f (new_AGEMA_signal_2841), .B1_t (new_AGEMA_signal_2842), .B1_f (new_AGEMA_signal_2843), .Z0_t (Output_s0_t[1]), .Z0_f (Output_s0_f[1]), .Z1_t (Output_s1_t[1]), .Z1_f (Output_s1_f[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_0_2_U1 ( .A0_t (MCOutput[2]), .A0_f (new_AGEMA_signal_3804), .A1_t (new_AGEMA_signal_3805), .A1_f (new_AGEMA_signal_3806), .B0_t (SelectedKey[2]), .B0_f (new_AGEMA_signal_2844), .B1_t (new_AGEMA_signal_2845), .B1_f (new_AGEMA_signal_2846), .Z0_t (Output_s0_t[2]), .Z0_f (Output_s0_f[2]), .Z1_t (Output_s1_t[2]), .Z1_f (Output_s1_f[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_0_3_U1 ( .A0_t (MCOutput[3]), .A0_f (new_AGEMA_signal_3618), .A1_t (new_AGEMA_signal_3619), .A1_f (new_AGEMA_signal_3620), .B0_t (SelectedKey[3]), .B0_f (new_AGEMA_signal_2847), .B1_t (new_AGEMA_signal_2848), .B1_f (new_AGEMA_signal_2849), .Z0_t (Output_s0_t[3]), .Z0_f (Output_s0_f[3]), .Z1_t (Output_s1_t[3]), .Z1_f (Output_s1_f[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_1_0_U1 ( .A0_t (MCOutput[4]), .A0_f (new_AGEMA_signal_3807), .A1_t (new_AGEMA_signal_3808), .A1_f (new_AGEMA_signal_3809), .B0_t (SelectedKey[4]), .B0_f (new_AGEMA_signal_2850), .B1_t (new_AGEMA_signal_2851), .B1_f (new_AGEMA_signal_2852), .Z0_t (Output_s0_t[4]), .Z0_f (Output_s0_f[4]), .Z1_t (Output_s1_t[4]), .Z1_f (Output_s1_f[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_1_1_U1 ( .A0_t (MCOutput[5]), .A0_f (new_AGEMA_signal_3624), .A1_t (new_AGEMA_signal_3625), .A1_f (new_AGEMA_signal_3626), .B0_t (SelectedKey[5]), .B0_f (new_AGEMA_signal_2853), .B1_t (new_AGEMA_signal_2854), .B1_f (new_AGEMA_signal_2855), .Z0_t (Output_s0_t[5]), .Z0_f (Output_s0_f[5]), .Z1_t (Output_s1_t[5]), .Z1_f (Output_s1_f[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_1_2_U1 ( .A0_t (MCOutput[6]), .A0_f (new_AGEMA_signal_3810), .A1_t (new_AGEMA_signal_3811), .A1_f (new_AGEMA_signal_3812), .B0_t (SelectedKey[6]), .B0_f (new_AGEMA_signal_2856), .B1_t (new_AGEMA_signal_2857), .B1_f (new_AGEMA_signal_2858), .Z0_t (Output_s0_t[6]), .Z0_f (Output_s0_f[6]), .Z1_t (Output_s1_t[6]), .Z1_f (Output_s1_f[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_1_3_U1 ( .A0_t (MCOutput[7]), .A0_f (new_AGEMA_signal_3630), .A1_t (new_AGEMA_signal_3631), .A1_f (new_AGEMA_signal_3632), .B0_t (SelectedKey[7]), .B0_f (new_AGEMA_signal_2859), .B1_t (new_AGEMA_signal_2860), .B1_f (new_AGEMA_signal_2861), .Z0_t (Output_s0_t[7]), .Z0_f (Output_s0_f[7]), .Z1_t (Output_s1_t[7]), .Z1_f (Output_s1_f[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_2_0_U1 ( .A0_t (MCOutput[8]), .A0_f (new_AGEMA_signal_3813), .A1_t (new_AGEMA_signal_3814), .A1_f (new_AGEMA_signal_3815), .B0_t (SelectedKey[8]), .B0_f (new_AGEMA_signal_2862), .B1_t (new_AGEMA_signal_2863), .B1_f (new_AGEMA_signal_2864), .Z0_t (Output_s0_t[8]), .Z0_f (Output_s0_f[8]), .Z1_t (Output_s1_t[8]), .Z1_f (Output_s1_f[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_2_1_U1 ( .A0_t (MCOutput[9]), .A0_f (new_AGEMA_signal_3636), .A1_t (new_AGEMA_signal_3637), .A1_f (new_AGEMA_signal_3638), .B0_t (SelectedKey[9]), .B0_f (new_AGEMA_signal_2865), .B1_t (new_AGEMA_signal_2866), .B1_f (new_AGEMA_signal_2867), .Z0_t (Output_s0_t[9]), .Z0_f (Output_s0_f[9]), .Z1_t (Output_s1_t[9]), .Z1_f (Output_s1_f[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_2_2_U1 ( .A0_t (MCOutput[10]), .A0_f (new_AGEMA_signal_3816), .A1_t (new_AGEMA_signal_3817), .A1_f (new_AGEMA_signal_3818), .B0_t (SelectedKey[10]), .B0_f (new_AGEMA_signal_2868), .B1_t (new_AGEMA_signal_2869), .B1_f (new_AGEMA_signal_2870), .Z0_t (Output_s0_t[10]), .Z0_f (Output_s0_f[10]), .Z1_t (Output_s1_t[10]), .Z1_f (Output_s1_f[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_2_3_U1 ( .A0_t (MCOutput[11]), .A0_f (new_AGEMA_signal_3642), .A1_t (new_AGEMA_signal_3643), .A1_f (new_AGEMA_signal_3644), .B0_t (SelectedKey[11]), .B0_f (new_AGEMA_signal_2871), .B1_t (new_AGEMA_signal_2872), .B1_f (new_AGEMA_signal_2873), .Z0_t (Output_s0_t[11]), .Z0_f (Output_s0_f[11]), .Z1_t (Output_s1_t[11]), .Z1_f (Output_s1_f[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_3_0_U1 ( .A0_t (MCOutput[12]), .A0_f (new_AGEMA_signal_3819), .A1_t (new_AGEMA_signal_3820), .A1_f (new_AGEMA_signal_3821), .B0_t (SelectedKey[12]), .B0_f (new_AGEMA_signal_2874), .B1_t (new_AGEMA_signal_2875), .B1_f (new_AGEMA_signal_2876), .Z0_t (Output_s0_t[12]), .Z0_f (Output_s0_f[12]), .Z1_t (Output_s1_t[12]), .Z1_f (Output_s1_f[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_3_1_U1 ( .A0_t (MCOutput[13]), .A0_f (new_AGEMA_signal_3648), .A1_t (new_AGEMA_signal_3649), .A1_f (new_AGEMA_signal_3650), .B0_t (SelectedKey[13]), .B0_f (new_AGEMA_signal_2877), .B1_t (new_AGEMA_signal_2878), .B1_f (new_AGEMA_signal_2879), .Z0_t (Output_s0_t[13]), .Z0_f (Output_s0_f[13]), .Z1_t (Output_s1_t[13]), .Z1_f (Output_s1_f[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_3_2_U1 ( .A0_t (MCOutput[14]), .A0_f (new_AGEMA_signal_3822), .A1_t (new_AGEMA_signal_3823), .A1_f (new_AGEMA_signal_3824), .B0_t (SelectedKey[14]), .B0_f (new_AGEMA_signal_2880), .B1_t (new_AGEMA_signal_2881), .B1_f (new_AGEMA_signal_2882), .Z0_t (Output_s0_t[14]), .Z0_f (Output_s0_f[14]), .Z1_t (Output_s1_t[14]), .Z1_f (Output_s1_f[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_3_3_U1 ( .A0_t (MCOutput[15]), .A0_f (new_AGEMA_signal_3654), .A1_t (new_AGEMA_signal_3655), .A1_f (new_AGEMA_signal_3656), .B0_t (SelectedKey[15]), .B0_f (new_AGEMA_signal_2883), .B1_t (new_AGEMA_signal_2884), .B1_f (new_AGEMA_signal_2885), .Z0_t (Output_s0_t[15]), .Z0_f (Output_s0_f[15]), .Z1_t (Output_s1_t[15]), .Z1_f (Output_s1_f[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_4_0_U1 ( .A0_t (MCOutput[16]), .A0_f (new_AGEMA_signal_3825), .A1_t (new_AGEMA_signal_3826), .A1_f (new_AGEMA_signal_3827), .B0_t (SelectedKey[16]), .B0_f (new_AGEMA_signal_2886), .B1_t (new_AGEMA_signal_2887), .B1_f (new_AGEMA_signal_2888), .Z0_t (Output_s0_t[16]), .Z0_f (Output_s0_f[16]), .Z1_t (Output_s1_t[16]), .Z1_f (Output_s1_f[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_4_1_U1 ( .A0_t (MCOutput[17]), .A0_f (new_AGEMA_signal_3660), .A1_t (new_AGEMA_signal_3661), .A1_f (new_AGEMA_signal_3662), .B0_t (SelectedKey[17]), .B0_f (new_AGEMA_signal_2889), .B1_t (new_AGEMA_signal_2890), .B1_f (new_AGEMA_signal_2891), .Z0_t (Output_s0_t[17]), .Z0_f (Output_s0_f[17]), .Z1_t (Output_s1_t[17]), .Z1_f (Output_s1_f[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_4_2_U1 ( .A0_t (MCOutput[18]), .A0_f (new_AGEMA_signal_3828), .A1_t (new_AGEMA_signal_3829), .A1_f (new_AGEMA_signal_3830), .B0_t (SelectedKey[18]), .B0_f (new_AGEMA_signal_2892), .B1_t (new_AGEMA_signal_2893), .B1_f (new_AGEMA_signal_2894), .Z0_t (Output_s0_t[18]), .Z0_f (Output_s0_f[18]), .Z1_t (Output_s1_t[18]), .Z1_f (Output_s1_f[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_4_3_U1 ( .A0_t (MCOutput[19]), .A0_f (new_AGEMA_signal_3666), .A1_t (new_AGEMA_signal_3667), .A1_f (new_AGEMA_signal_3668), .B0_t (SelectedKey[19]), .B0_f (new_AGEMA_signal_2895), .B1_t (new_AGEMA_signal_2896), .B1_f (new_AGEMA_signal_2897), .Z0_t (Output_s0_t[19]), .Z0_f (Output_s0_f[19]), .Z1_t (Output_s1_t[19]), .Z1_f (Output_s1_f[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_5_0_U1 ( .A0_t (MCOutput[20]), .A0_f (new_AGEMA_signal_3831), .A1_t (new_AGEMA_signal_3832), .A1_f (new_AGEMA_signal_3833), .B0_t (SelectedKey[20]), .B0_f (new_AGEMA_signal_2898), .B1_t (new_AGEMA_signal_2899), .B1_f (new_AGEMA_signal_2900), .Z0_t (Output_s0_t[20]), .Z0_f (Output_s0_f[20]), .Z1_t (Output_s1_t[20]), .Z1_f (Output_s1_f[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_5_1_U1 ( .A0_t (MCOutput[21]), .A0_f (new_AGEMA_signal_3672), .A1_t (new_AGEMA_signal_3673), .A1_f (new_AGEMA_signal_3674), .B0_t (SelectedKey[21]), .B0_f (new_AGEMA_signal_2901), .B1_t (new_AGEMA_signal_2902), .B1_f (new_AGEMA_signal_2903), .Z0_t (Output_s0_t[21]), .Z0_f (Output_s0_f[21]), .Z1_t (Output_s1_t[21]), .Z1_f (Output_s1_f[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_5_2_U1 ( .A0_t (MCOutput[22]), .A0_f (new_AGEMA_signal_3834), .A1_t (new_AGEMA_signal_3835), .A1_f (new_AGEMA_signal_3836), .B0_t (SelectedKey[22]), .B0_f (new_AGEMA_signal_2904), .B1_t (new_AGEMA_signal_2905), .B1_f (new_AGEMA_signal_2906), .Z0_t (Output_s0_t[22]), .Z0_f (Output_s0_f[22]), .Z1_t (Output_s1_t[22]), .Z1_f (Output_s1_f[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_5_3_U1 ( .A0_t (MCOutput[23]), .A0_f (new_AGEMA_signal_3678), .A1_t (new_AGEMA_signal_3679), .A1_f (new_AGEMA_signal_3680), .B0_t (SelectedKey[23]), .B0_f (new_AGEMA_signal_2907), .B1_t (new_AGEMA_signal_2908), .B1_f (new_AGEMA_signal_2909), .Z0_t (Output_s0_t[23]), .Z0_f (Output_s0_f[23]), .Z1_t (Output_s1_t[23]), .Z1_f (Output_s1_f[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_6_0_U1 ( .A0_t (MCOutput[24]), .A0_f (new_AGEMA_signal_3837), .A1_t (new_AGEMA_signal_3838), .A1_f (new_AGEMA_signal_3839), .B0_t (SelectedKey[24]), .B0_f (new_AGEMA_signal_2910), .B1_t (new_AGEMA_signal_2911), .B1_f (new_AGEMA_signal_2912), .Z0_t (Output_s0_t[24]), .Z0_f (Output_s0_f[24]), .Z1_t (Output_s1_t[24]), .Z1_f (Output_s1_f[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_6_1_U1 ( .A0_t (MCOutput[25]), .A0_f (new_AGEMA_signal_3684), .A1_t (new_AGEMA_signal_3685), .A1_f (new_AGEMA_signal_3686), .B0_t (SelectedKey[25]), .B0_f (new_AGEMA_signal_2913), .B1_t (new_AGEMA_signal_2914), .B1_f (new_AGEMA_signal_2915), .Z0_t (Output_s0_t[25]), .Z0_f (Output_s0_f[25]), .Z1_t (Output_s1_t[25]), .Z1_f (Output_s1_f[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_6_2_U1 ( .A0_t (MCOutput[26]), .A0_f (new_AGEMA_signal_3840), .A1_t (new_AGEMA_signal_3841), .A1_f (new_AGEMA_signal_3842), .B0_t (SelectedKey[26]), .B0_f (new_AGEMA_signal_2916), .B1_t (new_AGEMA_signal_2917), .B1_f (new_AGEMA_signal_2918), .Z0_t (Output_s0_t[26]), .Z0_f (Output_s0_f[26]), .Z1_t (Output_s1_t[26]), .Z1_f (Output_s1_f[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_6_3_U1 ( .A0_t (MCOutput[27]), .A0_f (new_AGEMA_signal_3690), .A1_t (new_AGEMA_signal_3691), .A1_f (new_AGEMA_signal_3692), .B0_t (SelectedKey[27]), .B0_f (new_AGEMA_signal_2919), .B1_t (new_AGEMA_signal_2920), .B1_f (new_AGEMA_signal_2921), .Z0_t (Output_s0_t[27]), .Z0_f (Output_s0_f[27]), .Z1_t (Output_s1_t[27]), .Z1_f (Output_s1_f[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_7_0_U1 ( .A0_t (MCOutput[28]), .A0_f (new_AGEMA_signal_3843), .A1_t (new_AGEMA_signal_3844), .A1_f (new_AGEMA_signal_3845), .B0_t (SelectedKey[28]), .B0_f (new_AGEMA_signal_2922), .B1_t (new_AGEMA_signal_2923), .B1_f (new_AGEMA_signal_2924), .Z0_t (Output_s0_t[28]), .Z0_f (Output_s0_f[28]), .Z1_t (Output_s1_t[28]), .Z1_f (Output_s1_f[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_7_1_U1 ( .A0_t (MCOutput[29]), .A0_f (new_AGEMA_signal_3696), .A1_t (new_AGEMA_signal_3697), .A1_f (new_AGEMA_signal_3698), .B0_t (SelectedKey[29]), .B0_f (new_AGEMA_signal_2925), .B1_t (new_AGEMA_signal_2926), .B1_f (new_AGEMA_signal_2927), .Z0_t (Output_s0_t[29]), .Z0_f (Output_s0_f[29]), .Z1_t (Output_s1_t[29]), .Z1_f (Output_s1_f[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_7_2_U1 ( .A0_t (MCOutput[30]), .A0_f (new_AGEMA_signal_3846), .A1_t (new_AGEMA_signal_3847), .A1_f (new_AGEMA_signal_3848), .B0_t (SelectedKey[30]), .B0_f (new_AGEMA_signal_2928), .B1_t (new_AGEMA_signal_2929), .B1_f (new_AGEMA_signal_2930), .Z0_t (Output_s0_t[30]), .Z0_f (Output_s0_f[30]), .Z1_t (Output_s1_t[30]), .Z1_f (Output_s1_f[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_7_3_U1 ( .A0_t (MCOutput[31]), .A0_f (new_AGEMA_signal_3702), .A1_t (new_AGEMA_signal_3703), .A1_f (new_AGEMA_signal_3704), .B0_t (SelectedKey[31]), .B0_f (new_AGEMA_signal_2931), .B1_t (new_AGEMA_signal_2932), .B1_f (new_AGEMA_signal_2933), .Z0_t (Output_s0_t[31]), .Z0_f (Output_s0_f[31]), .Z1_t (Output_s1_t[31]), .Z1_f (Output_s1_f[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_8_0_U1 ( .A0_t (MCOutput[32]), .A0_f (new_AGEMA_signal_3948), .A1_t (new_AGEMA_signal_3949), .A1_f (new_AGEMA_signal_3950), .B0_t (SelectedKey[32]), .B0_f (new_AGEMA_signal_2934), .B1_t (new_AGEMA_signal_2935), .B1_f (new_AGEMA_signal_2936), .Z0_t (Output_s0_t[32]), .Z0_f (Output_s0_f[32]), .Z1_t (Output_s1_t[32]), .Z1_f (Output_s1_f[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_8_1_U1 ( .A0_t (MCOutput[33]), .A0_f (new_AGEMA_signal_3900), .A1_t (new_AGEMA_signal_3901), .A1_f (new_AGEMA_signal_3902), .B0_t (SelectedKey[33]), .B0_f (new_AGEMA_signal_2937), .B1_t (new_AGEMA_signal_2938), .B1_f (new_AGEMA_signal_2939), .Z0_t (Output_s0_t[33]), .Z0_f (Output_s0_f[33]), .Z1_t (Output_s1_t[33]), .Z1_f (Output_s1_f[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_8_2_U1 ( .A0_t (MCOutput[34]), .A0_f (new_AGEMA_signal_3957), .A1_t (new_AGEMA_signal_3958), .A1_f (new_AGEMA_signal_3959), .B0_t (SelectedKey[34]), .B0_f (new_AGEMA_signal_2940), .B1_t (new_AGEMA_signal_2941), .B1_f (new_AGEMA_signal_2942), .Z0_t (Output_s0_t[34]), .Z0_f (Output_s0_f[34]), .Z1_t (Output_s1_t[34]), .Z1_f (Output_s1_f[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_8_3_U1 ( .A0_t (MCOutput[35]), .A0_f (new_AGEMA_signal_3906), .A1_t (new_AGEMA_signal_3907), .A1_f (new_AGEMA_signal_3908), .B0_t (SelectedKey[35]), .B0_f (new_AGEMA_signal_2943), .B1_t (new_AGEMA_signal_2944), .B1_f (new_AGEMA_signal_2945), .Z0_t (Output_s0_t[35]), .Z0_f (Output_s0_f[35]), .Z1_t (Output_s1_t[35]), .Z1_f (Output_s1_f[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_9_0_U1 ( .A0_t (MCOutput[36]), .A0_f (new_AGEMA_signal_3966), .A1_t (new_AGEMA_signal_3967), .A1_f (new_AGEMA_signal_3968), .B0_t (SelectedKey[36]), .B0_f (new_AGEMA_signal_2946), .B1_t (new_AGEMA_signal_2947), .B1_f (new_AGEMA_signal_2948), .Z0_t (Output_s0_t[36]), .Z0_f (Output_s0_f[36]), .Z1_t (Output_s1_t[36]), .Z1_f (Output_s1_f[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_9_1_U1 ( .A0_t (MCOutput[37]), .A0_f (new_AGEMA_signal_3912), .A1_t (new_AGEMA_signal_3913), .A1_f (new_AGEMA_signal_3914), .B0_t (SelectedKey[37]), .B0_f (new_AGEMA_signal_2949), .B1_t (new_AGEMA_signal_2950), .B1_f (new_AGEMA_signal_2951), .Z0_t (Output_s0_t[37]), .Z0_f (Output_s0_f[37]), .Z1_t (Output_s1_t[37]), .Z1_f (Output_s1_f[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_9_2_U1 ( .A0_t (MCOutput[38]), .A0_f (new_AGEMA_signal_3975), .A1_t (new_AGEMA_signal_3976), .A1_f (new_AGEMA_signal_3977), .B0_t (SelectedKey[38]), .B0_f (new_AGEMA_signal_2952), .B1_t (new_AGEMA_signal_2953), .B1_f (new_AGEMA_signal_2954), .Z0_t (Output_s0_t[38]), .Z0_f (Output_s0_f[38]), .Z1_t (Output_s1_t[38]), .Z1_f (Output_s1_f[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) AddKeyXOR2_XORInst_9_3_U1 ( .A0_t (MCOutput[39]), .A0_f (new_AGEMA_signal_3918), .A1_t (new_AGEMA_signal_3919), .A1_f (new_AGEMA_signal_3920), .B0_t (SelectedKey[39]), .B0_f (new_AGEMA_signal_2955), .B1_t (new_AGEMA_signal_2956), .B1_f (new_AGEMA_signal_2957), .Z0_t (Output_s0_t[39]), .Z0_f (Output_s0_f[39]), .Z1_t (Output_s1_t[39]), .Z1_f (Output_s1_f[39]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_U19 ( .A0_t (SubCellInst_SboxInst_0_n15), .A0_f (new_AGEMA_signal_2646), .A1_t (new_AGEMA_signal_2647), .A1_f (new_AGEMA_signal_2648), .B0_t (SubCellInst_SboxInst_0_n14), .B0_f (new_AGEMA_signal_1205), .B1_t (new_AGEMA_signal_1206), .B1_f (new_AGEMA_signal_1207), .Z0_t (Feedback[0]), .Z0_f (new_AGEMA_signal_3223), .Z1_t (new_AGEMA_signal_3224), .Z1_f (new_AGEMA_signal_3225) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_U18 ( .A0_t (Output_s0_t[61]), .A0_f (Output_s0_f[61]), .A1_t (Output_s1_t[61]), .A1_f (Output_s1_f[61]), .B0_t (SubCellInst_SboxInst_0_n13), .B0_f (new_AGEMA_signal_2211), .B1_t (new_AGEMA_signal_2212), .B1_f (new_AGEMA_signal_2213), .Z0_t (SubCellInst_SboxInst_0_n15), .Z0_f (new_AGEMA_signal_2646), .Z1_t (new_AGEMA_signal_2647), .Z1_f (new_AGEMA_signal_2648) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_U17 ( .A0_t (Output_s0_t[60]), .A0_f (Output_s0_f[60]), .A1_t (Output_s1_t[60]), .A1_f (Output_s1_f[60]), .B0_t (SubCellInst_SboxInst_0_n11), .B0_f (new_AGEMA_signal_1190), .B1_t (new_AGEMA_signal_1191), .B1_f (new_AGEMA_signal_1192), .Z0_t (SubCellInst_SboxInst_0_n13), .Z0_f (new_AGEMA_signal_2211), .Z1_t (new_AGEMA_signal_2212), .Z1_f (new_AGEMA_signal_2213) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_U16 ( .A0_t (Output_s0_t[62]), .A0_f (Output_s0_f[62]), .A1_t (Output_s1_t[62]), .A1_f (Output_s1_f[62]), .B0_t (Output_s0_t[63]), .B0_f (Output_s0_f[63]), .B1_t (Output_s1_t[63]), .B1_f (Output_s1_f[63]), .Z0_t (SubCellInst_SboxInst_0_n11), .Z0_f (new_AGEMA_signal_1190), .Z1_t (new_AGEMA_signal_1191), .Z1_f (new_AGEMA_signal_1192) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U15 ( .A0_t (SubCellInst_SboxInst_0_n10), .A0_f (new_AGEMA_signal_2214), .A1_t (new_AGEMA_signal_2215), .A1_f (new_AGEMA_signal_2216), .B0_t (SubCellInst_SboxInst_0_n9), .B0_f (new_AGEMA_signal_1196), .B1_t (new_AGEMA_signal_1197), .B1_f (new_AGEMA_signal_1198), .Z0_t (Feedback[1]), .Z0_f (new_AGEMA_signal_2649), .Z1_t (new_AGEMA_signal_2650), .Z1_f (new_AGEMA_signal_2651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U14 ( .A0_t (Output_s0_t[60]), .A0_f (Output_s0_f[60]), .A1_t (Output_s1_t[60]), .A1_f (Output_s1_f[60]), .B0_t (Output_s0_t[63]), .B0_f (Output_s0_f[63]), .B1_t (Output_s1_t[63]), .B1_f (Output_s1_f[63]), .Z0_t (SubCellInst_SboxInst_0_n9), .Z0_f (new_AGEMA_signal_1196), .Z1_t (new_AGEMA_signal_1197), .Z1_f (new_AGEMA_signal_1198) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U13 ( .A0_t (Output_s0_t[62]), .A0_f (Output_s0_f[62]), .A1_t (Output_s1_t[62]), .A1_f (Output_s1_f[62]), .B0_t (SubCellInst_SboxInst_0_n7), .B0_f (new_AGEMA_signal_1199), .B1_t (new_AGEMA_signal_1200), .B1_f (new_AGEMA_signal_1201), .Z0_t (SubCellInst_SboxInst_0_n10), .Z0_f (new_AGEMA_signal_2214), .Z1_t (new_AGEMA_signal_2215), .Z1_f (new_AGEMA_signal_2216) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U12 ( .A0_t (Output_s0_t[63]), .A0_f (Output_s0_f[63]), .A1_t (Output_s1_t[63]), .A1_f (Output_s1_f[63]), .B0_t (Output_s0_t[60]), .B0_f (Output_s0_f[60]), .B1_t (Output_s1_t[60]), .B1_f (Output_s1_f[60]), .Z0_t (SubCellInst_SboxInst_0_n7), .Z0_f (new_AGEMA_signal_1199), .Z1_t (new_AGEMA_signal_1200), .Z1_f (new_AGEMA_signal_1201) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U11 ( .A0_t (SubCellInst_SboxInst_0_n6), .A0_f (new_AGEMA_signal_2652), .A1_t (new_AGEMA_signal_2653), .A1_f (new_AGEMA_signal_2654), .B0_t (SubCellInst_SboxInst_0_n5), .B0_f (new_AGEMA_signal_1208), .B1_t (new_AGEMA_signal_1209), .B1_f (new_AGEMA_signal_1210), .Z0_t (Feedback[2]), .Z0_f (new_AGEMA_signal_3226), .Z1_t (new_AGEMA_signal_3227), .Z1_f (new_AGEMA_signal_3228) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U10 ( .A0_t (SubCellInst_SboxInst_0_n4), .A0_f (new_AGEMA_signal_2217), .A1_t (new_AGEMA_signal_2218), .A1_f (new_AGEMA_signal_2219), .B0_t (Output_s0_t[61]), .B0_f (Output_s0_f[61]), .B1_t (Output_s1_t[61]), .B1_f (Output_s1_f[61]), .Z0_t (SubCellInst_SboxInst_0_n6), .Z0_f (new_AGEMA_signal_2652), .Z1_t (new_AGEMA_signal_2653), .Z1_f (new_AGEMA_signal_2654) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U9 ( .A0_t (SubCellInst_SboxInst_0_n3), .A0_f (new_AGEMA_signal_1202), .A1_t (new_AGEMA_signal_1203), .A1_f (new_AGEMA_signal_1204), .B0_t (Output_s0_t[62]), .B0_f (Output_s0_f[62]), .B1_t (Output_s1_t[62]), .B1_f (Output_s1_f[62]), .Z0_t (SubCellInst_SboxInst_0_n4), .Z0_f (new_AGEMA_signal_2217), .Z1_t (new_AGEMA_signal_2218), .Z1_f (new_AGEMA_signal_2219) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U8 ( .A0_t (Output_s0_t[60]), .A0_f (Output_s0_f[60]), .A1_t (Output_s1_t[60]), .A1_f (Output_s1_f[60]), .B0_t (Output_s0_t[63]), .B0_f (Output_s0_f[63]), .B1_t (Output_s1_t[63]), .B1_f (Output_s1_f[63]), .Z0_t (SubCellInst_SboxInst_0_n3), .Z0_f (new_AGEMA_signal_1202), .Z1_t (new_AGEMA_signal_1203), .Z1_f (new_AGEMA_signal_1204) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U7 ( .A0_t (SubCellInst_SboxInst_0_n5), .A0_f (new_AGEMA_signal_1208), .A1_t (new_AGEMA_signal_1209), .A1_f (new_AGEMA_signal_1210), .B0_t (SubCellInst_SboxInst_0_n1), .B0_f (new_AGEMA_signal_2223), .B1_t (new_AGEMA_signal_2224), .B1_f (new_AGEMA_signal_2225), .Z0_t (Feedback[3]), .Z0_f (new_AGEMA_signal_2655), .Z1_t (new_AGEMA_signal_2656), .Z1_f (new_AGEMA_signal_2657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U6 ( .A0_t (Output_s0_t[61]), .A0_f (Output_s0_f[61]), .A1_t (Output_s1_t[61]), .A1_f (Output_s1_f[61]), .B0_t (SubCellInst_SboxInst_0_n14), .B0_f (new_AGEMA_signal_1205), .B1_t (new_AGEMA_signal_1206), .B1_f (new_AGEMA_signal_1207), .Z0_t (SubCellInst_SboxInst_0_n1), .Z0_f (new_AGEMA_signal_2223), .Z1_t (new_AGEMA_signal_2224), .Z1_f (new_AGEMA_signal_2225) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_U5 ( .A0_t (Output_s0_t[62]), .A0_f (Output_s0_f[62]), .A1_t (Output_s1_t[62]), .A1_f (Output_s1_f[62]), .B0_t (Output_s0_t[63]), .B0_f (Output_s0_f[63]), .B1_t (Output_s1_t[63]), .B1_f (Output_s1_f[63]), .Z0_t (SubCellInst_SboxInst_0_n14), .Z0_f (new_AGEMA_signal_1205), .Z1_t (new_AGEMA_signal_1206), .Z1_f (new_AGEMA_signal_1207) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_U3 ( .A0_t (Output_s0_t[63]), .A0_f (Output_s0_f[63]), .A1_t (Output_s1_t[63]), .A1_f (Output_s1_f[63]), .B0_t (Output_s0_t[60]), .B0_f (Output_s0_f[60]), .B1_t (Output_s1_t[60]), .B1_f (Output_s1_f[60]), .Z0_t (SubCellInst_SboxInst_0_n5), .Z0_f (new_AGEMA_signal_1208), .Z1_t (new_AGEMA_signal_1209), .Z1_f (new_AGEMA_signal_1210) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_U19 ( .A0_t (SubCellInst_SboxInst_1_n15), .A0_f (new_AGEMA_signal_2658), .A1_t (new_AGEMA_signal_2659), .A1_f (new_AGEMA_signal_2660), .B0_t (SubCellInst_SboxInst_1_n14), .B0_f (new_AGEMA_signal_1232), .B1_t (new_AGEMA_signal_1233), .B1_f (new_AGEMA_signal_1234), .Z0_t (Feedback[4]), .Z0_f (new_AGEMA_signal_3229), .Z1_t (new_AGEMA_signal_3230), .Z1_f (new_AGEMA_signal_3231) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_U18 ( .A0_t (Output_s0_t[49]), .A0_f (Output_s0_f[49]), .A1_t (Output_s1_t[49]), .A1_f (Output_s1_f[49]), .B0_t (SubCellInst_SboxInst_1_n13), .B0_f (new_AGEMA_signal_2226), .B1_t (new_AGEMA_signal_2227), .B1_f (new_AGEMA_signal_2228), .Z0_t (SubCellInst_SboxInst_1_n15), .Z0_f (new_AGEMA_signal_2658), .Z1_t (new_AGEMA_signal_2659), .Z1_f (new_AGEMA_signal_2660) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_U17 ( .A0_t (Output_s0_t[48]), .A0_f (Output_s0_f[48]), .A1_t (Output_s1_t[48]), .A1_f (Output_s1_f[48]), .B0_t (SubCellInst_SboxInst_1_n11), .B0_f (new_AGEMA_signal_1217), .B1_t (new_AGEMA_signal_1218), .B1_f (new_AGEMA_signal_1219), .Z0_t (SubCellInst_SboxInst_1_n13), .Z0_f (new_AGEMA_signal_2226), .Z1_t (new_AGEMA_signal_2227), .Z1_f (new_AGEMA_signal_2228) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_U16 ( .A0_t (Output_s0_t[50]), .A0_f (Output_s0_f[50]), .A1_t (Output_s1_t[50]), .A1_f (Output_s1_f[50]), .B0_t (Output_s0_t[51]), .B0_f (Output_s0_f[51]), .B1_t (Output_s1_t[51]), .B1_f (Output_s1_f[51]), .Z0_t (SubCellInst_SboxInst_1_n11), .Z0_f (new_AGEMA_signal_1217), .Z1_t (new_AGEMA_signal_1218), .Z1_f (new_AGEMA_signal_1219) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U15 ( .A0_t (SubCellInst_SboxInst_1_n10), .A0_f (new_AGEMA_signal_2229), .A1_t (new_AGEMA_signal_2230), .A1_f (new_AGEMA_signal_2231), .B0_t (SubCellInst_SboxInst_1_n9), .B0_f (new_AGEMA_signal_1223), .B1_t (new_AGEMA_signal_1224), .B1_f (new_AGEMA_signal_1225), .Z0_t (Feedback[5]), .Z0_f (new_AGEMA_signal_2661), .Z1_t (new_AGEMA_signal_2662), .Z1_f (new_AGEMA_signal_2663) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U14 ( .A0_t (Output_s0_t[48]), .A0_f (Output_s0_f[48]), .A1_t (Output_s1_t[48]), .A1_f (Output_s1_f[48]), .B0_t (Output_s0_t[51]), .B0_f (Output_s0_f[51]), .B1_t (Output_s1_t[51]), .B1_f (Output_s1_f[51]), .Z0_t (SubCellInst_SboxInst_1_n9), .Z0_f (new_AGEMA_signal_1223), .Z1_t (new_AGEMA_signal_1224), .Z1_f (new_AGEMA_signal_1225) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U13 ( .A0_t (Output_s0_t[50]), .A0_f (Output_s0_f[50]), .A1_t (Output_s1_t[50]), .A1_f (Output_s1_f[50]), .B0_t (SubCellInst_SboxInst_1_n7), .B0_f (new_AGEMA_signal_1226), .B1_t (new_AGEMA_signal_1227), .B1_f (new_AGEMA_signal_1228), .Z0_t (SubCellInst_SboxInst_1_n10), .Z0_f (new_AGEMA_signal_2229), .Z1_t (new_AGEMA_signal_2230), .Z1_f (new_AGEMA_signal_2231) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U12 ( .A0_t (Output_s0_t[51]), .A0_f (Output_s0_f[51]), .A1_t (Output_s1_t[51]), .A1_f (Output_s1_f[51]), .B0_t (Output_s0_t[48]), .B0_f (Output_s0_f[48]), .B1_t (Output_s1_t[48]), .B1_f (Output_s1_f[48]), .Z0_t (SubCellInst_SboxInst_1_n7), .Z0_f (new_AGEMA_signal_1226), .Z1_t (new_AGEMA_signal_1227), .Z1_f (new_AGEMA_signal_1228) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U11 ( .A0_t (SubCellInst_SboxInst_1_n6), .A0_f (new_AGEMA_signal_2664), .A1_t (new_AGEMA_signal_2665), .A1_f (new_AGEMA_signal_2666), .B0_t (SubCellInst_SboxInst_1_n5), .B0_f (new_AGEMA_signal_1235), .B1_t (new_AGEMA_signal_1236), .B1_f (new_AGEMA_signal_1237), .Z0_t (Feedback[6]), .Z0_f (new_AGEMA_signal_3232), .Z1_t (new_AGEMA_signal_3233), .Z1_f (new_AGEMA_signal_3234) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U10 ( .A0_t (SubCellInst_SboxInst_1_n4), .A0_f (new_AGEMA_signal_2232), .A1_t (new_AGEMA_signal_2233), .A1_f (new_AGEMA_signal_2234), .B0_t (Output_s0_t[49]), .B0_f (Output_s0_f[49]), .B1_t (Output_s1_t[49]), .B1_f (Output_s1_f[49]), .Z0_t (SubCellInst_SboxInst_1_n6), .Z0_f (new_AGEMA_signal_2664), .Z1_t (new_AGEMA_signal_2665), .Z1_f (new_AGEMA_signal_2666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U9 ( .A0_t (SubCellInst_SboxInst_1_n3), .A0_f (new_AGEMA_signal_1229), .A1_t (new_AGEMA_signal_1230), .A1_f (new_AGEMA_signal_1231), .B0_t (Output_s0_t[50]), .B0_f (Output_s0_f[50]), .B1_t (Output_s1_t[50]), .B1_f (Output_s1_f[50]), .Z0_t (SubCellInst_SboxInst_1_n4), .Z0_f (new_AGEMA_signal_2232), .Z1_t (new_AGEMA_signal_2233), .Z1_f (new_AGEMA_signal_2234) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U8 ( .A0_t (Output_s0_t[48]), .A0_f (Output_s0_f[48]), .A1_t (Output_s1_t[48]), .A1_f (Output_s1_f[48]), .B0_t (Output_s0_t[51]), .B0_f (Output_s0_f[51]), .B1_t (Output_s1_t[51]), .B1_f (Output_s1_f[51]), .Z0_t (SubCellInst_SboxInst_1_n3), .Z0_f (new_AGEMA_signal_1229), .Z1_t (new_AGEMA_signal_1230), .Z1_f (new_AGEMA_signal_1231) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U7 ( .A0_t (SubCellInst_SboxInst_1_n5), .A0_f (new_AGEMA_signal_1235), .A1_t (new_AGEMA_signal_1236), .A1_f (new_AGEMA_signal_1237), .B0_t (SubCellInst_SboxInst_1_n1), .B0_f (new_AGEMA_signal_2238), .B1_t (new_AGEMA_signal_2239), .B1_f (new_AGEMA_signal_2240), .Z0_t (Feedback[7]), .Z0_f (new_AGEMA_signal_2667), .Z1_t (new_AGEMA_signal_2668), .Z1_f (new_AGEMA_signal_2669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U6 ( .A0_t (Output_s0_t[49]), .A0_f (Output_s0_f[49]), .A1_t (Output_s1_t[49]), .A1_f (Output_s1_f[49]), .B0_t (SubCellInst_SboxInst_1_n14), .B0_f (new_AGEMA_signal_1232), .B1_t (new_AGEMA_signal_1233), .B1_f (new_AGEMA_signal_1234), .Z0_t (SubCellInst_SboxInst_1_n1), .Z0_f (new_AGEMA_signal_2238), .Z1_t (new_AGEMA_signal_2239), .Z1_f (new_AGEMA_signal_2240) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_U5 ( .A0_t (Output_s0_t[50]), .A0_f (Output_s0_f[50]), .A1_t (Output_s1_t[50]), .A1_f (Output_s1_f[50]), .B0_t (Output_s0_t[51]), .B0_f (Output_s0_f[51]), .B1_t (Output_s1_t[51]), .B1_f (Output_s1_f[51]), .Z0_t (SubCellInst_SboxInst_1_n14), .Z0_f (new_AGEMA_signal_1232), .Z1_t (new_AGEMA_signal_1233), .Z1_f (new_AGEMA_signal_1234) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_U3 ( .A0_t (Output_s0_t[51]), .A0_f (Output_s0_f[51]), .A1_t (Output_s1_t[51]), .A1_f (Output_s1_f[51]), .B0_t (Output_s0_t[48]), .B0_f (Output_s0_f[48]), .B1_t (Output_s1_t[48]), .B1_f (Output_s1_f[48]), .Z0_t (SubCellInst_SboxInst_1_n5), .Z0_f (new_AGEMA_signal_1235), .Z1_t (new_AGEMA_signal_1236), .Z1_f (new_AGEMA_signal_1237) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_U19 ( .A0_t (SubCellInst_SboxInst_2_n15), .A0_f (new_AGEMA_signal_2670), .A1_t (new_AGEMA_signal_2671), .A1_f (new_AGEMA_signal_2672), .B0_t (SubCellInst_SboxInst_2_n14), .B0_f (new_AGEMA_signal_1259), .B1_t (new_AGEMA_signal_1260), .B1_f (new_AGEMA_signal_1261), .Z0_t (Feedback[8]), .Z0_f (new_AGEMA_signal_3235), .Z1_t (new_AGEMA_signal_3236), .Z1_f (new_AGEMA_signal_3237) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_U18 ( .A0_t (Output_s0_t[53]), .A0_f (Output_s0_f[53]), .A1_t (Output_s1_t[53]), .A1_f (Output_s1_f[53]), .B0_t (SubCellInst_SboxInst_2_n13), .B0_f (new_AGEMA_signal_2241), .B1_t (new_AGEMA_signal_2242), .B1_f (new_AGEMA_signal_2243), .Z0_t (SubCellInst_SboxInst_2_n15), .Z0_f (new_AGEMA_signal_2670), .Z1_t (new_AGEMA_signal_2671), .Z1_f (new_AGEMA_signal_2672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_U17 ( .A0_t (Output_s0_t[52]), .A0_f (Output_s0_f[52]), .A1_t (Output_s1_t[52]), .A1_f (Output_s1_f[52]), .B0_t (SubCellInst_SboxInst_2_n11), .B0_f (new_AGEMA_signal_1244), .B1_t (new_AGEMA_signal_1245), .B1_f (new_AGEMA_signal_1246), .Z0_t (SubCellInst_SboxInst_2_n13), .Z0_f (new_AGEMA_signal_2241), .Z1_t (new_AGEMA_signal_2242), .Z1_f (new_AGEMA_signal_2243) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_U16 ( .A0_t (Output_s0_t[54]), .A0_f (Output_s0_f[54]), .A1_t (Output_s1_t[54]), .A1_f (Output_s1_f[54]), .B0_t (Output_s0_t[55]), .B0_f (Output_s0_f[55]), .B1_t (Output_s1_t[55]), .B1_f (Output_s1_f[55]), .Z0_t (SubCellInst_SboxInst_2_n11), .Z0_f (new_AGEMA_signal_1244), .Z1_t (new_AGEMA_signal_1245), .Z1_f (new_AGEMA_signal_1246) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U15 ( .A0_t (SubCellInst_SboxInst_2_n10), .A0_f (new_AGEMA_signal_2244), .A1_t (new_AGEMA_signal_2245), .A1_f (new_AGEMA_signal_2246), .B0_t (SubCellInst_SboxInst_2_n9), .B0_f (new_AGEMA_signal_1250), .B1_t (new_AGEMA_signal_1251), .B1_f (new_AGEMA_signal_1252), .Z0_t (Feedback[9]), .Z0_f (new_AGEMA_signal_2673), .Z1_t (new_AGEMA_signal_2674), .Z1_f (new_AGEMA_signal_2675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U14 ( .A0_t (Output_s0_t[52]), .A0_f (Output_s0_f[52]), .A1_t (Output_s1_t[52]), .A1_f (Output_s1_f[52]), .B0_t (Output_s0_t[55]), .B0_f (Output_s0_f[55]), .B1_t (Output_s1_t[55]), .B1_f (Output_s1_f[55]), .Z0_t (SubCellInst_SboxInst_2_n9), .Z0_f (new_AGEMA_signal_1250), .Z1_t (new_AGEMA_signal_1251), .Z1_f (new_AGEMA_signal_1252) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U13 ( .A0_t (Output_s0_t[54]), .A0_f (Output_s0_f[54]), .A1_t (Output_s1_t[54]), .A1_f (Output_s1_f[54]), .B0_t (SubCellInst_SboxInst_2_n7), .B0_f (new_AGEMA_signal_1253), .B1_t (new_AGEMA_signal_1254), .B1_f (new_AGEMA_signal_1255), .Z0_t (SubCellInst_SboxInst_2_n10), .Z0_f (new_AGEMA_signal_2244), .Z1_t (new_AGEMA_signal_2245), .Z1_f (new_AGEMA_signal_2246) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U12 ( .A0_t (Output_s0_t[55]), .A0_f (Output_s0_f[55]), .A1_t (Output_s1_t[55]), .A1_f (Output_s1_f[55]), .B0_t (Output_s0_t[52]), .B0_f (Output_s0_f[52]), .B1_t (Output_s1_t[52]), .B1_f (Output_s1_f[52]), .Z0_t (SubCellInst_SboxInst_2_n7), .Z0_f (new_AGEMA_signal_1253), .Z1_t (new_AGEMA_signal_1254), .Z1_f (new_AGEMA_signal_1255) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U11 ( .A0_t (SubCellInst_SboxInst_2_n6), .A0_f (new_AGEMA_signal_2676), .A1_t (new_AGEMA_signal_2677), .A1_f (new_AGEMA_signal_2678), .B0_t (SubCellInst_SboxInst_2_n5), .B0_f (new_AGEMA_signal_1262), .B1_t (new_AGEMA_signal_1263), .B1_f (new_AGEMA_signal_1264), .Z0_t (Feedback[10]), .Z0_f (new_AGEMA_signal_3238), .Z1_t (new_AGEMA_signal_3239), .Z1_f (new_AGEMA_signal_3240) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U10 ( .A0_t (SubCellInst_SboxInst_2_n4), .A0_f (new_AGEMA_signal_2247), .A1_t (new_AGEMA_signal_2248), .A1_f (new_AGEMA_signal_2249), .B0_t (Output_s0_t[53]), .B0_f (Output_s0_f[53]), .B1_t (Output_s1_t[53]), .B1_f (Output_s1_f[53]), .Z0_t (SubCellInst_SboxInst_2_n6), .Z0_f (new_AGEMA_signal_2676), .Z1_t (new_AGEMA_signal_2677), .Z1_f (new_AGEMA_signal_2678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U9 ( .A0_t (SubCellInst_SboxInst_2_n3), .A0_f (new_AGEMA_signal_1256), .A1_t (new_AGEMA_signal_1257), .A1_f (new_AGEMA_signal_1258), .B0_t (Output_s0_t[54]), .B0_f (Output_s0_f[54]), .B1_t (Output_s1_t[54]), .B1_f (Output_s1_f[54]), .Z0_t (SubCellInst_SboxInst_2_n4), .Z0_f (new_AGEMA_signal_2247), .Z1_t (new_AGEMA_signal_2248), .Z1_f (new_AGEMA_signal_2249) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U8 ( .A0_t (Output_s0_t[52]), .A0_f (Output_s0_f[52]), .A1_t (Output_s1_t[52]), .A1_f (Output_s1_f[52]), .B0_t (Output_s0_t[55]), .B0_f (Output_s0_f[55]), .B1_t (Output_s1_t[55]), .B1_f (Output_s1_f[55]), .Z0_t (SubCellInst_SboxInst_2_n3), .Z0_f (new_AGEMA_signal_1256), .Z1_t (new_AGEMA_signal_1257), .Z1_f (new_AGEMA_signal_1258) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U7 ( .A0_t (SubCellInst_SboxInst_2_n5), .A0_f (new_AGEMA_signal_1262), .A1_t (new_AGEMA_signal_1263), .A1_f (new_AGEMA_signal_1264), .B0_t (SubCellInst_SboxInst_2_n1), .B0_f (new_AGEMA_signal_2253), .B1_t (new_AGEMA_signal_2254), .B1_f (new_AGEMA_signal_2255), .Z0_t (Feedback[11]), .Z0_f (new_AGEMA_signal_2679), .Z1_t (new_AGEMA_signal_2680), .Z1_f (new_AGEMA_signal_2681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U6 ( .A0_t (Output_s0_t[53]), .A0_f (Output_s0_f[53]), .A1_t (Output_s1_t[53]), .A1_f (Output_s1_f[53]), .B0_t (SubCellInst_SboxInst_2_n14), .B0_f (new_AGEMA_signal_1259), .B1_t (new_AGEMA_signal_1260), .B1_f (new_AGEMA_signal_1261), .Z0_t (SubCellInst_SboxInst_2_n1), .Z0_f (new_AGEMA_signal_2253), .Z1_t (new_AGEMA_signal_2254), .Z1_f (new_AGEMA_signal_2255) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_U5 ( .A0_t (Output_s0_t[54]), .A0_f (Output_s0_f[54]), .A1_t (Output_s1_t[54]), .A1_f (Output_s1_f[54]), .B0_t (Output_s0_t[55]), .B0_f (Output_s0_f[55]), .B1_t (Output_s1_t[55]), .B1_f (Output_s1_f[55]), .Z0_t (SubCellInst_SboxInst_2_n14), .Z0_f (new_AGEMA_signal_1259), .Z1_t (new_AGEMA_signal_1260), .Z1_f (new_AGEMA_signal_1261) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_U3 ( .A0_t (Output_s0_t[55]), .A0_f (Output_s0_f[55]), .A1_t (Output_s1_t[55]), .A1_f (Output_s1_f[55]), .B0_t (Output_s0_t[52]), .B0_f (Output_s0_f[52]), .B1_t (Output_s1_t[52]), .B1_f (Output_s1_f[52]), .Z0_t (SubCellInst_SboxInst_2_n5), .Z0_f (new_AGEMA_signal_1262), .Z1_t (new_AGEMA_signal_1263), .Z1_f (new_AGEMA_signal_1264) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_U19 ( .A0_t (SubCellInst_SboxInst_3_n15), .A0_f (new_AGEMA_signal_2682), .A1_t (new_AGEMA_signal_2683), .A1_f (new_AGEMA_signal_2684), .B0_t (SubCellInst_SboxInst_3_n14), .B0_f (new_AGEMA_signal_1286), .B1_t (new_AGEMA_signal_1287), .B1_f (new_AGEMA_signal_1288), .Z0_t (Feedback[12]), .Z0_f (new_AGEMA_signal_3241), .Z1_t (new_AGEMA_signal_3242), .Z1_f (new_AGEMA_signal_3243) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_U18 ( .A0_t (Output_s0_t[57]), .A0_f (Output_s0_f[57]), .A1_t (Output_s1_t[57]), .A1_f (Output_s1_f[57]), .B0_t (SubCellInst_SboxInst_3_n13), .B0_f (new_AGEMA_signal_2256), .B1_t (new_AGEMA_signal_2257), .B1_f (new_AGEMA_signal_2258), .Z0_t (SubCellInst_SboxInst_3_n15), .Z0_f (new_AGEMA_signal_2682), .Z1_t (new_AGEMA_signal_2683), .Z1_f (new_AGEMA_signal_2684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_U17 ( .A0_t (Output_s0_t[56]), .A0_f (Output_s0_f[56]), .A1_t (Output_s1_t[56]), .A1_f (Output_s1_f[56]), .B0_t (SubCellInst_SboxInst_3_n11), .B0_f (new_AGEMA_signal_1271), .B1_t (new_AGEMA_signal_1272), .B1_f (new_AGEMA_signal_1273), .Z0_t (SubCellInst_SboxInst_3_n13), .Z0_f (new_AGEMA_signal_2256), .Z1_t (new_AGEMA_signal_2257), .Z1_f (new_AGEMA_signal_2258) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_U16 ( .A0_t (Output_s0_t[58]), .A0_f (Output_s0_f[58]), .A1_t (Output_s1_t[58]), .A1_f (Output_s1_f[58]), .B0_t (Output_s0_t[59]), .B0_f (Output_s0_f[59]), .B1_t (Output_s1_t[59]), .B1_f (Output_s1_f[59]), .Z0_t (SubCellInst_SboxInst_3_n11), .Z0_f (new_AGEMA_signal_1271), .Z1_t (new_AGEMA_signal_1272), .Z1_f (new_AGEMA_signal_1273) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U15 ( .A0_t (SubCellInst_SboxInst_3_n10), .A0_f (new_AGEMA_signal_2259), .A1_t (new_AGEMA_signal_2260), .A1_f (new_AGEMA_signal_2261), .B0_t (SubCellInst_SboxInst_3_n9), .B0_f (new_AGEMA_signal_1277), .B1_t (new_AGEMA_signal_1278), .B1_f (new_AGEMA_signal_1279), .Z0_t (Feedback[13]), .Z0_f (new_AGEMA_signal_2685), .Z1_t (new_AGEMA_signal_2686), .Z1_f (new_AGEMA_signal_2687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U14 ( .A0_t (Output_s0_t[56]), .A0_f (Output_s0_f[56]), .A1_t (Output_s1_t[56]), .A1_f (Output_s1_f[56]), .B0_t (Output_s0_t[59]), .B0_f (Output_s0_f[59]), .B1_t (Output_s1_t[59]), .B1_f (Output_s1_f[59]), .Z0_t (SubCellInst_SboxInst_3_n9), .Z0_f (new_AGEMA_signal_1277), .Z1_t (new_AGEMA_signal_1278), .Z1_f (new_AGEMA_signal_1279) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U13 ( .A0_t (Output_s0_t[58]), .A0_f (Output_s0_f[58]), .A1_t (Output_s1_t[58]), .A1_f (Output_s1_f[58]), .B0_t (SubCellInst_SboxInst_3_n7), .B0_f (new_AGEMA_signal_1280), .B1_t (new_AGEMA_signal_1281), .B1_f (new_AGEMA_signal_1282), .Z0_t (SubCellInst_SboxInst_3_n10), .Z0_f (new_AGEMA_signal_2259), .Z1_t (new_AGEMA_signal_2260), .Z1_f (new_AGEMA_signal_2261) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U12 ( .A0_t (Output_s0_t[59]), .A0_f (Output_s0_f[59]), .A1_t (Output_s1_t[59]), .A1_f (Output_s1_f[59]), .B0_t (Output_s0_t[56]), .B0_f (Output_s0_f[56]), .B1_t (Output_s1_t[56]), .B1_f (Output_s1_f[56]), .Z0_t (SubCellInst_SboxInst_3_n7), .Z0_f (new_AGEMA_signal_1280), .Z1_t (new_AGEMA_signal_1281), .Z1_f (new_AGEMA_signal_1282) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U11 ( .A0_t (SubCellInst_SboxInst_3_n6), .A0_f (new_AGEMA_signal_2688), .A1_t (new_AGEMA_signal_2689), .A1_f (new_AGEMA_signal_2690), .B0_t (SubCellInst_SboxInst_3_n5), .B0_f (new_AGEMA_signal_1289), .B1_t (new_AGEMA_signal_1290), .B1_f (new_AGEMA_signal_1291), .Z0_t (Feedback[14]), .Z0_f (new_AGEMA_signal_3244), .Z1_t (new_AGEMA_signal_3245), .Z1_f (new_AGEMA_signal_3246) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U10 ( .A0_t (SubCellInst_SboxInst_3_n4), .A0_f (new_AGEMA_signal_2262), .A1_t (new_AGEMA_signal_2263), .A1_f (new_AGEMA_signal_2264), .B0_t (Output_s0_t[57]), .B0_f (Output_s0_f[57]), .B1_t (Output_s1_t[57]), .B1_f (Output_s1_f[57]), .Z0_t (SubCellInst_SboxInst_3_n6), .Z0_f (new_AGEMA_signal_2688), .Z1_t (new_AGEMA_signal_2689), .Z1_f (new_AGEMA_signal_2690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U9 ( .A0_t (SubCellInst_SboxInst_3_n3), .A0_f (new_AGEMA_signal_1283), .A1_t (new_AGEMA_signal_1284), .A1_f (new_AGEMA_signal_1285), .B0_t (Output_s0_t[58]), .B0_f (Output_s0_f[58]), .B1_t (Output_s1_t[58]), .B1_f (Output_s1_f[58]), .Z0_t (SubCellInst_SboxInst_3_n4), .Z0_f (new_AGEMA_signal_2262), .Z1_t (new_AGEMA_signal_2263), .Z1_f (new_AGEMA_signal_2264) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U8 ( .A0_t (Output_s0_t[56]), .A0_f (Output_s0_f[56]), .A1_t (Output_s1_t[56]), .A1_f (Output_s1_f[56]), .B0_t (Output_s0_t[59]), .B0_f (Output_s0_f[59]), .B1_t (Output_s1_t[59]), .B1_f (Output_s1_f[59]), .Z0_t (SubCellInst_SboxInst_3_n3), .Z0_f (new_AGEMA_signal_1283), .Z1_t (new_AGEMA_signal_1284), .Z1_f (new_AGEMA_signal_1285) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U7 ( .A0_t (SubCellInst_SboxInst_3_n5), .A0_f (new_AGEMA_signal_1289), .A1_t (new_AGEMA_signal_1290), .A1_f (new_AGEMA_signal_1291), .B0_t (SubCellInst_SboxInst_3_n1), .B0_f (new_AGEMA_signal_2268), .B1_t (new_AGEMA_signal_2269), .B1_f (new_AGEMA_signal_2270), .Z0_t (Feedback[15]), .Z0_f (new_AGEMA_signal_2691), .Z1_t (new_AGEMA_signal_2692), .Z1_f (new_AGEMA_signal_2693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U6 ( .A0_t (Output_s0_t[57]), .A0_f (Output_s0_f[57]), .A1_t (Output_s1_t[57]), .A1_f (Output_s1_f[57]), .B0_t (SubCellInst_SboxInst_3_n14), .B0_f (new_AGEMA_signal_1286), .B1_t (new_AGEMA_signal_1287), .B1_f (new_AGEMA_signal_1288), .Z0_t (SubCellInst_SboxInst_3_n1), .Z0_f (new_AGEMA_signal_2268), .Z1_t (new_AGEMA_signal_2269), .Z1_f (new_AGEMA_signal_2270) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_U5 ( .A0_t (Output_s0_t[58]), .A0_f (Output_s0_f[58]), .A1_t (Output_s1_t[58]), .A1_f (Output_s1_f[58]), .B0_t (Output_s0_t[59]), .B0_f (Output_s0_f[59]), .B1_t (Output_s1_t[59]), .B1_f (Output_s1_f[59]), .Z0_t (SubCellInst_SboxInst_3_n14), .Z0_f (new_AGEMA_signal_1286), .Z1_t (new_AGEMA_signal_1287), .Z1_f (new_AGEMA_signal_1288) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_U3 ( .A0_t (Output_s0_t[59]), .A0_f (Output_s0_f[59]), .A1_t (Output_s1_t[59]), .A1_f (Output_s1_f[59]), .B0_t (Output_s0_t[56]), .B0_f (Output_s0_f[56]), .B1_t (Output_s1_t[56]), .B1_f (Output_s1_f[56]), .Z0_t (SubCellInst_SboxInst_3_n5), .Z0_f (new_AGEMA_signal_1289), .Z1_t (new_AGEMA_signal_1290), .Z1_f (new_AGEMA_signal_1291) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U19 ( .A0_t (SubCellInst_SboxInst_4_n15), .A0_f (new_AGEMA_signal_1301), .A1_t (new_AGEMA_signal_1302), .A1_f (new_AGEMA_signal_1303), .B0_t (SubCellInst_SboxInst_4_n14), .B0_f (new_AGEMA_signal_2271), .B1_t (new_AGEMA_signal_2272), .B1_f (new_AGEMA_signal_2273), .Z0_t (Feedback[17]), .Z0_f (new_AGEMA_signal_2694), .Z1_t (new_AGEMA_signal_2695), .Z1_f (new_AGEMA_signal_2696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U18 ( .A0_t (Output_s0_t[34]), .A0_f (Output_s0_f[34]), .A1_t (Output_s1_t[34]), .A1_f (Output_s1_f[34]), .B0_t (SubCellInst_SboxInst_4_n13), .B0_f (new_AGEMA_signal_1298), .B1_t (new_AGEMA_signal_1299), .B1_f (new_AGEMA_signal_1300), .Z0_t (SubCellInst_SboxInst_4_n14), .Z0_f (new_AGEMA_signal_2271), .Z1_t (new_AGEMA_signal_2272), .Z1_f (new_AGEMA_signal_2273) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U17 ( .A0_t (Output_s0_t[35]), .A0_f (Output_s0_f[35]), .A1_t (Output_s1_t[35]), .A1_f (Output_s1_f[35]), .B0_t (Output_s0_t[32]), .B0_f (Output_s0_f[32]), .B1_t (Output_s1_t[32]), .B1_f (Output_s1_f[32]), .Z0_t (SubCellInst_SboxInst_4_n13), .Z0_f (new_AGEMA_signal_1298), .Z1_t (new_AGEMA_signal_1299), .Z1_f (new_AGEMA_signal_1300) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U16 ( .A0_t (Output_s0_t[32]), .A0_f (Output_s0_f[32]), .A1_t (Output_s1_t[32]), .A1_f (Output_s1_f[32]), .B0_t (Output_s0_t[35]), .B0_f (Output_s0_f[35]), .B1_t (Output_s1_t[35]), .B1_f (Output_s1_f[35]), .Z0_t (SubCellInst_SboxInst_4_n15), .Z0_f (new_AGEMA_signal_1301), .Z1_t (new_AGEMA_signal_1302), .Z1_f (new_AGEMA_signal_1303) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U15 ( .A0_t (SubCellInst_SboxInst_4_n10), .A0_f (new_AGEMA_signal_1316), .A1_t (new_AGEMA_signal_1317), .A1_f (new_AGEMA_signal_1318), .B0_t (SubCellInst_SboxInst_4_n9), .B0_f (new_AGEMA_signal_2277), .B1_t (new_AGEMA_signal_2278), .B1_f (new_AGEMA_signal_2279), .Z0_t (Feedback[19]), .Z0_f (new_AGEMA_signal_2697), .Z1_t (new_AGEMA_signal_2698), .Z1_f (new_AGEMA_signal_2699) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U14 ( .A0_t (Output_s0_t[33]), .A0_f (Output_s0_f[33]), .A1_t (Output_s1_t[33]), .A1_f (Output_s1_f[33]), .B0_t (SubCellInst_SboxInst_4_n8), .B0_f (new_AGEMA_signal_1310), .B1_t (new_AGEMA_signal_1311), .B1_f (new_AGEMA_signal_1312), .Z0_t (SubCellInst_SboxInst_4_n9), .Z0_f (new_AGEMA_signal_2277), .Z1_t (new_AGEMA_signal_2278), .Z1_f (new_AGEMA_signal_2279) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_U13 ( .A0_t (SubCellInst_SboxInst_4_n8), .A0_f (new_AGEMA_signal_1310), .A1_t (new_AGEMA_signal_1311), .A1_f (new_AGEMA_signal_1312), .B0_t (SubCellInst_SboxInst_4_n7), .B0_f (new_AGEMA_signal_2700), .B1_t (new_AGEMA_signal_2701), .B1_f (new_AGEMA_signal_2702), .Z0_t (Feedback[16]), .Z0_f (new_AGEMA_signal_3247), .Z1_t (new_AGEMA_signal_3248), .Z1_f (new_AGEMA_signal_3249) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_U12 ( .A0_t (Output_s0_t[33]), .A0_f (Output_s0_f[33]), .A1_t (Output_s1_t[33]), .A1_f (Output_s1_f[33]), .B0_t (SubCellInst_SboxInst_4_n6), .B0_f (new_AGEMA_signal_2280), .B1_t (new_AGEMA_signal_2281), .B1_f (new_AGEMA_signal_2282), .Z0_t (SubCellInst_SboxInst_4_n7), .Z0_f (new_AGEMA_signal_2700), .Z1_t (new_AGEMA_signal_2701), .Z1_f (new_AGEMA_signal_2702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_U11 ( .A0_t (Output_s0_t[32]), .A0_f (Output_s0_f[32]), .A1_t (Output_s1_t[32]), .A1_f (Output_s1_f[32]), .B0_t (SubCellInst_SboxInst_4_n5), .B0_f (new_AGEMA_signal_1307), .B1_t (new_AGEMA_signal_1308), .B1_f (new_AGEMA_signal_1309), .Z0_t (SubCellInst_SboxInst_4_n6), .Z0_f (new_AGEMA_signal_2280), .Z1_t (new_AGEMA_signal_2281), .Z1_f (new_AGEMA_signal_2282) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_U10 ( .A0_t (Output_s0_t[35]), .A0_f (Output_s0_f[35]), .A1_t (Output_s1_t[35]), .A1_f (Output_s1_f[35]), .B0_t (Output_s0_t[34]), .B0_f (Output_s0_f[34]), .B1_t (Output_s1_t[34]), .B1_f (Output_s1_f[34]), .Z0_t (SubCellInst_SboxInst_4_n5), .Z0_f (new_AGEMA_signal_1307), .Z1_t (new_AGEMA_signal_1308), .Z1_f (new_AGEMA_signal_1309) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_U9 ( .A0_t (Output_s0_t[35]), .A0_f (Output_s0_f[35]), .A1_t (Output_s1_t[35]), .A1_f (Output_s1_f[35]), .B0_t (Output_s0_t[34]), .B0_f (Output_s0_f[34]), .B1_t (Output_s1_t[34]), .B1_f (Output_s1_f[34]), .Z0_t (SubCellInst_SboxInst_4_n8), .Z0_f (new_AGEMA_signal_1310), .Z1_t (new_AGEMA_signal_1311), .Z1_f (new_AGEMA_signal_1312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U8 ( .A0_t (SubCellInst_SboxInst_4_n10), .A0_f (new_AGEMA_signal_1316), .A1_t (new_AGEMA_signal_1317), .A1_f (new_AGEMA_signal_1318), .B0_t (SubCellInst_SboxInst_4_n3), .B0_f (new_AGEMA_signal_2703), .B1_t (new_AGEMA_signal_2704), .B1_f (new_AGEMA_signal_2705), .Z0_t (Feedback[18]), .Z0_f (new_AGEMA_signal_3250), .Z1_t (new_AGEMA_signal_3251), .Z1_f (new_AGEMA_signal_3252) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U7 ( .A0_t (SubCellInst_SboxInst_4_n2), .A0_f (new_AGEMA_signal_2283), .A1_t (new_AGEMA_signal_2284), .A1_f (new_AGEMA_signal_2285), .B0_t (Output_s0_t[33]), .B0_f (Output_s0_f[33]), .B1_t (Output_s1_t[33]), .B1_f (Output_s1_f[33]), .Z0_t (SubCellInst_SboxInst_4_n3), .Z0_f (new_AGEMA_signal_2703), .Z1_t (new_AGEMA_signal_2704), .Z1_f (new_AGEMA_signal_2705) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U6 ( .A0_t (SubCellInst_SboxInst_4_n1), .A0_f (new_AGEMA_signal_1313), .A1_t (new_AGEMA_signal_1314), .A1_f (new_AGEMA_signal_1315), .B0_t (Output_s0_t[34]), .B0_f (Output_s0_f[34]), .B1_t (Output_s1_t[34]), .B1_f (Output_s1_f[34]), .Z0_t (SubCellInst_SboxInst_4_n2), .Z0_f (new_AGEMA_signal_2283), .Z1_t (new_AGEMA_signal_2284), .Z1_f (new_AGEMA_signal_2285) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U4 ( .A0_t (Output_s0_t[35]), .A0_f (Output_s0_f[35]), .A1_t (Output_s1_t[35]), .A1_f (Output_s1_f[35]), .B0_t (Output_s0_t[32]), .B0_f (Output_s0_f[32]), .B1_t (Output_s1_t[32]), .B1_f (Output_s1_f[32]), .Z0_t (SubCellInst_SboxInst_4_n1), .Z0_f (new_AGEMA_signal_1313), .Z1_t (new_AGEMA_signal_1314), .Z1_f (new_AGEMA_signal_1315) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_U3 ( .A0_t (Output_s0_t[32]), .A0_f (Output_s0_f[32]), .A1_t (Output_s1_t[32]), .A1_f (Output_s1_f[32]), .B0_t (Output_s0_t[35]), .B0_f (Output_s0_f[35]), .B1_t (Output_s1_t[35]), .B1_f (Output_s1_f[35]), .Z0_t (SubCellInst_SboxInst_4_n10), .Z0_f (new_AGEMA_signal_1316), .Z1_t (new_AGEMA_signal_1317), .Z1_f (new_AGEMA_signal_1318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U19 ( .A0_t (SubCellInst_SboxInst_5_n15), .A0_f (new_AGEMA_signal_1328), .A1_t (new_AGEMA_signal_1329), .A1_f (new_AGEMA_signal_1330), .B0_t (SubCellInst_SboxInst_5_n14), .B0_f (new_AGEMA_signal_2286), .B1_t (new_AGEMA_signal_2287), .B1_f (new_AGEMA_signal_2288), .Z0_t (Feedback[21]), .Z0_f (new_AGEMA_signal_2706), .Z1_t (new_AGEMA_signal_2707), .Z1_f (new_AGEMA_signal_2708) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U18 ( .A0_t (Output_s0_t[46]), .A0_f (Output_s0_f[46]), .A1_t (Output_s1_t[46]), .A1_f (Output_s1_f[46]), .B0_t (SubCellInst_SboxInst_5_n13), .B0_f (new_AGEMA_signal_1325), .B1_t (new_AGEMA_signal_1326), .B1_f (new_AGEMA_signal_1327), .Z0_t (SubCellInst_SboxInst_5_n14), .Z0_f (new_AGEMA_signal_2286), .Z1_t (new_AGEMA_signal_2287), .Z1_f (new_AGEMA_signal_2288) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U17 ( .A0_t (Output_s0_t[47]), .A0_f (Output_s0_f[47]), .A1_t (Output_s1_t[47]), .A1_f (Output_s1_f[47]), .B0_t (Output_s0_t[44]), .B0_f (Output_s0_f[44]), .B1_t (Output_s1_t[44]), .B1_f (Output_s1_f[44]), .Z0_t (SubCellInst_SboxInst_5_n13), .Z0_f (new_AGEMA_signal_1325), .Z1_t (new_AGEMA_signal_1326), .Z1_f (new_AGEMA_signal_1327) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U16 ( .A0_t (Output_s0_t[44]), .A0_f (Output_s0_f[44]), .A1_t (Output_s1_t[44]), .A1_f (Output_s1_f[44]), .B0_t (Output_s0_t[47]), .B0_f (Output_s0_f[47]), .B1_t (Output_s1_t[47]), .B1_f (Output_s1_f[47]), .Z0_t (SubCellInst_SboxInst_5_n15), .Z0_f (new_AGEMA_signal_1328), .Z1_t (new_AGEMA_signal_1329), .Z1_f (new_AGEMA_signal_1330) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U15 ( .A0_t (SubCellInst_SboxInst_5_n10), .A0_f (new_AGEMA_signal_1343), .A1_t (new_AGEMA_signal_1344), .A1_f (new_AGEMA_signal_1345), .B0_t (SubCellInst_SboxInst_5_n9), .B0_f (new_AGEMA_signal_2292), .B1_t (new_AGEMA_signal_2293), .B1_f (new_AGEMA_signal_2294), .Z0_t (Feedback[23]), .Z0_f (new_AGEMA_signal_2709), .Z1_t (new_AGEMA_signal_2710), .Z1_f (new_AGEMA_signal_2711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U14 ( .A0_t (Output_s0_t[45]), .A0_f (Output_s0_f[45]), .A1_t (Output_s1_t[45]), .A1_f (Output_s1_f[45]), .B0_t (SubCellInst_SboxInst_5_n8), .B0_f (new_AGEMA_signal_1337), .B1_t (new_AGEMA_signal_1338), .B1_f (new_AGEMA_signal_1339), .Z0_t (SubCellInst_SboxInst_5_n9), .Z0_f (new_AGEMA_signal_2292), .Z1_t (new_AGEMA_signal_2293), .Z1_f (new_AGEMA_signal_2294) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_U13 ( .A0_t (SubCellInst_SboxInst_5_n8), .A0_f (new_AGEMA_signal_1337), .A1_t (new_AGEMA_signal_1338), .A1_f (new_AGEMA_signal_1339), .B0_t (SubCellInst_SboxInst_5_n7), .B0_f (new_AGEMA_signal_2712), .B1_t (new_AGEMA_signal_2713), .B1_f (new_AGEMA_signal_2714), .Z0_t (Feedback[20]), .Z0_f (new_AGEMA_signal_3253), .Z1_t (new_AGEMA_signal_3254), .Z1_f (new_AGEMA_signal_3255) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_U12 ( .A0_t (Output_s0_t[45]), .A0_f (Output_s0_f[45]), .A1_t (Output_s1_t[45]), .A1_f (Output_s1_f[45]), .B0_t (SubCellInst_SboxInst_5_n6), .B0_f (new_AGEMA_signal_2295), .B1_t (new_AGEMA_signal_2296), .B1_f (new_AGEMA_signal_2297), .Z0_t (SubCellInst_SboxInst_5_n7), .Z0_f (new_AGEMA_signal_2712), .Z1_t (new_AGEMA_signal_2713), .Z1_f (new_AGEMA_signal_2714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_U11 ( .A0_t (Output_s0_t[44]), .A0_f (Output_s0_f[44]), .A1_t (Output_s1_t[44]), .A1_f (Output_s1_f[44]), .B0_t (SubCellInst_SboxInst_5_n5), .B0_f (new_AGEMA_signal_1334), .B1_t (new_AGEMA_signal_1335), .B1_f (new_AGEMA_signal_1336), .Z0_t (SubCellInst_SboxInst_5_n6), .Z0_f (new_AGEMA_signal_2295), .Z1_t (new_AGEMA_signal_2296), .Z1_f (new_AGEMA_signal_2297) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_U10 ( .A0_t (Output_s0_t[47]), .A0_f (Output_s0_f[47]), .A1_t (Output_s1_t[47]), .A1_f (Output_s1_f[47]), .B0_t (Output_s0_t[46]), .B0_f (Output_s0_f[46]), .B1_t (Output_s1_t[46]), .B1_f (Output_s1_f[46]), .Z0_t (SubCellInst_SboxInst_5_n5), .Z0_f (new_AGEMA_signal_1334), .Z1_t (new_AGEMA_signal_1335), .Z1_f (new_AGEMA_signal_1336) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_U9 ( .A0_t (Output_s0_t[47]), .A0_f (Output_s0_f[47]), .A1_t (Output_s1_t[47]), .A1_f (Output_s1_f[47]), .B0_t (Output_s0_t[46]), .B0_f (Output_s0_f[46]), .B1_t (Output_s1_t[46]), .B1_f (Output_s1_f[46]), .Z0_t (SubCellInst_SboxInst_5_n8), .Z0_f (new_AGEMA_signal_1337), .Z1_t (new_AGEMA_signal_1338), .Z1_f (new_AGEMA_signal_1339) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U8 ( .A0_t (SubCellInst_SboxInst_5_n10), .A0_f (new_AGEMA_signal_1343), .A1_t (new_AGEMA_signal_1344), .A1_f (new_AGEMA_signal_1345), .B0_t (SubCellInst_SboxInst_5_n3), .B0_f (new_AGEMA_signal_2715), .B1_t (new_AGEMA_signal_2716), .B1_f (new_AGEMA_signal_2717), .Z0_t (Feedback[22]), .Z0_f (new_AGEMA_signal_3256), .Z1_t (new_AGEMA_signal_3257), .Z1_f (new_AGEMA_signal_3258) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U7 ( .A0_t (SubCellInst_SboxInst_5_n2), .A0_f (new_AGEMA_signal_2298), .A1_t (new_AGEMA_signal_2299), .A1_f (new_AGEMA_signal_2300), .B0_t (Output_s0_t[45]), .B0_f (Output_s0_f[45]), .B1_t (Output_s1_t[45]), .B1_f (Output_s1_f[45]), .Z0_t (SubCellInst_SboxInst_5_n3), .Z0_f (new_AGEMA_signal_2715), .Z1_t (new_AGEMA_signal_2716), .Z1_f (new_AGEMA_signal_2717) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U6 ( .A0_t (SubCellInst_SboxInst_5_n1), .A0_f (new_AGEMA_signal_1340), .A1_t (new_AGEMA_signal_1341), .A1_f (new_AGEMA_signal_1342), .B0_t (Output_s0_t[46]), .B0_f (Output_s0_f[46]), .B1_t (Output_s1_t[46]), .B1_f (Output_s1_f[46]), .Z0_t (SubCellInst_SboxInst_5_n2), .Z0_f (new_AGEMA_signal_2298), .Z1_t (new_AGEMA_signal_2299), .Z1_f (new_AGEMA_signal_2300) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U4 ( .A0_t (Output_s0_t[47]), .A0_f (Output_s0_f[47]), .A1_t (Output_s1_t[47]), .A1_f (Output_s1_f[47]), .B0_t (Output_s0_t[44]), .B0_f (Output_s0_f[44]), .B1_t (Output_s1_t[44]), .B1_f (Output_s1_f[44]), .Z0_t (SubCellInst_SboxInst_5_n1), .Z0_f (new_AGEMA_signal_1340), .Z1_t (new_AGEMA_signal_1341), .Z1_f (new_AGEMA_signal_1342) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_U3 ( .A0_t (Output_s0_t[44]), .A0_f (Output_s0_f[44]), .A1_t (Output_s1_t[44]), .A1_f (Output_s1_f[44]), .B0_t (Output_s0_t[47]), .B0_f (Output_s0_f[47]), .B1_t (Output_s1_t[47]), .B1_f (Output_s1_f[47]), .Z0_t (SubCellInst_SboxInst_5_n10), .Z0_f (new_AGEMA_signal_1343), .Z1_t (new_AGEMA_signal_1344), .Z1_f (new_AGEMA_signal_1345) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U19 ( .A0_t (SubCellInst_SboxInst_6_n15), .A0_f (new_AGEMA_signal_1355), .A1_t (new_AGEMA_signal_1356), .A1_f (new_AGEMA_signal_1357), .B0_t (SubCellInst_SboxInst_6_n14), .B0_f (new_AGEMA_signal_2301), .B1_t (new_AGEMA_signal_2302), .B1_f (new_AGEMA_signal_2303), .Z0_t (Feedback[25]), .Z0_f (new_AGEMA_signal_2718), .Z1_t (new_AGEMA_signal_2719), .Z1_f (new_AGEMA_signal_2720) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U18 ( .A0_t (Output_s0_t[42]), .A0_f (Output_s0_f[42]), .A1_t (Output_s1_t[42]), .A1_f (Output_s1_f[42]), .B0_t (SubCellInst_SboxInst_6_n13), .B0_f (new_AGEMA_signal_1352), .B1_t (new_AGEMA_signal_1353), .B1_f (new_AGEMA_signal_1354), .Z0_t (SubCellInst_SboxInst_6_n14), .Z0_f (new_AGEMA_signal_2301), .Z1_t (new_AGEMA_signal_2302), .Z1_f (new_AGEMA_signal_2303) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U17 ( .A0_t (Output_s0_t[43]), .A0_f (Output_s0_f[43]), .A1_t (Output_s1_t[43]), .A1_f (Output_s1_f[43]), .B0_t (Output_s0_t[40]), .B0_f (Output_s0_f[40]), .B1_t (Output_s1_t[40]), .B1_f (Output_s1_f[40]), .Z0_t (SubCellInst_SboxInst_6_n13), .Z0_f (new_AGEMA_signal_1352), .Z1_t (new_AGEMA_signal_1353), .Z1_f (new_AGEMA_signal_1354) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U16 ( .A0_t (Output_s0_t[40]), .A0_f (Output_s0_f[40]), .A1_t (Output_s1_t[40]), .A1_f (Output_s1_f[40]), .B0_t (Output_s0_t[43]), .B0_f (Output_s0_f[43]), .B1_t (Output_s1_t[43]), .B1_f (Output_s1_f[43]), .Z0_t (SubCellInst_SboxInst_6_n15), .Z0_f (new_AGEMA_signal_1355), .Z1_t (new_AGEMA_signal_1356), .Z1_f (new_AGEMA_signal_1357) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U15 ( .A0_t (SubCellInst_SboxInst_6_n10), .A0_f (new_AGEMA_signal_1370), .A1_t (new_AGEMA_signal_1371), .A1_f (new_AGEMA_signal_1372), .B0_t (SubCellInst_SboxInst_6_n9), .B0_f (new_AGEMA_signal_2307), .B1_t (new_AGEMA_signal_2308), .B1_f (new_AGEMA_signal_2309), .Z0_t (Feedback[27]), .Z0_f (new_AGEMA_signal_2721), .Z1_t (new_AGEMA_signal_2722), .Z1_f (new_AGEMA_signal_2723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U14 ( .A0_t (Output_s0_t[41]), .A0_f (Output_s0_f[41]), .A1_t (Output_s1_t[41]), .A1_f (Output_s1_f[41]), .B0_t (SubCellInst_SboxInst_6_n8), .B0_f (new_AGEMA_signal_1364), .B1_t (new_AGEMA_signal_1365), .B1_f (new_AGEMA_signal_1366), .Z0_t (SubCellInst_SboxInst_6_n9), .Z0_f (new_AGEMA_signal_2307), .Z1_t (new_AGEMA_signal_2308), .Z1_f (new_AGEMA_signal_2309) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_U13 ( .A0_t (SubCellInst_SboxInst_6_n8), .A0_f (new_AGEMA_signal_1364), .A1_t (new_AGEMA_signal_1365), .A1_f (new_AGEMA_signal_1366), .B0_t (SubCellInst_SboxInst_6_n7), .B0_f (new_AGEMA_signal_2724), .B1_t (new_AGEMA_signal_2725), .B1_f (new_AGEMA_signal_2726), .Z0_t (Feedback[24]), .Z0_f (new_AGEMA_signal_3259), .Z1_t (new_AGEMA_signal_3260), .Z1_f (new_AGEMA_signal_3261) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_U12 ( .A0_t (Output_s0_t[41]), .A0_f (Output_s0_f[41]), .A1_t (Output_s1_t[41]), .A1_f (Output_s1_f[41]), .B0_t (SubCellInst_SboxInst_6_n6), .B0_f (new_AGEMA_signal_2310), .B1_t (new_AGEMA_signal_2311), .B1_f (new_AGEMA_signal_2312), .Z0_t (SubCellInst_SboxInst_6_n7), .Z0_f (new_AGEMA_signal_2724), .Z1_t (new_AGEMA_signal_2725), .Z1_f (new_AGEMA_signal_2726) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_U11 ( .A0_t (Output_s0_t[40]), .A0_f (Output_s0_f[40]), .A1_t (Output_s1_t[40]), .A1_f (Output_s1_f[40]), .B0_t (SubCellInst_SboxInst_6_n5), .B0_f (new_AGEMA_signal_1361), .B1_t (new_AGEMA_signal_1362), .B1_f (new_AGEMA_signal_1363), .Z0_t (SubCellInst_SboxInst_6_n6), .Z0_f (new_AGEMA_signal_2310), .Z1_t (new_AGEMA_signal_2311), .Z1_f (new_AGEMA_signal_2312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_U10 ( .A0_t (Output_s0_t[43]), .A0_f (Output_s0_f[43]), .A1_t (Output_s1_t[43]), .A1_f (Output_s1_f[43]), .B0_t (Output_s0_t[42]), .B0_f (Output_s0_f[42]), .B1_t (Output_s1_t[42]), .B1_f (Output_s1_f[42]), .Z0_t (SubCellInst_SboxInst_6_n5), .Z0_f (new_AGEMA_signal_1361), .Z1_t (new_AGEMA_signal_1362), .Z1_f (new_AGEMA_signal_1363) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_U9 ( .A0_t (Output_s0_t[43]), .A0_f (Output_s0_f[43]), .A1_t (Output_s1_t[43]), .A1_f (Output_s1_f[43]), .B0_t (Output_s0_t[42]), .B0_f (Output_s0_f[42]), .B1_t (Output_s1_t[42]), .B1_f (Output_s1_f[42]), .Z0_t (SubCellInst_SboxInst_6_n8), .Z0_f (new_AGEMA_signal_1364), .Z1_t (new_AGEMA_signal_1365), .Z1_f (new_AGEMA_signal_1366) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U8 ( .A0_t (SubCellInst_SboxInst_6_n10), .A0_f (new_AGEMA_signal_1370), .A1_t (new_AGEMA_signal_1371), .A1_f (new_AGEMA_signal_1372), .B0_t (SubCellInst_SboxInst_6_n3), .B0_f (new_AGEMA_signal_2727), .B1_t (new_AGEMA_signal_2728), .B1_f (new_AGEMA_signal_2729), .Z0_t (Feedback[26]), .Z0_f (new_AGEMA_signal_3262), .Z1_t (new_AGEMA_signal_3263), .Z1_f (new_AGEMA_signal_3264) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U7 ( .A0_t (SubCellInst_SboxInst_6_n2), .A0_f (new_AGEMA_signal_2313), .A1_t (new_AGEMA_signal_2314), .A1_f (new_AGEMA_signal_2315), .B0_t (Output_s0_t[41]), .B0_f (Output_s0_f[41]), .B1_t (Output_s1_t[41]), .B1_f (Output_s1_f[41]), .Z0_t (SubCellInst_SboxInst_6_n3), .Z0_f (new_AGEMA_signal_2727), .Z1_t (new_AGEMA_signal_2728), .Z1_f (new_AGEMA_signal_2729) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U6 ( .A0_t (SubCellInst_SboxInst_6_n1), .A0_f (new_AGEMA_signal_1367), .A1_t (new_AGEMA_signal_1368), .A1_f (new_AGEMA_signal_1369), .B0_t (Output_s0_t[42]), .B0_f (Output_s0_f[42]), .B1_t (Output_s1_t[42]), .B1_f (Output_s1_f[42]), .Z0_t (SubCellInst_SboxInst_6_n2), .Z0_f (new_AGEMA_signal_2313), .Z1_t (new_AGEMA_signal_2314), .Z1_f (new_AGEMA_signal_2315) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U4 ( .A0_t (Output_s0_t[43]), .A0_f (Output_s0_f[43]), .A1_t (Output_s1_t[43]), .A1_f (Output_s1_f[43]), .B0_t (Output_s0_t[40]), .B0_f (Output_s0_f[40]), .B1_t (Output_s1_t[40]), .B1_f (Output_s1_f[40]), .Z0_t (SubCellInst_SboxInst_6_n1), .Z0_f (new_AGEMA_signal_1367), .Z1_t (new_AGEMA_signal_1368), .Z1_f (new_AGEMA_signal_1369) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_U3 ( .A0_t (Output_s0_t[40]), .A0_f (Output_s0_f[40]), .A1_t (Output_s1_t[40]), .A1_f (Output_s1_f[40]), .B0_t (Output_s0_t[43]), .B0_f (Output_s0_f[43]), .B1_t (Output_s1_t[43]), .B1_f (Output_s1_f[43]), .Z0_t (SubCellInst_SboxInst_6_n10), .Z0_f (new_AGEMA_signal_1370), .Z1_t (new_AGEMA_signal_1371), .Z1_f (new_AGEMA_signal_1372) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U19 ( .A0_t (SubCellInst_SboxInst_7_n15), .A0_f (new_AGEMA_signal_1382), .A1_t (new_AGEMA_signal_1383), .A1_f (new_AGEMA_signal_1384), .B0_t (SubCellInst_SboxInst_7_n14), .B0_f (new_AGEMA_signal_2316), .B1_t (new_AGEMA_signal_2317), .B1_f (new_AGEMA_signal_2318), .Z0_t (Feedback[29]), .Z0_f (new_AGEMA_signal_2730), .Z1_t (new_AGEMA_signal_2731), .Z1_f (new_AGEMA_signal_2732) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U18 ( .A0_t (Output_s0_t[38]), .A0_f (Output_s0_f[38]), .A1_t (Output_s1_t[38]), .A1_f (Output_s1_f[38]), .B0_t (SubCellInst_SboxInst_7_n13), .B0_f (new_AGEMA_signal_1379), .B1_t (new_AGEMA_signal_1380), .B1_f (new_AGEMA_signal_1381), .Z0_t (SubCellInst_SboxInst_7_n14), .Z0_f (new_AGEMA_signal_2316), .Z1_t (new_AGEMA_signal_2317), .Z1_f (new_AGEMA_signal_2318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U17 ( .A0_t (Output_s0_t[39]), .A0_f (Output_s0_f[39]), .A1_t (Output_s1_t[39]), .A1_f (Output_s1_f[39]), .B0_t (Output_s0_t[36]), .B0_f (Output_s0_f[36]), .B1_t (Output_s1_t[36]), .B1_f (Output_s1_f[36]), .Z0_t (SubCellInst_SboxInst_7_n13), .Z0_f (new_AGEMA_signal_1379), .Z1_t (new_AGEMA_signal_1380), .Z1_f (new_AGEMA_signal_1381) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U16 ( .A0_t (Output_s0_t[36]), .A0_f (Output_s0_f[36]), .A1_t (Output_s1_t[36]), .A1_f (Output_s1_f[36]), .B0_t (Output_s0_t[39]), .B0_f (Output_s0_f[39]), .B1_t (Output_s1_t[39]), .B1_f (Output_s1_f[39]), .Z0_t (SubCellInst_SboxInst_7_n15), .Z0_f (new_AGEMA_signal_1382), .Z1_t (new_AGEMA_signal_1383), .Z1_f (new_AGEMA_signal_1384) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U15 ( .A0_t (SubCellInst_SboxInst_7_n10), .A0_f (new_AGEMA_signal_1397), .A1_t (new_AGEMA_signal_1398), .A1_f (new_AGEMA_signal_1399), .B0_t (SubCellInst_SboxInst_7_n9), .B0_f (new_AGEMA_signal_2322), .B1_t (new_AGEMA_signal_2323), .B1_f (new_AGEMA_signal_2324), .Z0_t (Feedback[31]), .Z0_f (new_AGEMA_signal_2733), .Z1_t (new_AGEMA_signal_2734), .Z1_f (new_AGEMA_signal_2735) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U14 ( .A0_t (Output_s0_t[37]), .A0_f (Output_s0_f[37]), .A1_t (Output_s1_t[37]), .A1_f (Output_s1_f[37]), .B0_t (SubCellInst_SboxInst_7_n8), .B0_f (new_AGEMA_signal_1391), .B1_t (new_AGEMA_signal_1392), .B1_f (new_AGEMA_signal_1393), .Z0_t (SubCellInst_SboxInst_7_n9), .Z0_f (new_AGEMA_signal_2322), .Z1_t (new_AGEMA_signal_2323), .Z1_f (new_AGEMA_signal_2324) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_U13 ( .A0_t (SubCellInst_SboxInst_7_n8), .A0_f (new_AGEMA_signal_1391), .A1_t (new_AGEMA_signal_1392), .A1_f (new_AGEMA_signal_1393), .B0_t (SubCellInst_SboxInst_7_n7), .B0_f (new_AGEMA_signal_2736), .B1_t (new_AGEMA_signal_2737), .B1_f (new_AGEMA_signal_2738), .Z0_t (Feedback[28]), .Z0_f (new_AGEMA_signal_3265), .Z1_t (new_AGEMA_signal_3266), .Z1_f (new_AGEMA_signal_3267) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_U12 ( .A0_t (Output_s0_t[37]), .A0_f (Output_s0_f[37]), .A1_t (Output_s1_t[37]), .A1_f (Output_s1_f[37]), .B0_t (SubCellInst_SboxInst_7_n6), .B0_f (new_AGEMA_signal_2325), .B1_t (new_AGEMA_signal_2326), .B1_f (new_AGEMA_signal_2327), .Z0_t (SubCellInst_SboxInst_7_n7), .Z0_f (new_AGEMA_signal_2736), .Z1_t (new_AGEMA_signal_2737), .Z1_f (new_AGEMA_signal_2738) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_U11 ( .A0_t (Output_s0_t[36]), .A0_f (Output_s0_f[36]), .A1_t (Output_s1_t[36]), .A1_f (Output_s1_f[36]), .B0_t (SubCellInst_SboxInst_7_n5), .B0_f (new_AGEMA_signal_1388), .B1_t (new_AGEMA_signal_1389), .B1_f (new_AGEMA_signal_1390), .Z0_t (SubCellInst_SboxInst_7_n6), .Z0_f (new_AGEMA_signal_2325), .Z1_t (new_AGEMA_signal_2326), .Z1_f (new_AGEMA_signal_2327) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_U10 ( .A0_t (Output_s0_t[39]), .A0_f (Output_s0_f[39]), .A1_t (Output_s1_t[39]), .A1_f (Output_s1_f[39]), .B0_t (Output_s0_t[38]), .B0_f (Output_s0_f[38]), .B1_t (Output_s1_t[38]), .B1_f (Output_s1_f[38]), .Z0_t (SubCellInst_SboxInst_7_n5), .Z0_f (new_AGEMA_signal_1388), .Z1_t (new_AGEMA_signal_1389), .Z1_f (new_AGEMA_signal_1390) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_U9 ( .A0_t (Output_s0_t[39]), .A0_f (Output_s0_f[39]), .A1_t (Output_s1_t[39]), .A1_f (Output_s1_f[39]), .B0_t (Output_s0_t[38]), .B0_f (Output_s0_f[38]), .B1_t (Output_s1_t[38]), .B1_f (Output_s1_f[38]), .Z0_t (SubCellInst_SboxInst_7_n8), .Z0_f (new_AGEMA_signal_1391), .Z1_t (new_AGEMA_signal_1392), .Z1_f (new_AGEMA_signal_1393) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U8 ( .A0_t (SubCellInst_SboxInst_7_n10), .A0_f (new_AGEMA_signal_1397), .A1_t (new_AGEMA_signal_1398), .A1_f (new_AGEMA_signal_1399), .B0_t (SubCellInst_SboxInst_7_n3), .B0_f (new_AGEMA_signal_2739), .B1_t (new_AGEMA_signal_2740), .B1_f (new_AGEMA_signal_2741), .Z0_t (Feedback[30]), .Z0_f (new_AGEMA_signal_3268), .Z1_t (new_AGEMA_signal_3269), .Z1_f (new_AGEMA_signal_3270) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U7 ( .A0_t (SubCellInst_SboxInst_7_n2), .A0_f (new_AGEMA_signal_2328), .A1_t (new_AGEMA_signal_2329), .A1_f (new_AGEMA_signal_2330), .B0_t (Output_s0_t[37]), .B0_f (Output_s0_f[37]), .B1_t (Output_s1_t[37]), .B1_f (Output_s1_f[37]), .Z0_t (SubCellInst_SboxInst_7_n3), .Z0_f (new_AGEMA_signal_2739), .Z1_t (new_AGEMA_signal_2740), .Z1_f (new_AGEMA_signal_2741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U6 ( .A0_t (SubCellInst_SboxInst_7_n1), .A0_f (new_AGEMA_signal_1394), .A1_t (new_AGEMA_signal_1395), .A1_f (new_AGEMA_signal_1396), .B0_t (Output_s0_t[38]), .B0_f (Output_s0_f[38]), .B1_t (Output_s1_t[38]), .B1_f (Output_s1_f[38]), .Z0_t (SubCellInst_SboxInst_7_n2), .Z0_f (new_AGEMA_signal_2328), .Z1_t (new_AGEMA_signal_2329), .Z1_f (new_AGEMA_signal_2330) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U4 ( .A0_t (Output_s0_t[39]), .A0_f (Output_s0_f[39]), .A1_t (Output_s1_t[39]), .A1_f (Output_s1_f[39]), .B0_t (Output_s0_t[36]), .B0_f (Output_s0_f[36]), .B1_t (Output_s1_t[36]), .B1_f (Output_s1_f[36]), .Z0_t (SubCellInst_SboxInst_7_n1), .Z0_f (new_AGEMA_signal_1394), .Z1_t (new_AGEMA_signal_1395), .Z1_f (new_AGEMA_signal_1396) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_U3 ( .A0_t (Output_s0_t[36]), .A0_f (Output_s0_f[36]), .A1_t (Output_s1_t[36]), .A1_f (Output_s1_f[36]), .B0_t (Output_s0_t[39]), .B0_f (Output_s0_f[39]), .B1_t (Output_s1_t[39]), .B1_f (Output_s1_f[39]), .Z0_t (SubCellInst_SboxInst_7_n10), .Z0_f (new_AGEMA_signal_1397), .Z1_t (new_AGEMA_signal_1398), .Z1_f (new_AGEMA_signal_1399) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U19 ( .A0_t (SubCellInst_SboxInst_8_n15), .A0_f (new_AGEMA_signal_1409), .A1_t (new_AGEMA_signal_1410), .A1_f (new_AGEMA_signal_1411), .B0_t (SubCellInst_SboxInst_8_n14), .B0_f (new_AGEMA_signal_2331), .B1_t (new_AGEMA_signal_2332), .B1_f (new_AGEMA_signal_2333), .Z0_t (Feedback[33]), .Z0_f (new_AGEMA_signal_2742), .Z1_t (new_AGEMA_signal_2743), .Z1_f (new_AGEMA_signal_2744) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U18 ( .A0_t (Output_s0_t[16]), .A0_f (Output_s0_f[16]), .A1_t (Output_s1_t[16]), .A1_f (Output_s1_f[16]), .B0_t (SubCellInst_SboxInst_8_n13), .B0_f (new_AGEMA_signal_1406), .B1_t (new_AGEMA_signal_1407), .B1_f (new_AGEMA_signal_1408), .Z0_t (SubCellInst_SboxInst_8_n14), .Z0_f (new_AGEMA_signal_2331), .Z1_t (new_AGEMA_signal_2332), .Z1_f (new_AGEMA_signal_2333) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U17 ( .A0_t (Output_s0_t[19]), .A0_f (Output_s0_f[19]), .A1_t (Output_s1_t[19]), .A1_f (Output_s1_f[19]), .B0_t (Output_s0_t[18]), .B0_f (Output_s0_f[18]), .B1_t (Output_s1_t[18]), .B1_f (Output_s1_f[18]), .Z0_t (SubCellInst_SboxInst_8_n13), .Z0_f (new_AGEMA_signal_1406), .Z1_t (new_AGEMA_signal_1407), .Z1_f (new_AGEMA_signal_1408) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U16 ( .A0_t (Output_s0_t[18]), .A0_f (Output_s0_f[18]), .A1_t (Output_s1_t[18]), .A1_f (Output_s1_f[18]), .B0_t (Output_s0_t[19]), .B0_f (Output_s0_f[19]), .B1_t (Output_s1_t[19]), .B1_f (Output_s1_f[19]), .Z0_t (SubCellInst_SboxInst_8_n15), .Z0_f (new_AGEMA_signal_1409), .Z1_t (new_AGEMA_signal_1410), .Z1_f (new_AGEMA_signal_1411) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U15 ( .A0_t (SubCellInst_SboxInst_8_n10), .A0_f (new_AGEMA_signal_1418), .A1_t (new_AGEMA_signal_1419), .A1_f (new_AGEMA_signal_1420), .B0_t (SubCellInst_SboxInst_8_n9), .B0_f (new_AGEMA_signal_2337), .B1_t (new_AGEMA_signal_2338), .B1_f (new_AGEMA_signal_2339), .Z0_t (Feedback[35]), .Z0_f (new_AGEMA_signal_2745), .Z1_t (new_AGEMA_signal_2746), .Z1_f (new_AGEMA_signal_2747) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U14 ( .A0_t (SubCellInst_SboxInst_8_n8), .A0_f (new_AGEMA_signal_1424), .A1_t (new_AGEMA_signal_1425), .A1_f (new_AGEMA_signal_1426), .B0_t (Output_s0_t[17]), .B0_f (Output_s0_f[17]), .B1_t (Output_s1_t[17]), .B1_f (Output_s1_f[17]), .Z0_t (SubCellInst_SboxInst_8_n9), .Z0_f (new_AGEMA_signal_2337), .Z1_t (new_AGEMA_signal_2338), .Z1_f (new_AGEMA_signal_2339) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U13 ( .A0_t (SubCellInst_SboxInst_8_n10), .A0_f (new_AGEMA_signal_1418), .A1_t (new_AGEMA_signal_1419), .A1_f (new_AGEMA_signal_1420), .B0_t (SubCellInst_SboxInst_8_n7), .B0_f (new_AGEMA_signal_2748), .B1_t (new_AGEMA_signal_2749), .B1_f (new_AGEMA_signal_2750), .Z0_t (Feedback[34]), .Z0_f (new_AGEMA_signal_3271), .Z1_t (new_AGEMA_signal_3272), .Z1_f (new_AGEMA_signal_3273) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U12 ( .A0_t (SubCellInst_SboxInst_8_n6), .A0_f (new_AGEMA_signal_2340), .A1_t (new_AGEMA_signal_2341), .A1_f (new_AGEMA_signal_2342), .B0_t (Output_s0_t[17]), .B0_f (Output_s0_f[17]), .B1_t (Output_s1_t[17]), .B1_f (Output_s1_f[17]), .Z0_t (SubCellInst_SboxInst_8_n7), .Z0_f (new_AGEMA_signal_2748), .Z1_t (new_AGEMA_signal_2749), .Z1_f (new_AGEMA_signal_2750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U11 ( .A0_t (SubCellInst_SboxInst_8_n5), .A0_f (new_AGEMA_signal_1415), .A1_t (new_AGEMA_signal_1416), .A1_f (new_AGEMA_signal_1417), .B0_t (Output_s0_t[18]), .B0_f (Output_s0_f[18]), .B1_t (Output_s1_t[18]), .B1_f (Output_s1_f[18]), .Z0_t (SubCellInst_SboxInst_8_n6), .Z0_f (new_AGEMA_signal_2340), .Z1_t (new_AGEMA_signal_2341), .Z1_f (new_AGEMA_signal_2342) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U10 ( .A0_t (Output_s0_t[16]), .A0_f (Output_s0_f[16]), .A1_t (Output_s1_t[16]), .A1_f (Output_s1_f[16]), .B0_t (Output_s0_t[19]), .B0_f (Output_s0_f[19]), .B1_t (Output_s1_t[19]), .B1_f (Output_s1_f[19]), .Z0_t (SubCellInst_SboxInst_8_n5), .Z0_f (new_AGEMA_signal_1415), .Z1_t (new_AGEMA_signal_1416), .Z1_f (new_AGEMA_signal_1417) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_U9 ( .A0_t (Output_s0_t[19]), .A0_f (Output_s0_f[19]), .A1_t (Output_s1_t[19]), .A1_f (Output_s1_f[19]), .B0_t (Output_s0_t[16]), .B0_f (Output_s0_f[16]), .B1_t (Output_s1_t[16]), .B1_f (Output_s1_f[16]), .Z0_t (SubCellInst_SboxInst_8_n10), .Z0_f (new_AGEMA_signal_1418), .Z1_t (new_AGEMA_signal_1419), .Z1_f (new_AGEMA_signal_1420) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_U8 ( .A0_t (SubCellInst_SboxInst_8_n8), .A0_f (new_AGEMA_signal_1424), .A1_t (new_AGEMA_signal_1425), .A1_f (new_AGEMA_signal_1426), .B0_t (SubCellInst_SboxInst_8_n3), .B0_f (new_AGEMA_signal_2751), .B1_t (new_AGEMA_signal_2752), .B1_f (new_AGEMA_signal_2753), .Z0_t (Feedback[32]), .Z0_f (new_AGEMA_signal_3274), .Z1_t (new_AGEMA_signal_3275), .Z1_f (new_AGEMA_signal_3276) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_U7 ( .A0_t (Output_s0_t[17]), .A0_f (Output_s0_f[17]), .A1_t (Output_s1_t[17]), .A1_f (Output_s1_f[17]), .B0_t (SubCellInst_SboxInst_8_n2), .B0_f (new_AGEMA_signal_2343), .B1_t (new_AGEMA_signal_2344), .B1_f (new_AGEMA_signal_2345), .Z0_t (SubCellInst_SboxInst_8_n3), .Z0_f (new_AGEMA_signal_2751), .Z1_t (new_AGEMA_signal_2752), .Z1_f (new_AGEMA_signal_2753) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_U6 ( .A0_t (Output_s0_t[16]), .A0_f (Output_s0_f[16]), .A1_t (Output_s1_t[16]), .A1_f (Output_s1_f[16]), .B0_t (SubCellInst_SboxInst_8_n1), .B0_f (new_AGEMA_signal_1421), .B1_t (new_AGEMA_signal_1422), .B1_f (new_AGEMA_signal_1423), .Z0_t (SubCellInst_SboxInst_8_n2), .Z0_f (new_AGEMA_signal_2343), .Z1_t (new_AGEMA_signal_2344), .Z1_f (new_AGEMA_signal_2345) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_U5 ( .A0_t (Output_s0_t[18]), .A0_f (Output_s0_f[18]), .A1_t (Output_s1_t[18]), .A1_f (Output_s1_f[18]), .B0_t (Output_s0_t[19]), .B0_f (Output_s0_f[19]), .B1_t (Output_s1_t[19]), .B1_f (Output_s1_f[19]), .Z0_t (SubCellInst_SboxInst_8_n1), .Z0_f (new_AGEMA_signal_1421), .Z1_t (new_AGEMA_signal_1422), .Z1_f (new_AGEMA_signal_1423) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_U3 ( .A0_t (Output_s0_t[18]), .A0_f (Output_s0_f[18]), .A1_t (Output_s1_t[18]), .A1_f (Output_s1_f[18]), .B0_t (Output_s0_t[19]), .B0_f (Output_s0_f[19]), .B1_t (Output_s1_t[19]), .B1_f (Output_s1_f[19]), .Z0_t (SubCellInst_SboxInst_8_n8), .Z0_f (new_AGEMA_signal_1424), .Z1_t (new_AGEMA_signal_1425), .Z1_f (new_AGEMA_signal_1426) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U19 ( .A0_t (SubCellInst_SboxInst_9_n15), .A0_f (new_AGEMA_signal_1436), .A1_t (new_AGEMA_signal_1437), .A1_f (new_AGEMA_signal_1438), .B0_t (SubCellInst_SboxInst_9_n14), .B0_f (new_AGEMA_signal_2346), .B1_t (new_AGEMA_signal_2347), .B1_f (new_AGEMA_signal_2348), .Z0_t (Feedback[37]), .Z0_f (new_AGEMA_signal_2754), .Z1_t (new_AGEMA_signal_2755), .Z1_f (new_AGEMA_signal_2756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U18 ( .A0_t (Output_s0_t[28]), .A0_f (Output_s0_f[28]), .A1_t (Output_s1_t[28]), .A1_f (Output_s1_f[28]), .B0_t (SubCellInst_SboxInst_9_n13), .B0_f (new_AGEMA_signal_1433), .B1_t (new_AGEMA_signal_1434), .B1_f (new_AGEMA_signal_1435), .Z0_t (SubCellInst_SboxInst_9_n14), .Z0_f (new_AGEMA_signal_2346), .Z1_t (new_AGEMA_signal_2347), .Z1_f (new_AGEMA_signal_2348) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U17 ( .A0_t (Output_s0_t[31]), .A0_f (Output_s0_f[31]), .A1_t (Output_s1_t[31]), .A1_f (Output_s1_f[31]), .B0_t (Output_s0_t[30]), .B0_f (Output_s0_f[30]), .B1_t (Output_s1_t[30]), .B1_f (Output_s1_f[30]), .Z0_t (SubCellInst_SboxInst_9_n13), .Z0_f (new_AGEMA_signal_1433), .Z1_t (new_AGEMA_signal_1434), .Z1_f (new_AGEMA_signal_1435) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U16 ( .A0_t (Output_s0_t[30]), .A0_f (Output_s0_f[30]), .A1_t (Output_s1_t[30]), .A1_f (Output_s1_f[30]), .B0_t (Output_s0_t[31]), .B0_f (Output_s0_f[31]), .B1_t (Output_s1_t[31]), .B1_f (Output_s1_f[31]), .Z0_t (SubCellInst_SboxInst_9_n15), .Z0_f (new_AGEMA_signal_1436), .Z1_t (new_AGEMA_signal_1437), .Z1_f (new_AGEMA_signal_1438) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U15 ( .A0_t (SubCellInst_SboxInst_9_n10), .A0_f (new_AGEMA_signal_1445), .A1_t (new_AGEMA_signal_1446), .A1_f (new_AGEMA_signal_1447), .B0_t (SubCellInst_SboxInst_9_n9), .B0_f (new_AGEMA_signal_2352), .B1_t (new_AGEMA_signal_2353), .B1_f (new_AGEMA_signal_2354), .Z0_t (Feedback[39]), .Z0_f (new_AGEMA_signal_2757), .Z1_t (new_AGEMA_signal_2758), .Z1_f (new_AGEMA_signal_2759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U14 ( .A0_t (SubCellInst_SboxInst_9_n8), .A0_f (new_AGEMA_signal_1451), .A1_t (new_AGEMA_signal_1452), .A1_f (new_AGEMA_signal_1453), .B0_t (Output_s0_t[29]), .B0_f (Output_s0_f[29]), .B1_t (Output_s1_t[29]), .B1_f (Output_s1_f[29]), .Z0_t (SubCellInst_SboxInst_9_n9), .Z0_f (new_AGEMA_signal_2352), .Z1_t (new_AGEMA_signal_2353), .Z1_f (new_AGEMA_signal_2354) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U13 ( .A0_t (SubCellInst_SboxInst_9_n10), .A0_f (new_AGEMA_signal_1445), .A1_t (new_AGEMA_signal_1446), .A1_f (new_AGEMA_signal_1447), .B0_t (SubCellInst_SboxInst_9_n7), .B0_f (new_AGEMA_signal_2760), .B1_t (new_AGEMA_signal_2761), .B1_f (new_AGEMA_signal_2762), .Z0_t (Feedback[38]), .Z0_f (new_AGEMA_signal_3277), .Z1_t (new_AGEMA_signal_3278), .Z1_f (new_AGEMA_signal_3279) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U12 ( .A0_t (SubCellInst_SboxInst_9_n6), .A0_f (new_AGEMA_signal_2355), .A1_t (new_AGEMA_signal_2356), .A1_f (new_AGEMA_signal_2357), .B0_t (Output_s0_t[29]), .B0_f (Output_s0_f[29]), .B1_t (Output_s1_t[29]), .B1_f (Output_s1_f[29]), .Z0_t (SubCellInst_SboxInst_9_n7), .Z0_f (new_AGEMA_signal_2760), .Z1_t (new_AGEMA_signal_2761), .Z1_f (new_AGEMA_signal_2762) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U11 ( .A0_t (SubCellInst_SboxInst_9_n5), .A0_f (new_AGEMA_signal_1442), .A1_t (new_AGEMA_signal_1443), .A1_f (new_AGEMA_signal_1444), .B0_t (Output_s0_t[30]), .B0_f (Output_s0_f[30]), .B1_t (Output_s1_t[30]), .B1_f (Output_s1_f[30]), .Z0_t (SubCellInst_SboxInst_9_n6), .Z0_f (new_AGEMA_signal_2355), .Z1_t (new_AGEMA_signal_2356), .Z1_f (new_AGEMA_signal_2357) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U10 ( .A0_t (Output_s0_t[28]), .A0_f (Output_s0_f[28]), .A1_t (Output_s1_t[28]), .A1_f (Output_s1_f[28]), .B0_t (Output_s0_t[31]), .B0_f (Output_s0_f[31]), .B1_t (Output_s1_t[31]), .B1_f (Output_s1_f[31]), .Z0_t (SubCellInst_SboxInst_9_n5), .Z0_f (new_AGEMA_signal_1442), .Z1_t (new_AGEMA_signal_1443), .Z1_f (new_AGEMA_signal_1444) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_U9 ( .A0_t (Output_s0_t[31]), .A0_f (Output_s0_f[31]), .A1_t (Output_s1_t[31]), .A1_f (Output_s1_f[31]), .B0_t (Output_s0_t[28]), .B0_f (Output_s0_f[28]), .B1_t (Output_s1_t[28]), .B1_f (Output_s1_f[28]), .Z0_t (SubCellInst_SboxInst_9_n10), .Z0_f (new_AGEMA_signal_1445), .Z1_t (new_AGEMA_signal_1446), .Z1_f (new_AGEMA_signal_1447) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_U8 ( .A0_t (SubCellInst_SboxInst_9_n8), .A0_f (new_AGEMA_signal_1451), .A1_t (new_AGEMA_signal_1452), .A1_f (new_AGEMA_signal_1453), .B0_t (SubCellInst_SboxInst_9_n3), .B0_f (new_AGEMA_signal_2763), .B1_t (new_AGEMA_signal_2764), .B1_f (new_AGEMA_signal_2765), .Z0_t (Feedback[36]), .Z0_f (new_AGEMA_signal_3280), .Z1_t (new_AGEMA_signal_3281), .Z1_f (new_AGEMA_signal_3282) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_U7 ( .A0_t (Output_s0_t[29]), .A0_f (Output_s0_f[29]), .A1_t (Output_s1_t[29]), .A1_f (Output_s1_f[29]), .B0_t (SubCellInst_SboxInst_9_n2), .B0_f (new_AGEMA_signal_2358), .B1_t (new_AGEMA_signal_2359), .B1_f (new_AGEMA_signal_2360), .Z0_t (SubCellInst_SboxInst_9_n3), .Z0_f (new_AGEMA_signal_2763), .Z1_t (new_AGEMA_signal_2764), .Z1_f (new_AGEMA_signal_2765) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_U6 ( .A0_t (Output_s0_t[28]), .A0_f (Output_s0_f[28]), .A1_t (Output_s1_t[28]), .A1_f (Output_s1_f[28]), .B0_t (SubCellInst_SboxInst_9_n1), .B0_f (new_AGEMA_signal_1448), .B1_t (new_AGEMA_signal_1449), .B1_f (new_AGEMA_signal_1450), .Z0_t (SubCellInst_SboxInst_9_n2), .Z0_f (new_AGEMA_signal_2358), .Z1_t (new_AGEMA_signal_2359), .Z1_f (new_AGEMA_signal_2360) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_U5 ( .A0_t (Output_s0_t[30]), .A0_f (Output_s0_f[30]), .A1_t (Output_s1_t[30]), .A1_f (Output_s1_f[30]), .B0_t (Output_s0_t[31]), .B0_f (Output_s0_f[31]), .B1_t (Output_s1_t[31]), .B1_f (Output_s1_f[31]), .Z0_t (SubCellInst_SboxInst_9_n1), .Z0_f (new_AGEMA_signal_1448), .Z1_t (new_AGEMA_signal_1449), .Z1_f (new_AGEMA_signal_1450) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_U3 ( .A0_t (Output_s0_t[30]), .A0_f (Output_s0_f[30]), .A1_t (Output_s1_t[30]), .A1_f (Output_s1_f[30]), .B0_t (Output_s0_t[31]), .B0_f (Output_s0_f[31]), .B1_t (Output_s1_t[31]), .B1_f (Output_s1_f[31]), .Z0_t (SubCellInst_SboxInst_9_n8), .Z0_f (new_AGEMA_signal_1451), .Z1_t (new_AGEMA_signal_1452), .Z1_f (new_AGEMA_signal_1453) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U19 ( .A0_t (SubCellInst_SboxInst_10_n15), .A0_f (new_AGEMA_signal_1463), .A1_t (new_AGEMA_signal_1464), .A1_f (new_AGEMA_signal_1465), .B0_t (SubCellInst_SboxInst_10_n14), .B0_f (new_AGEMA_signal_2361), .B1_t (new_AGEMA_signal_2362), .B1_f (new_AGEMA_signal_2363), .Z0_t (Feedback[41]), .Z0_f (new_AGEMA_signal_2766), .Z1_t (new_AGEMA_signal_2767), .Z1_f (new_AGEMA_signal_2768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U18 ( .A0_t (Output_s0_t[24]), .A0_f (Output_s0_f[24]), .A1_t (Output_s1_t[24]), .A1_f (Output_s1_f[24]), .B0_t (SubCellInst_SboxInst_10_n13), .B0_f (new_AGEMA_signal_1460), .B1_t (new_AGEMA_signal_1461), .B1_f (new_AGEMA_signal_1462), .Z0_t (SubCellInst_SboxInst_10_n14), .Z0_f (new_AGEMA_signal_2361), .Z1_t (new_AGEMA_signal_2362), .Z1_f (new_AGEMA_signal_2363) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U17 ( .A0_t (Output_s0_t[27]), .A0_f (Output_s0_f[27]), .A1_t (Output_s1_t[27]), .A1_f (Output_s1_f[27]), .B0_t (Output_s0_t[26]), .B0_f (Output_s0_f[26]), .B1_t (Output_s1_t[26]), .B1_f (Output_s1_f[26]), .Z0_t (SubCellInst_SboxInst_10_n13), .Z0_f (new_AGEMA_signal_1460), .Z1_t (new_AGEMA_signal_1461), .Z1_f (new_AGEMA_signal_1462) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U16 ( .A0_t (Output_s0_t[26]), .A0_f (Output_s0_f[26]), .A1_t (Output_s1_t[26]), .A1_f (Output_s1_f[26]), .B0_t (Output_s0_t[27]), .B0_f (Output_s0_f[27]), .B1_t (Output_s1_t[27]), .B1_f (Output_s1_f[27]), .Z0_t (SubCellInst_SboxInst_10_n15), .Z0_f (new_AGEMA_signal_1463), .Z1_t (new_AGEMA_signal_1464), .Z1_f (new_AGEMA_signal_1465) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U15 ( .A0_t (SubCellInst_SboxInst_10_n10), .A0_f (new_AGEMA_signal_1472), .A1_t (new_AGEMA_signal_1473), .A1_f (new_AGEMA_signal_1474), .B0_t (SubCellInst_SboxInst_10_n9), .B0_f (new_AGEMA_signal_2367), .B1_t (new_AGEMA_signal_2368), .B1_f (new_AGEMA_signal_2369), .Z0_t (Feedback[43]), .Z0_f (new_AGEMA_signal_2769), .Z1_t (new_AGEMA_signal_2770), .Z1_f (new_AGEMA_signal_2771) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U14 ( .A0_t (SubCellInst_SboxInst_10_n8), .A0_f (new_AGEMA_signal_1478), .A1_t (new_AGEMA_signal_1479), .A1_f (new_AGEMA_signal_1480), .B0_t (Output_s0_t[25]), .B0_f (Output_s0_f[25]), .B1_t (Output_s1_t[25]), .B1_f (Output_s1_f[25]), .Z0_t (SubCellInst_SboxInst_10_n9), .Z0_f (new_AGEMA_signal_2367), .Z1_t (new_AGEMA_signal_2368), .Z1_f (new_AGEMA_signal_2369) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U13 ( .A0_t (SubCellInst_SboxInst_10_n10), .A0_f (new_AGEMA_signal_1472), .A1_t (new_AGEMA_signal_1473), .A1_f (new_AGEMA_signal_1474), .B0_t (SubCellInst_SboxInst_10_n7), .B0_f (new_AGEMA_signal_2772), .B1_t (new_AGEMA_signal_2773), .B1_f (new_AGEMA_signal_2774), .Z0_t (Feedback[42]), .Z0_f (new_AGEMA_signal_3283), .Z1_t (new_AGEMA_signal_3284), .Z1_f (new_AGEMA_signal_3285) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U12 ( .A0_t (SubCellInst_SboxInst_10_n6), .A0_f (new_AGEMA_signal_2370), .A1_t (new_AGEMA_signal_2371), .A1_f (new_AGEMA_signal_2372), .B0_t (Output_s0_t[25]), .B0_f (Output_s0_f[25]), .B1_t (Output_s1_t[25]), .B1_f (Output_s1_f[25]), .Z0_t (SubCellInst_SboxInst_10_n7), .Z0_f (new_AGEMA_signal_2772), .Z1_t (new_AGEMA_signal_2773), .Z1_f (new_AGEMA_signal_2774) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U11 ( .A0_t (SubCellInst_SboxInst_10_n5), .A0_f (new_AGEMA_signal_1469), .A1_t (new_AGEMA_signal_1470), .A1_f (new_AGEMA_signal_1471), .B0_t (Output_s0_t[26]), .B0_f (Output_s0_f[26]), .B1_t (Output_s1_t[26]), .B1_f (Output_s1_f[26]), .Z0_t (SubCellInst_SboxInst_10_n6), .Z0_f (new_AGEMA_signal_2370), .Z1_t (new_AGEMA_signal_2371), .Z1_f (new_AGEMA_signal_2372) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U10 ( .A0_t (Output_s0_t[24]), .A0_f (Output_s0_f[24]), .A1_t (Output_s1_t[24]), .A1_f (Output_s1_f[24]), .B0_t (Output_s0_t[27]), .B0_f (Output_s0_f[27]), .B1_t (Output_s1_t[27]), .B1_f (Output_s1_f[27]), .Z0_t (SubCellInst_SboxInst_10_n5), .Z0_f (new_AGEMA_signal_1469), .Z1_t (new_AGEMA_signal_1470), .Z1_f (new_AGEMA_signal_1471) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_U9 ( .A0_t (Output_s0_t[27]), .A0_f (Output_s0_f[27]), .A1_t (Output_s1_t[27]), .A1_f (Output_s1_f[27]), .B0_t (Output_s0_t[24]), .B0_f (Output_s0_f[24]), .B1_t (Output_s1_t[24]), .B1_f (Output_s1_f[24]), .Z0_t (SubCellInst_SboxInst_10_n10), .Z0_f (new_AGEMA_signal_1472), .Z1_t (new_AGEMA_signal_1473), .Z1_f (new_AGEMA_signal_1474) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_U8 ( .A0_t (SubCellInst_SboxInst_10_n8), .A0_f (new_AGEMA_signal_1478), .A1_t (new_AGEMA_signal_1479), .A1_f (new_AGEMA_signal_1480), .B0_t (SubCellInst_SboxInst_10_n3), .B0_f (new_AGEMA_signal_2775), .B1_t (new_AGEMA_signal_2776), .B1_f (new_AGEMA_signal_2777), .Z0_t (Feedback[40]), .Z0_f (new_AGEMA_signal_3286), .Z1_t (new_AGEMA_signal_3287), .Z1_f (new_AGEMA_signal_3288) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_U7 ( .A0_t (Output_s0_t[25]), .A0_f (Output_s0_f[25]), .A1_t (Output_s1_t[25]), .A1_f (Output_s1_f[25]), .B0_t (SubCellInst_SboxInst_10_n2), .B0_f (new_AGEMA_signal_2373), .B1_t (new_AGEMA_signal_2374), .B1_f (new_AGEMA_signal_2375), .Z0_t (SubCellInst_SboxInst_10_n3), .Z0_f (new_AGEMA_signal_2775), .Z1_t (new_AGEMA_signal_2776), .Z1_f (new_AGEMA_signal_2777) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_U6 ( .A0_t (Output_s0_t[24]), .A0_f (Output_s0_f[24]), .A1_t (Output_s1_t[24]), .A1_f (Output_s1_f[24]), .B0_t (SubCellInst_SboxInst_10_n1), .B0_f (new_AGEMA_signal_1475), .B1_t (new_AGEMA_signal_1476), .B1_f (new_AGEMA_signal_1477), .Z0_t (SubCellInst_SboxInst_10_n2), .Z0_f (new_AGEMA_signal_2373), .Z1_t (new_AGEMA_signal_2374), .Z1_f (new_AGEMA_signal_2375) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_U5 ( .A0_t (Output_s0_t[26]), .A0_f (Output_s0_f[26]), .A1_t (Output_s1_t[26]), .A1_f (Output_s1_f[26]), .B0_t (Output_s0_t[27]), .B0_f (Output_s0_f[27]), .B1_t (Output_s1_t[27]), .B1_f (Output_s1_f[27]), .Z0_t (SubCellInst_SboxInst_10_n1), .Z0_f (new_AGEMA_signal_1475), .Z1_t (new_AGEMA_signal_1476), .Z1_f (new_AGEMA_signal_1477) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_U3 ( .A0_t (Output_s0_t[26]), .A0_f (Output_s0_f[26]), .A1_t (Output_s1_t[26]), .A1_f (Output_s1_f[26]), .B0_t (Output_s0_t[27]), .B0_f (Output_s0_f[27]), .B1_t (Output_s1_t[27]), .B1_f (Output_s1_f[27]), .Z0_t (SubCellInst_SboxInst_10_n8), .Z0_f (new_AGEMA_signal_1478), .Z1_t (new_AGEMA_signal_1479), .Z1_f (new_AGEMA_signal_1480) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U19 ( .A0_t (SubCellInst_SboxInst_11_n15), .A0_f (new_AGEMA_signal_1490), .A1_t (new_AGEMA_signal_1491), .A1_f (new_AGEMA_signal_1492), .B0_t (SubCellInst_SboxInst_11_n14), .B0_f (new_AGEMA_signal_2376), .B1_t (new_AGEMA_signal_2377), .B1_f (new_AGEMA_signal_2378), .Z0_t (Feedback[45]), .Z0_f (new_AGEMA_signal_2778), .Z1_t (new_AGEMA_signal_2779), .Z1_f (new_AGEMA_signal_2780) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U18 ( .A0_t (Output_s0_t[20]), .A0_f (Output_s0_f[20]), .A1_t (Output_s1_t[20]), .A1_f (Output_s1_f[20]), .B0_t (SubCellInst_SboxInst_11_n13), .B0_f (new_AGEMA_signal_1487), .B1_t (new_AGEMA_signal_1488), .B1_f (new_AGEMA_signal_1489), .Z0_t (SubCellInst_SboxInst_11_n14), .Z0_f (new_AGEMA_signal_2376), .Z1_t (new_AGEMA_signal_2377), .Z1_f (new_AGEMA_signal_2378) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U17 ( .A0_t (Output_s0_t[23]), .A0_f (Output_s0_f[23]), .A1_t (Output_s1_t[23]), .A1_f (Output_s1_f[23]), .B0_t (Output_s0_t[22]), .B0_f (Output_s0_f[22]), .B1_t (Output_s1_t[22]), .B1_f (Output_s1_f[22]), .Z0_t (SubCellInst_SboxInst_11_n13), .Z0_f (new_AGEMA_signal_1487), .Z1_t (new_AGEMA_signal_1488), .Z1_f (new_AGEMA_signal_1489) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U16 ( .A0_t (Output_s0_t[22]), .A0_f (Output_s0_f[22]), .A1_t (Output_s1_t[22]), .A1_f (Output_s1_f[22]), .B0_t (Output_s0_t[23]), .B0_f (Output_s0_f[23]), .B1_t (Output_s1_t[23]), .B1_f (Output_s1_f[23]), .Z0_t (SubCellInst_SboxInst_11_n15), .Z0_f (new_AGEMA_signal_1490), .Z1_t (new_AGEMA_signal_1491), .Z1_f (new_AGEMA_signal_1492) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U15 ( .A0_t (SubCellInst_SboxInst_11_n10), .A0_f (new_AGEMA_signal_1499), .A1_t (new_AGEMA_signal_1500), .A1_f (new_AGEMA_signal_1501), .B0_t (SubCellInst_SboxInst_11_n9), .B0_f (new_AGEMA_signal_2382), .B1_t (new_AGEMA_signal_2383), .B1_f (new_AGEMA_signal_2384), .Z0_t (Feedback[47]), .Z0_f (new_AGEMA_signal_2781), .Z1_t (new_AGEMA_signal_2782), .Z1_f (new_AGEMA_signal_2783) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U14 ( .A0_t (SubCellInst_SboxInst_11_n8), .A0_f (new_AGEMA_signal_1505), .A1_t (new_AGEMA_signal_1506), .A1_f (new_AGEMA_signal_1507), .B0_t (Output_s0_t[21]), .B0_f (Output_s0_f[21]), .B1_t (Output_s1_t[21]), .B1_f (Output_s1_f[21]), .Z0_t (SubCellInst_SboxInst_11_n9), .Z0_f (new_AGEMA_signal_2382), .Z1_t (new_AGEMA_signal_2383), .Z1_f (new_AGEMA_signal_2384) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U13 ( .A0_t (SubCellInst_SboxInst_11_n10), .A0_f (new_AGEMA_signal_1499), .A1_t (new_AGEMA_signal_1500), .A1_f (new_AGEMA_signal_1501), .B0_t (SubCellInst_SboxInst_11_n7), .B0_f (new_AGEMA_signal_2784), .B1_t (new_AGEMA_signal_2785), .B1_f (new_AGEMA_signal_2786), .Z0_t (Feedback[46]), .Z0_f (new_AGEMA_signal_3289), .Z1_t (new_AGEMA_signal_3290), .Z1_f (new_AGEMA_signal_3291) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U12 ( .A0_t (SubCellInst_SboxInst_11_n6), .A0_f (new_AGEMA_signal_2385), .A1_t (new_AGEMA_signal_2386), .A1_f (new_AGEMA_signal_2387), .B0_t (Output_s0_t[21]), .B0_f (Output_s0_f[21]), .B1_t (Output_s1_t[21]), .B1_f (Output_s1_f[21]), .Z0_t (SubCellInst_SboxInst_11_n7), .Z0_f (new_AGEMA_signal_2784), .Z1_t (new_AGEMA_signal_2785), .Z1_f (new_AGEMA_signal_2786) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U11 ( .A0_t (SubCellInst_SboxInst_11_n5), .A0_f (new_AGEMA_signal_1496), .A1_t (new_AGEMA_signal_1497), .A1_f (new_AGEMA_signal_1498), .B0_t (Output_s0_t[22]), .B0_f (Output_s0_f[22]), .B1_t (Output_s1_t[22]), .B1_f (Output_s1_f[22]), .Z0_t (SubCellInst_SboxInst_11_n6), .Z0_f (new_AGEMA_signal_2385), .Z1_t (new_AGEMA_signal_2386), .Z1_f (new_AGEMA_signal_2387) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U10 ( .A0_t (Output_s0_t[20]), .A0_f (Output_s0_f[20]), .A1_t (Output_s1_t[20]), .A1_f (Output_s1_f[20]), .B0_t (Output_s0_t[23]), .B0_f (Output_s0_f[23]), .B1_t (Output_s1_t[23]), .B1_f (Output_s1_f[23]), .Z0_t (SubCellInst_SboxInst_11_n5), .Z0_f (new_AGEMA_signal_1496), .Z1_t (new_AGEMA_signal_1497), .Z1_f (new_AGEMA_signal_1498) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_U9 ( .A0_t (Output_s0_t[23]), .A0_f (Output_s0_f[23]), .A1_t (Output_s1_t[23]), .A1_f (Output_s1_f[23]), .B0_t (Output_s0_t[20]), .B0_f (Output_s0_f[20]), .B1_t (Output_s1_t[20]), .B1_f (Output_s1_f[20]), .Z0_t (SubCellInst_SboxInst_11_n10), .Z0_f (new_AGEMA_signal_1499), .Z1_t (new_AGEMA_signal_1500), .Z1_f (new_AGEMA_signal_1501) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_U8 ( .A0_t (SubCellInst_SboxInst_11_n8), .A0_f (new_AGEMA_signal_1505), .A1_t (new_AGEMA_signal_1506), .A1_f (new_AGEMA_signal_1507), .B0_t (SubCellInst_SboxInst_11_n3), .B0_f (new_AGEMA_signal_2787), .B1_t (new_AGEMA_signal_2788), .B1_f (new_AGEMA_signal_2789), .Z0_t (Feedback[44]), .Z0_f (new_AGEMA_signal_3292), .Z1_t (new_AGEMA_signal_3293), .Z1_f (new_AGEMA_signal_3294) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_U7 ( .A0_t (Output_s0_t[21]), .A0_f (Output_s0_f[21]), .A1_t (Output_s1_t[21]), .A1_f (Output_s1_f[21]), .B0_t (SubCellInst_SboxInst_11_n2), .B0_f (new_AGEMA_signal_2388), .B1_t (new_AGEMA_signal_2389), .B1_f (new_AGEMA_signal_2390), .Z0_t (SubCellInst_SboxInst_11_n3), .Z0_f (new_AGEMA_signal_2787), .Z1_t (new_AGEMA_signal_2788), .Z1_f (new_AGEMA_signal_2789) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_U6 ( .A0_t (Output_s0_t[20]), .A0_f (Output_s0_f[20]), .A1_t (Output_s1_t[20]), .A1_f (Output_s1_f[20]), .B0_t (SubCellInst_SboxInst_11_n1), .B0_f (new_AGEMA_signal_1502), .B1_t (new_AGEMA_signal_1503), .B1_f (new_AGEMA_signal_1504), .Z0_t (SubCellInst_SboxInst_11_n2), .Z0_f (new_AGEMA_signal_2388), .Z1_t (new_AGEMA_signal_2389), .Z1_f (new_AGEMA_signal_2390) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_U5 ( .A0_t (Output_s0_t[22]), .A0_f (Output_s0_f[22]), .A1_t (Output_s1_t[22]), .A1_f (Output_s1_f[22]), .B0_t (Output_s0_t[23]), .B0_f (Output_s0_f[23]), .B1_t (Output_s1_t[23]), .B1_f (Output_s1_f[23]), .Z0_t (SubCellInst_SboxInst_11_n1), .Z0_f (new_AGEMA_signal_1502), .Z1_t (new_AGEMA_signal_1503), .Z1_f (new_AGEMA_signal_1504) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_U3 ( .A0_t (Output_s0_t[22]), .A0_f (Output_s0_f[22]), .A1_t (Output_s1_t[22]), .A1_f (Output_s1_f[22]), .B0_t (Output_s0_t[23]), .B0_f (Output_s0_f[23]), .B1_t (Output_s1_t[23]), .B1_f (Output_s1_f[23]), .Z0_t (SubCellInst_SboxInst_11_n8), .Z0_f (new_AGEMA_signal_1505), .Z1_t (new_AGEMA_signal_1506), .Z1_f (new_AGEMA_signal_1507) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U19 ( .A0_t (SubCellInst_SboxInst_12_n15), .A0_f (new_AGEMA_signal_1517), .A1_t (new_AGEMA_signal_1518), .A1_f (new_AGEMA_signal_1519), .B0_t (SubCellInst_SboxInst_12_n14), .B0_f (new_AGEMA_signal_2391), .B1_t (new_AGEMA_signal_2392), .B1_f (new_AGEMA_signal_2393), .Z0_t (Feedback[49]), .Z0_f (new_AGEMA_signal_2790), .Z1_t (new_AGEMA_signal_2791), .Z1_f (new_AGEMA_signal_2792) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U18 ( .A0_t (Output_s0_t[4]), .A0_f (Output_s0_f[4]), .A1_t (Output_s1_t[4]), .A1_f (Output_s1_f[4]), .B0_t (SubCellInst_SboxInst_12_n13), .B0_f (new_AGEMA_signal_1514), .B1_t (new_AGEMA_signal_1515), .B1_f (new_AGEMA_signal_1516), .Z0_t (SubCellInst_SboxInst_12_n14), .Z0_f (new_AGEMA_signal_2391), .Z1_t (new_AGEMA_signal_2392), .Z1_f (new_AGEMA_signal_2393) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U17 ( .A0_t (Output_s0_t[7]), .A0_f (Output_s0_f[7]), .A1_t (Output_s1_t[7]), .A1_f (Output_s1_f[7]), .B0_t (Output_s0_t[6]), .B0_f (Output_s0_f[6]), .B1_t (Output_s1_t[6]), .B1_f (Output_s1_f[6]), .Z0_t (SubCellInst_SboxInst_12_n13), .Z0_f (new_AGEMA_signal_1514), .Z1_t (new_AGEMA_signal_1515), .Z1_f (new_AGEMA_signal_1516) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U16 ( .A0_t (Output_s0_t[6]), .A0_f (Output_s0_f[6]), .A1_t (Output_s1_t[6]), .A1_f (Output_s1_f[6]), .B0_t (Output_s0_t[7]), .B0_f (Output_s0_f[7]), .B1_t (Output_s1_t[7]), .B1_f (Output_s1_f[7]), .Z0_t (SubCellInst_SboxInst_12_n15), .Z0_f (new_AGEMA_signal_1517), .Z1_t (new_AGEMA_signal_1518), .Z1_f (new_AGEMA_signal_1519) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U15 ( .A0_t (SubCellInst_SboxInst_12_n10), .A0_f (new_AGEMA_signal_1526), .A1_t (new_AGEMA_signal_1527), .A1_f (new_AGEMA_signal_1528), .B0_t (SubCellInst_SboxInst_12_n9), .B0_f (new_AGEMA_signal_2397), .B1_t (new_AGEMA_signal_2398), .B1_f (new_AGEMA_signal_2399), .Z0_t (Feedback[51]), .Z0_f (new_AGEMA_signal_2793), .Z1_t (new_AGEMA_signal_2794), .Z1_f (new_AGEMA_signal_2795) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U14 ( .A0_t (SubCellInst_SboxInst_12_n8), .A0_f (new_AGEMA_signal_1532), .A1_t (new_AGEMA_signal_1533), .A1_f (new_AGEMA_signal_1534), .B0_t (Output_s0_t[5]), .B0_f (Output_s0_f[5]), .B1_t (Output_s1_t[5]), .B1_f (Output_s1_f[5]), .Z0_t (SubCellInst_SboxInst_12_n9), .Z0_f (new_AGEMA_signal_2397), .Z1_t (new_AGEMA_signal_2398), .Z1_f (new_AGEMA_signal_2399) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U13 ( .A0_t (SubCellInst_SboxInst_12_n10), .A0_f (new_AGEMA_signal_1526), .A1_t (new_AGEMA_signal_1527), .A1_f (new_AGEMA_signal_1528), .B0_t (SubCellInst_SboxInst_12_n7), .B0_f (new_AGEMA_signal_2796), .B1_t (new_AGEMA_signal_2797), .B1_f (new_AGEMA_signal_2798), .Z0_t (Feedback[50]), .Z0_f (new_AGEMA_signal_3295), .Z1_t (new_AGEMA_signal_3296), .Z1_f (new_AGEMA_signal_3297) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U12 ( .A0_t (SubCellInst_SboxInst_12_n6), .A0_f (new_AGEMA_signal_2400), .A1_t (new_AGEMA_signal_2401), .A1_f (new_AGEMA_signal_2402), .B0_t (Output_s0_t[5]), .B0_f (Output_s0_f[5]), .B1_t (Output_s1_t[5]), .B1_f (Output_s1_f[5]), .Z0_t (SubCellInst_SboxInst_12_n7), .Z0_f (new_AGEMA_signal_2796), .Z1_t (new_AGEMA_signal_2797), .Z1_f (new_AGEMA_signal_2798) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U11 ( .A0_t (SubCellInst_SboxInst_12_n5), .A0_f (new_AGEMA_signal_1523), .A1_t (new_AGEMA_signal_1524), .A1_f (new_AGEMA_signal_1525), .B0_t (Output_s0_t[6]), .B0_f (Output_s0_f[6]), .B1_t (Output_s1_t[6]), .B1_f (Output_s1_f[6]), .Z0_t (SubCellInst_SboxInst_12_n6), .Z0_f (new_AGEMA_signal_2400), .Z1_t (new_AGEMA_signal_2401), .Z1_f (new_AGEMA_signal_2402) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U10 ( .A0_t (Output_s0_t[4]), .A0_f (Output_s0_f[4]), .A1_t (Output_s1_t[4]), .A1_f (Output_s1_f[4]), .B0_t (Output_s0_t[7]), .B0_f (Output_s0_f[7]), .B1_t (Output_s1_t[7]), .B1_f (Output_s1_f[7]), .Z0_t (SubCellInst_SboxInst_12_n5), .Z0_f (new_AGEMA_signal_1523), .Z1_t (new_AGEMA_signal_1524), .Z1_f (new_AGEMA_signal_1525) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_U9 ( .A0_t (Output_s0_t[7]), .A0_f (Output_s0_f[7]), .A1_t (Output_s1_t[7]), .A1_f (Output_s1_f[7]), .B0_t (Output_s0_t[4]), .B0_f (Output_s0_f[4]), .B1_t (Output_s1_t[4]), .B1_f (Output_s1_f[4]), .Z0_t (SubCellInst_SboxInst_12_n10), .Z0_f (new_AGEMA_signal_1526), .Z1_t (new_AGEMA_signal_1527), .Z1_f (new_AGEMA_signal_1528) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_U8 ( .A0_t (SubCellInst_SboxInst_12_n8), .A0_f (new_AGEMA_signal_1532), .A1_t (new_AGEMA_signal_1533), .A1_f (new_AGEMA_signal_1534), .B0_t (SubCellInst_SboxInst_12_n3), .B0_f (new_AGEMA_signal_2799), .B1_t (new_AGEMA_signal_2800), .B1_f (new_AGEMA_signal_2801), .Z0_t (Feedback[48]), .Z0_f (new_AGEMA_signal_3298), .Z1_t (new_AGEMA_signal_3299), .Z1_f (new_AGEMA_signal_3300) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_U7 ( .A0_t (Output_s0_t[5]), .A0_f (Output_s0_f[5]), .A1_t (Output_s1_t[5]), .A1_f (Output_s1_f[5]), .B0_t (SubCellInst_SboxInst_12_n2), .B0_f (new_AGEMA_signal_2403), .B1_t (new_AGEMA_signal_2404), .B1_f (new_AGEMA_signal_2405), .Z0_t (SubCellInst_SboxInst_12_n3), .Z0_f (new_AGEMA_signal_2799), .Z1_t (new_AGEMA_signal_2800), .Z1_f (new_AGEMA_signal_2801) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_U6 ( .A0_t (Output_s0_t[4]), .A0_f (Output_s0_f[4]), .A1_t (Output_s1_t[4]), .A1_f (Output_s1_f[4]), .B0_t (SubCellInst_SboxInst_12_n1), .B0_f (new_AGEMA_signal_1529), .B1_t (new_AGEMA_signal_1530), .B1_f (new_AGEMA_signal_1531), .Z0_t (SubCellInst_SboxInst_12_n2), .Z0_f (new_AGEMA_signal_2403), .Z1_t (new_AGEMA_signal_2404), .Z1_f (new_AGEMA_signal_2405) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_U5 ( .A0_t (Output_s0_t[6]), .A0_f (Output_s0_f[6]), .A1_t (Output_s1_t[6]), .A1_f (Output_s1_f[6]), .B0_t (Output_s0_t[7]), .B0_f (Output_s0_f[7]), .B1_t (Output_s1_t[7]), .B1_f (Output_s1_f[7]), .Z0_t (SubCellInst_SboxInst_12_n1), .Z0_f (new_AGEMA_signal_1529), .Z1_t (new_AGEMA_signal_1530), .Z1_f (new_AGEMA_signal_1531) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_U3 ( .A0_t (Output_s0_t[6]), .A0_f (Output_s0_f[6]), .A1_t (Output_s1_t[6]), .A1_f (Output_s1_f[6]), .B0_t (Output_s0_t[7]), .B0_f (Output_s0_f[7]), .B1_t (Output_s1_t[7]), .B1_f (Output_s1_f[7]), .Z0_t (SubCellInst_SboxInst_12_n8), .Z0_f (new_AGEMA_signal_1532), .Z1_t (new_AGEMA_signal_1533), .Z1_f (new_AGEMA_signal_1534) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U19 ( .A0_t (SubCellInst_SboxInst_13_n15), .A0_f (new_AGEMA_signal_1544), .A1_t (new_AGEMA_signal_1545), .A1_f (new_AGEMA_signal_1546), .B0_t (SubCellInst_SboxInst_13_n14), .B0_f (new_AGEMA_signal_2406), .B1_t (new_AGEMA_signal_2407), .B1_f (new_AGEMA_signal_2408), .Z0_t (Feedback[53]), .Z0_f (new_AGEMA_signal_2802), .Z1_t (new_AGEMA_signal_2803), .Z1_f (new_AGEMA_signal_2804) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U18 ( .A0_t (Output_s0_t[8]), .A0_f (Output_s0_f[8]), .A1_t (Output_s1_t[8]), .A1_f (Output_s1_f[8]), .B0_t (SubCellInst_SboxInst_13_n13), .B0_f (new_AGEMA_signal_1541), .B1_t (new_AGEMA_signal_1542), .B1_f (new_AGEMA_signal_1543), .Z0_t (SubCellInst_SboxInst_13_n14), .Z0_f (new_AGEMA_signal_2406), .Z1_t (new_AGEMA_signal_2407), .Z1_f (new_AGEMA_signal_2408) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U17 ( .A0_t (Output_s0_t[11]), .A0_f (Output_s0_f[11]), .A1_t (Output_s1_t[11]), .A1_f (Output_s1_f[11]), .B0_t (Output_s0_t[10]), .B0_f (Output_s0_f[10]), .B1_t (Output_s1_t[10]), .B1_f (Output_s1_f[10]), .Z0_t (SubCellInst_SboxInst_13_n13), .Z0_f (new_AGEMA_signal_1541), .Z1_t (new_AGEMA_signal_1542), .Z1_f (new_AGEMA_signal_1543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U16 ( .A0_t (Output_s0_t[10]), .A0_f (Output_s0_f[10]), .A1_t (Output_s1_t[10]), .A1_f (Output_s1_f[10]), .B0_t (Output_s0_t[11]), .B0_f (Output_s0_f[11]), .B1_t (Output_s1_t[11]), .B1_f (Output_s1_f[11]), .Z0_t (SubCellInst_SboxInst_13_n15), .Z0_f (new_AGEMA_signal_1544), .Z1_t (new_AGEMA_signal_1545), .Z1_f (new_AGEMA_signal_1546) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U15 ( .A0_t (SubCellInst_SboxInst_13_n10), .A0_f (new_AGEMA_signal_1553), .A1_t (new_AGEMA_signal_1554), .A1_f (new_AGEMA_signal_1555), .B0_t (SubCellInst_SboxInst_13_n9), .B0_f (new_AGEMA_signal_2412), .B1_t (new_AGEMA_signal_2413), .B1_f (new_AGEMA_signal_2414), .Z0_t (Feedback[55]), .Z0_f (new_AGEMA_signal_2805), .Z1_t (new_AGEMA_signal_2806), .Z1_f (new_AGEMA_signal_2807) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U14 ( .A0_t (SubCellInst_SboxInst_13_n8), .A0_f (new_AGEMA_signal_1559), .A1_t (new_AGEMA_signal_1560), .A1_f (new_AGEMA_signal_1561), .B0_t (Output_s0_t[9]), .B0_f (Output_s0_f[9]), .B1_t (Output_s1_t[9]), .B1_f (Output_s1_f[9]), .Z0_t (SubCellInst_SboxInst_13_n9), .Z0_f (new_AGEMA_signal_2412), .Z1_t (new_AGEMA_signal_2413), .Z1_f (new_AGEMA_signal_2414) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U13 ( .A0_t (SubCellInst_SboxInst_13_n10), .A0_f (new_AGEMA_signal_1553), .A1_t (new_AGEMA_signal_1554), .A1_f (new_AGEMA_signal_1555), .B0_t (SubCellInst_SboxInst_13_n7), .B0_f (new_AGEMA_signal_2808), .B1_t (new_AGEMA_signal_2809), .B1_f (new_AGEMA_signal_2810), .Z0_t (Feedback[54]), .Z0_f (new_AGEMA_signal_3301), .Z1_t (new_AGEMA_signal_3302), .Z1_f (new_AGEMA_signal_3303) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U12 ( .A0_t (SubCellInst_SboxInst_13_n6), .A0_f (new_AGEMA_signal_2415), .A1_t (new_AGEMA_signal_2416), .A1_f (new_AGEMA_signal_2417), .B0_t (Output_s0_t[9]), .B0_f (Output_s0_f[9]), .B1_t (Output_s1_t[9]), .B1_f (Output_s1_f[9]), .Z0_t (SubCellInst_SboxInst_13_n7), .Z0_f (new_AGEMA_signal_2808), .Z1_t (new_AGEMA_signal_2809), .Z1_f (new_AGEMA_signal_2810) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U11 ( .A0_t (SubCellInst_SboxInst_13_n5), .A0_f (new_AGEMA_signal_1550), .A1_t (new_AGEMA_signal_1551), .A1_f (new_AGEMA_signal_1552), .B0_t (Output_s0_t[10]), .B0_f (Output_s0_f[10]), .B1_t (Output_s1_t[10]), .B1_f (Output_s1_f[10]), .Z0_t (SubCellInst_SboxInst_13_n6), .Z0_f (new_AGEMA_signal_2415), .Z1_t (new_AGEMA_signal_2416), .Z1_f (new_AGEMA_signal_2417) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U10 ( .A0_t (Output_s0_t[8]), .A0_f (Output_s0_f[8]), .A1_t (Output_s1_t[8]), .A1_f (Output_s1_f[8]), .B0_t (Output_s0_t[11]), .B0_f (Output_s0_f[11]), .B1_t (Output_s1_t[11]), .B1_f (Output_s1_f[11]), .Z0_t (SubCellInst_SboxInst_13_n5), .Z0_f (new_AGEMA_signal_1550), .Z1_t (new_AGEMA_signal_1551), .Z1_f (new_AGEMA_signal_1552) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_U9 ( .A0_t (Output_s0_t[11]), .A0_f (Output_s0_f[11]), .A1_t (Output_s1_t[11]), .A1_f (Output_s1_f[11]), .B0_t (Output_s0_t[8]), .B0_f (Output_s0_f[8]), .B1_t (Output_s1_t[8]), .B1_f (Output_s1_f[8]), .Z0_t (SubCellInst_SboxInst_13_n10), .Z0_f (new_AGEMA_signal_1553), .Z1_t (new_AGEMA_signal_1554), .Z1_f (new_AGEMA_signal_1555) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_U8 ( .A0_t (SubCellInst_SboxInst_13_n8), .A0_f (new_AGEMA_signal_1559), .A1_t (new_AGEMA_signal_1560), .A1_f (new_AGEMA_signal_1561), .B0_t (SubCellInst_SboxInst_13_n3), .B0_f (new_AGEMA_signal_2811), .B1_t (new_AGEMA_signal_2812), .B1_f (new_AGEMA_signal_2813), .Z0_t (Feedback[52]), .Z0_f (new_AGEMA_signal_3304), .Z1_t (new_AGEMA_signal_3305), .Z1_f (new_AGEMA_signal_3306) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_U7 ( .A0_t (Output_s0_t[9]), .A0_f (Output_s0_f[9]), .A1_t (Output_s1_t[9]), .A1_f (Output_s1_f[9]), .B0_t (SubCellInst_SboxInst_13_n2), .B0_f (new_AGEMA_signal_2418), .B1_t (new_AGEMA_signal_2419), .B1_f (new_AGEMA_signal_2420), .Z0_t (SubCellInst_SboxInst_13_n3), .Z0_f (new_AGEMA_signal_2811), .Z1_t (new_AGEMA_signal_2812), .Z1_f (new_AGEMA_signal_2813) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_U6 ( .A0_t (Output_s0_t[8]), .A0_f (Output_s0_f[8]), .A1_t (Output_s1_t[8]), .A1_f (Output_s1_f[8]), .B0_t (SubCellInst_SboxInst_13_n1), .B0_f (new_AGEMA_signal_1556), .B1_t (new_AGEMA_signal_1557), .B1_f (new_AGEMA_signal_1558), .Z0_t (SubCellInst_SboxInst_13_n2), .Z0_f (new_AGEMA_signal_2418), .Z1_t (new_AGEMA_signal_2419), .Z1_f (new_AGEMA_signal_2420) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_U5 ( .A0_t (Output_s0_t[10]), .A0_f (Output_s0_f[10]), .A1_t (Output_s1_t[10]), .A1_f (Output_s1_f[10]), .B0_t (Output_s0_t[11]), .B0_f (Output_s0_f[11]), .B1_t (Output_s1_t[11]), .B1_f (Output_s1_f[11]), .Z0_t (SubCellInst_SboxInst_13_n1), .Z0_f (new_AGEMA_signal_1556), .Z1_t (new_AGEMA_signal_1557), .Z1_f (new_AGEMA_signal_1558) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_U3 ( .A0_t (Output_s0_t[10]), .A0_f (Output_s0_f[10]), .A1_t (Output_s1_t[10]), .A1_f (Output_s1_f[10]), .B0_t (Output_s0_t[11]), .B0_f (Output_s0_f[11]), .B1_t (Output_s1_t[11]), .B1_f (Output_s1_f[11]), .Z0_t (SubCellInst_SboxInst_13_n8), .Z0_f (new_AGEMA_signal_1559), .Z1_t (new_AGEMA_signal_1560), .Z1_f (new_AGEMA_signal_1561) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U19 ( .A0_t (SubCellInst_SboxInst_14_n15), .A0_f (new_AGEMA_signal_1571), .A1_t (new_AGEMA_signal_1572), .A1_f (new_AGEMA_signal_1573), .B0_t (SubCellInst_SboxInst_14_n14), .B0_f (new_AGEMA_signal_2421), .B1_t (new_AGEMA_signal_2422), .B1_f (new_AGEMA_signal_2423), .Z0_t (Feedback[57]), .Z0_f (new_AGEMA_signal_2814), .Z1_t (new_AGEMA_signal_2815), .Z1_f (new_AGEMA_signal_2816) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U18 ( .A0_t (Output_s0_t[12]), .A0_f (Output_s0_f[12]), .A1_t (Output_s1_t[12]), .A1_f (Output_s1_f[12]), .B0_t (SubCellInst_SboxInst_14_n13), .B0_f (new_AGEMA_signal_1568), .B1_t (new_AGEMA_signal_1569), .B1_f (new_AGEMA_signal_1570), .Z0_t (SubCellInst_SboxInst_14_n14), .Z0_f (new_AGEMA_signal_2421), .Z1_t (new_AGEMA_signal_2422), .Z1_f (new_AGEMA_signal_2423) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U17 ( .A0_t (Output_s0_t[15]), .A0_f (Output_s0_f[15]), .A1_t (Output_s1_t[15]), .A1_f (Output_s1_f[15]), .B0_t (Output_s0_t[14]), .B0_f (Output_s0_f[14]), .B1_t (Output_s1_t[14]), .B1_f (Output_s1_f[14]), .Z0_t (SubCellInst_SboxInst_14_n13), .Z0_f (new_AGEMA_signal_1568), .Z1_t (new_AGEMA_signal_1569), .Z1_f (new_AGEMA_signal_1570) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U16 ( .A0_t (Output_s0_t[14]), .A0_f (Output_s0_f[14]), .A1_t (Output_s1_t[14]), .A1_f (Output_s1_f[14]), .B0_t (Output_s0_t[15]), .B0_f (Output_s0_f[15]), .B1_t (Output_s1_t[15]), .B1_f (Output_s1_f[15]), .Z0_t (SubCellInst_SboxInst_14_n15), .Z0_f (new_AGEMA_signal_1571), .Z1_t (new_AGEMA_signal_1572), .Z1_f (new_AGEMA_signal_1573) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U15 ( .A0_t (SubCellInst_SboxInst_14_n10), .A0_f (new_AGEMA_signal_1580), .A1_t (new_AGEMA_signal_1581), .A1_f (new_AGEMA_signal_1582), .B0_t (SubCellInst_SboxInst_14_n9), .B0_f (new_AGEMA_signal_2427), .B1_t (new_AGEMA_signal_2428), .B1_f (new_AGEMA_signal_2429), .Z0_t (Feedback[59]), .Z0_f (new_AGEMA_signal_2817), .Z1_t (new_AGEMA_signal_2818), .Z1_f (new_AGEMA_signal_2819) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U14 ( .A0_t (SubCellInst_SboxInst_14_n8), .A0_f (new_AGEMA_signal_1586), .A1_t (new_AGEMA_signal_1587), .A1_f (new_AGEMA_signal_1588), .B0_t (Output_s0_t[13]), .B0_f (Output_s0_f[13]), .B1_t (Output_s1_t[13]), .B1_f (Output_s1_f[13]), .Z0_t (SubCellInst_SboxInst_14_n9), .Z0_f (new_AGEMA_signal_2427), .Z1_t (new_AGEMA_signal_2428), .Z1_f (new_AGEMA_signal_2429) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U13 ( .A0_t (SubCellInst_SboxInst_14_n10), .A0_f (new_AGEMA_signal_1580), .A1_t (new_AGEMA_signal_1581), .A1_f (new_AGEMA_signal_1582), .B0_t (SubCellInst_SboxInst_14_n7), .B0_f (new_AGEMA_signal_2820), .B1_t (new_AGEMA_signal_2821), .B1_f (new_AGEMA_signal_2822), .Z0_t (Feedback[58]), .Z0_f (new_AGEMA_signal_3307), .Z1_t (new_AGEMA_signal_3308), .Z1_f (new_AGEMA_signal_3309) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U12 ( .A0_t (SubCellInst_SboxInst_14_n6), .A0_f (new_AGEMA_signal_2430), .A1_t (new_AGEMA_signal_2431), .A1_f (new_AGEMA_signal_2432), .B0_t (Output_s0_t[13]), .B0_f (Output_s0_f[13]), .B1_t (Output_s1_t[13]), .B1_f (Output_s1_f[13]), .Z0_t (SubCellInst_SboxInst_14_n7), .Z0_f (new_AGEMA_signal_2820), .Z1_t (new_AGEMA_signal_2821), .Z1_f (new_AGEMA_signal_2822) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U11 ( .A0_t (SubCellInst_SboxInst_14_n5), .A0_f (new_AGEMA_signal_1577), .A1_t (new_AGEMA_signal_1578), .A1_f (new_AGEMA_signal_1579), .B0_t (Output_s0_t[14]), .B0_f (Output_s0_f[14]), .B1_t (Output_s1_t[14]), .B1_f (Output_s1_f[14]), .Z0_t (SubCellInst_SboxInst_14_n6), .Z0_f (new_AGEMA_signal_2430), .Z1_t (new_AGEMA_signal_2431), .Z1_f (new_AGEMA_signal_2432) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U10 ( .A0_t (Output_s0_t[12]), .A0_f (Output_s0_f[12]), .A1_t (Output_s1_t[12]), .A1_f (Output_s1_f[12]), .B0_t (Output_s0_t[15]), .B0_f (Output_s0_f[15]), .B1_t (Output_s1_t[15]), .B1_f (Output_s1_f[15]), .Z0_t (SubCellInst_SboxInst_14_n5), .Z0_f (new_AGEMA_signal_1577), .Z1_t (new_AGEMA_signal_1578), .Z1_f (new_AGEMA_signal_1579) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_U9 ( .A0_t (Output_s0_t[15]), .A0_f (Output_s0_f[15]), .A1_t (Output_s1_t[15]), .A1_f (Output_s1_f[15]), .B0_t (Output_s0_t[12]), .B0_f (Output_s0_f[12]), .B1_t (Output_s1_t[12]), .B1_f (Output_s1_f[12]), .Z0_t (SubCellInst_SboxInst_14_n10), .Z0_f (new_AGEMA_signal_1580), .Z1_t (new_AGEMA_signal_1581), .Z1_f (new_AGEMA_signal_1582) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_U8 ( .A0_t (SubCellInst_SboxInst_14_n8), .A0_f (new_AGEMA_signal_1586), .A1_t (new_AGEMA_signal_1587), .A1_f (new_AGEMA_signal_1588), .B0_t (SubCellInst_SboxInst_14_n3), .B0_f (new_AGEMA_signal_2823), .B1_t (new_AGEMA_signal_2824), .B1_f (new_AGEMA_signal_2825), .Z0_t (Feedback[56]), .Z0_f (new_AGEMA_signal_3310), .Z1_t (new_AGEMA_signal_3311), .Z1_f (new_AGEMA_signal_3312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_U7 ( .A0_t (Output_s0_t[13]), .A0_f (Output_s0_f[13]), .A1_t (Output_s1_t[13]), .A1_f (Output_s1_f[13]), .B0_t (SubCellInst_SboxInst_14_n2), .B0_f (new_AGEMA_signal_2433), .B1_t (new_AGEMA_signal_2434), .B1_f (new_AGEMA_signal_2435), .Z0_t (SubCellInst_SboxInst_14_n3), .Z0_f (new_AGEMA_signal_2823), .Z1_t (new_AGEMA_signal_2824), .Z1_f (new_AGEMA_signal_2825) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_U6 ( .A0_t (Output_s0_t[12]), .A0_f (Output_s0_f[12]), .A1_t (Output_s1_t[12]), .A1_f (Output_s1_f[12]), .B0_t (SubCellInst_SboxInst_14_n1), .B0_f (new_AGEMA_signal_1583), .B1_t (new_AGEMA_signal_1584), .B1_f (new_AGEMA_signal_1585), .Z0_t (SubCellInst_SboxInst_14_n2), .Z0_f (new_AGEMA_signal_2433), .Z1_t (new_AGEMA_signal_2434), .Z1_f (new_AGEMA_signal_2435) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_U5 ( .A0_t (Output_s0_t[14]), .A0_f (Output_s0_f[14]), .A1_t (Output_s1_t[14]), .A1_f (Output_s1_f[14]), .B0_t (Output_s0_t[15]), .B0_f (Output_s0_f[15]), .B1_t (Output_s1_t[15]), .B1_f (Output_s1_f[15]), .Z0_t (SubCellInst_SboxInst_14_n1), .Z0_f (new_AGEMA_signal_1583), .Z1_t (new_AGEMA_signal_1584), .Z1_f (new_AGEMA_signal_1585) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_U3 ( .A0_t (Output_s0_t[14]), .A0_f (Output_s0_f[14]), .A1_t (Output_s1_t[14]), .A1_f (Output_s1_f[14]), .B0_t (Output_s0_t[15]), .B0_f (Output_s0_f[15]), .B1_t (Output_s1_t[15]), .B1_f (Output_s1_f[15]), .Z0_t (SubCellInst_SboxInst_14_n8), .Z0_f (new_AGEMA_signal_1586), .Z1_t (new_AGEMA_signal_1587), .Z1_f (new_AGEMA_signal_1588) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U19 ( .A0_t (SubCellInst_SboxInst_15_n15), .A0_f (new_AGEMA_signal_1598), .A1_t (new_AGEMA_signal_1599), .A1_f (new_AGEMA_signal_1600), .B0_t (SubCellInst_SboxInst_15_n14), .B0_f (new_AGEMA_signal_2436), .B1_t (new_AGEMA_signal_2437), .B1_f (new_AGEMA_signal_2438), .Z0_t (Feedback[61]), .Z0_f (new_AGEMA_signal_2826), .Z1_t (new_AGEMA_signal_2827), .Z1_f (new_AGEMA_signal_2828) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U18 ( .A0_t (Output_s0_t[0]), .A0_f (Output_s0_f[0]), .A1_t (Output_s1_t[0]), .A1_f (Output_s1_f[0]), .B0_t (SubCellInst_SboxInst_15_n13), .B0_f (new_AGEMA_signal_1595), .B1_t (new_AGEMA_signal_1596), .B1_f (new_AGEMA_signal_1597), .Z0_t (SubCellInst_SboxInst_15_n14), .Z0_f (new_AGEMA_signal_2436), .Z1_t (new_AGEMA_signal_2437), .Z1_f (new_AGEMA_signal_2438) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U17 ( .A0_t (Output_s0_t[3]), .A0_f (Output_s0_f[3]), .A1_t (Output_s1_t[3]), .A1_f (Output_s1_f[3]), .B0_t (Output_s0_t[2]), .B0_f (Output_s0_f[2]), .B1_t (Output_s1_t[2]), .B1_f (Output_s1_f[2]), .Z0_t (SubCellInst_SboxInst_15_n13), .Z0_f (new_AGEMA_signal_1595), .Z1_t (new_AGEMA_signal_1596), .Z1_f (new_AGEMA_signal_1597) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U16 ( .A0_t (Output_s0_t[2]), .A0_f (Output_s0_f[2]), .A1_t (Output_s1_t[2]), .A1_f (Output_s1_f[2]), .B0_t (Output_s0_t[3]), .B0_f (Output_s0_f[3]), .B1_t (Output_s1_t[3]), .B1_f (Output_s1_f[3]), .Z0_t (SubCellInst_SboxInst_15_n15), .Z0_f (new_AGEMA_signal_1598), .Z1_t (new_AGEMA_signal_1599), .Z1_f (new_AGEMA_signal_1600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U15 ( .A0_t (SubCellInst_SboxInst_15_n10), .A0_f (new_AGEMA_signal_1607), .A1_t (new_AGEMA_signal_1608), .A1_f (new_AGEMA_signal_1609), .B0_t (SubCellInst_SboxInst_15_n9), .B0_f (new_AGEMA_signal_2442), .B1_t (new_AGEMA_signal_2443), .B1_f (new_AGEMA_signal_2444), .Z0_t (Feedback[63]), .Z0_f (new_AGEMA_signal_2829), .Z1_t (new_AGEMA_signal_2830), .Z1_f (new_AGEMA_signal_2831) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U14 ( .A0_t (SubCellInst_SboxInst_15_n8), .A0_f (new_AGEMA_signal_1613), .A1_t (new_AGEMA_signal_1614), .A1_f (new_AGEMA_signal_1615), .B0_t (Output_s0_t[1]), .B0_f (Output_s0_f[1]), .B1_t (Output_s1_t[1]), .B1_f (Output_s1_f[1]), .Z0_t (SubCellInst_SboxInst_15_n9), .Z0_f (new_AGEMA_signal_2442), .Z1_t (new_AGEMA_signal_2443), .Z1_f (new_AGEMA_signal_2444) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U13 ( .A0_t (SubCellInst_SboxInst_15_n10), .A0_f (new_AGEMA_signal_1607), .A1_t (new_AGEMA_signal_1608), .A1_f (new_AGEMA_signal_1609), .B0_t (SubCellInst_SboxInst_15_n7), .B0_f (new_AGEMA_signal_2832), .B1_t (new_AGEMA_signal_2833), .B1_f (new_AGEMA_signal_2834), .Z0_t (Feedback[62]), .Z0_f (new_AGEMA_signal_3313), .Z1_t (new_AGEMA_signal_3314), .Z1_f (new_AGEMA_signal_3315) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U12 ( .A0_t (SubCellInst_SboxInst_15_n6), .A0_f (new_AGEMA_signal_2445), .A1_t (new_AGEMA_signal_2446), .A1_f (new_AGEMA_signal_2447), .B0_t (Output_s0_t[1]), .B0_f (Output_s0_f[1]), .B1_t (Output_s1_t[1]), .B1_f (Output_s1_f[1]), .Z0_t (SubCellInst_SboxInst_15_n7), .Z0_f (new_AGEMA_signal_2832), .Z1_t (new_AGEMA_signal_2833), .Z1_f (new_AGEMA_signal_2834) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U11 ( .A0_t (SubCellInst_SboxInst_15_n5), .A0_f (new_AGEMA_signal_1604), .A1_t (new_AGEMA_signal_1605), .A1_f (new_AGEMA_signal_1606), .B0_t (Output_s0_t[2]), .B0_f (Output_s0_f[2]), .B1_t (Output_s1_t[2]), .B1_f (Output_s1_f[2]), .Z0_t (SubCellInst_SboxInst_15_n6), .Z0_f (new_AGEMA_signal_2445), .Z1_t (new_AGEMA_signal_2446), .Z1_f (new_AGEMA_signal_2447) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U10 ( .A0_t (Output_s0_t[0]), .A0_f (Output_s0_f[0]), .A1_t (Output_s1_t[0]), .A1_f (Output_s1_f[0]), .B0_t (Output_s0_t[3]), .B0_f (Output_s0_f[3]), .B1_t (Output_s1_t[3]), .B1_f (Output_s1_f[3]), .Z0_t (SubCellInst_SboxInst_15_n5), .Z0_f (new_AGEMA_signal_1604), .Z1_t (new_AGEMA_signal_1605), .Z1_f (new_AGEMA_signal_1606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_U9 ( .A0_t (Output_s0_t[3]), .A0_f (Output_s0_f[3]), .A1_t (Output_s1_t[3]), .A1_f (Output_s1_f[3]), .B0_t (Output_s0_t[0]), .B0_f (Output_s0_f[0]), .B1_t (Output_s1_t[0]), .B1_f (Output_s1_f[0]), .Z0_t (SubCellInst_SboxInst_15_n10), .Z0_f (new_AGEMA_signal_1607), .Z1_t (new_AGEMA_signal_1608), .Z1_f (new_AGEMA_signal_1609) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_U8 ( .A0_t (SubCellInst_SboxInst_15_n8), .A0_f (new_AGEMA_signal_1613), .A1_t (new_AGEMA_signal_1614), .A1_f (new_AGEMA_signal_1615), .B0_t (SubCellInst_SboxInst_15_n3), .B0_f (new_AGEMA_signal_2835), .B1_t (new_AGEMA_signal_2836), .B1_f (new_AGEMA_signal_2837), .Z0_t (Feedback[60]), .Z0_f (new_AGEMA_signal_3316), .Z1_t (new_AGEMA_signal_3317), .Z1_f (new_AGEMA_signal_3318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_U7 ( .A0_t (Output_s0_t[1]), .A0_f (Output_s0_f[1]), .A1_t (Output_s1_t[1]), .A1_f (Output_s1_f[1]), .B0_t (SubCellInst_SboxInst_15_n2), .B0_f (new_AGEMA_signal_2448), .B1_t (new_AGEMA_signal_2449), .B1_f (new_AGEMA_signal_2450), .Z0_t (SubCellInst_SboxInst_15_n3), .Z0_f (new_AGEMA_signal_2835), .Z1_t (new_AGEMA_signal_2836), .Z1_f (new_AGEMA_signal_2837) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_U6 ( .A0_t (Output_s0_t[0]), .A0_f (Output_s0_f[0]), .A1_t (Output_s1_t[0]), .A1_f (Output_s1_f[0]), .B0_t (SubCellInst_SboxInst_15_n1), .B0_f (new_AGEMA_signal_1610), .B1_t (new_AGEMA_signal_1611), .B1_f (new_AGEMA_signal_1612), .Z0_t (SubCellInst_SboxInst_15_n2), .Z0_f (new_AGEMA_signal_2448), .Z1_t (new_AGEMA_signal_2449), .Z1_f (new_AGEMA_signal_2450) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_U5 ( .A0_t (Output_s0_t[2]), .A0_f (Output_s0_f[2]), .A1_t (Output_s1_t[2]), .A1_f (Output_s1_f[2]), .B0_t (Output_s0_t[3]), .B0_f (Output_s0_f[3]), .B1_t (Output_s1_t[3]), .B1_f (Output_s1_f[3]), .Z0_t (SubCellInst_SboxInst_15_n1), .Z0_f (new_AGEMA_signal_1610), .Z1_t (new_AGEMA_signal_1611), .Z1_f (new_AGEMA_signal_1612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_U3 ( .A0_t (Output_s0_t[2]), .A0_f (Output_s0_f[2]), .A1_t (Output_s1_t[2]), .A1_f (Output_s1_f[2]), .B0_t (Output_s0_t[3]), .B0_f (Output_s0_f[3]), .B1_t (Output_s1_t[3]), .B1_f (Output_s1_f[3]), .Z0_t (SubCellInst_SboxInst_15_n8), .Z0_f (new_AGEMA_signal_1613), .Z1_t (new_AGEMA_signal_1614), .Z1_f (new_AGEMA_signal_1615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_0_U1_XOR1_U1 ( .A0_t (Key_s0_t[64]), .A0_f (Key_s0_f[64]), .A1_t (Key_s1_t[64]), .A1_f (Key_s1_f[64]), .B0_t (Key_s0_t[0]), .B0_f (Key_s0_f[0]), .B1_t (Key_s1_t[0]), .B1_f (Key_s1_f[0]), .Z0_t (KeyMUX_MUXInst_0_U1_X), .Z0_f (new_AGEMA_signal_1622), .Z1_t (new_AGEMA_signal_1623), .Z1_f (new_AGEMA_signal_1624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_0_U1_X), .B0_f (new_AGEMA_signal_1622), .B1_t (new_AGEMA_signal_1623), .B1_f (new_AGEMA_signal_1624), .Z0_t (KeyMUX_MUXInst_0_U1_Y), .Z0_f (new_AGEMA_signal_2451), .Z1_t (new_AGEMA_signal_2452), .Z1_f (new_AGEMA_signal_2453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_0_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_0_U1_Y), .A0_f (new_AGEMA_signal_2451), .A1_t (new_AGEMA_signal_2452), .A1_f (new_AGEMA_signal_2453), .B0_t (Key_s0_t[64]), .B0_f (Key_s0_f[64]), .B1_t (Key_s1_t[64]), .B1_f (Key_s1_f[64]), .Z0_t (SelectedKey[0]), .Z0_f (new_AGEMA_signal_2838), .Z1_t (new_AGEMA_signal_2839), .Z1_f (new_AGEMA_signal_2840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_1_U1_XOR1_U1 ( .A0_t (Key_s0_t[65]), .A0_f (Key_s0_f[65]), .A1_t (Key_s1_t[65]), .A1_f (Key_s1_f[65]), .B0_t (Key_s0_t[1]), .B0_f (Key_s0_f[1]), .B1_t (Key_s1_t[1]), .B1_f (Key_s1_f[1]), .Z0_t (KeyMUX_MUXInst_1_U1_X), .Z0_f (new_AGEMA_signal_1631), .Z1_t (new_AGEMA_signal_1632), .Z1_f (new_AGEMA_signal_1633) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_1_U1_X), .B0_f (new_AGEMA_signal_1631), .B1_t (new_AGEMA_signal_1632), .B1_f (new_AGEMA_signal_1633), .Z0_t (KeyMUX_MUXInst_1_U1_Y), .Z0_f (new_AGEMA_signal_2454), .Z1_t (new_AGEMA_signal_2455), .Z1_f (new_AGEMA_signal_2456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_1_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_1_U1_Y), .A0_f (new_AGEMA_signal_2454), .A1_t (new_AGEMA_signal_2455), .A1_f (new_AGEMA_signal_2456), .B0_t (Key_s0_t[65]), .B0_f (Key_s0_f[65]), .B1_t (Key_s1_t[65]), .B1_f (Key_s1_f[65]), .Z0_t (SelectedKey[1]), .Z0_f (new_AGEMA_signal_2841), .Z1_t (new_AGEMA_signal_2842), .Z1_f (new_AGEMA_signal_2843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_2_U1_XOR1_U1 ( .A0_t (Key_s0_t[66]), .A0_f (Key_s0_f[66]), .A1_t (Key_s1_t[66]), .A1_f (Key_s1_f[66]), .B0_t (Key_s0_t[2]), .B0_f (Key_s0_f[2]), .B1_t (Key_s1_t[2]), .B1_f (Key_s1_f[2]), .Z0_t (KeyMUX_MUXInst_2_U1_X), .Z0_f (new_AGEMA_signal_1640), .Z1_t (new_AGEMA_signal_1641), .Z1_f (new_AGEMA_signal_1642) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_2_U1_X), .B0_f (new_AGEMA_signal_1640), .B1_t (new_AGEMA_signal_1641), .B1_f (new_AGEMA_signal_1642), .Z0_t (KeyMUX_MUXInst_2_U1_Y), .Z0_f (new_AGEMA_signal_2457), .Z1_t (new_AGEMA_signal_2458), .Z1_f (new_AGEMA_signal_2459) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_2_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_2_U1_Y), .A0_f (new_AGEMA_signal_2457), .A1_t (new_AGEMA_signal_2458), .A1_f (new_AGEMA_signal_2459), .B0_t (Key_s0_t[66]), .B0_f (Key_s0_f[66]), .B1_t (Key_s1_t[66]), .B1_f (Key_s1_f[66]), .Z0_t (SelectedKey[2]), .Z0_f (new_AGEMA_signal_2844), .Z1_t (new_AGEMA_signal_2845), .Z1_f (new_AGEMA_signal_2846) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_3_U1_XOR1_U1 ( .A0_t (Key_s0_t[67]), .A0_f (Key_s0_f[67]), .A1_t (Key_s1_t[67]), .A1_f (Key_s1_f[67]), .B0_t (Key_s0_t[3]), .B0_f (Key_s0_f[3]), .B1_t (Key_s1_t[3]), .B1_f (Key_s1_f[3]), .Z0_t (KeyMUX_MUXInst_3_U1_X), .Z0_f (new_AGEMA_signal_1649), .Z1_t (new_AGEMA_signal_1650), .Z1_f (new_AGEMA_signal_1651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_3_U1_X), .B0_f (new_AGEMA_signal_1649), .B1_t (new_AGEMA_signal_1650), .B1_f (new_AGEMA_signal_1651), .Z0_t (KeyMUX_MUXInst_3_U1_Y), .Z0_f (new_AGEMA_signal_2460), .Z1_t (new_AGEMA_signal_2461), .Z1_f (new_AGEMA_signal_2462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_3_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_3_U1_Y), .A0_f (new_AGEMA_signal_2460), .A1_t (new_AGEMA_signal_2461), .A1_f (new_AGEMA_signal_2462), .B0_t (Key_s0_t[67]), .B0_f (Key_s0_f[67]), .B1_t (Key_s1_t[67]), .B1_f (Key_s1_f[67]), .Z0_t (SelectedKey[3]), .Z0_f (new_AGEMA_signal_2847), .Z1_t (new_AGEMA_signal_2848), .Z1_f (new_AGEMA_signal_2849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_4_U1_XOR1_U1 ( .A0_t (Key_s0_t[68]), .A0_f (Key_s0_f[68]), .A1_t (Key_s1_t[68]), .A1_f (Key_s1_f[68]), .B0_t (Key_s0_t[4]), .B0_f (Key_s0_f[4]), .B1_t (Key_s1_t[4]), .B1_f (Key_s1_f[4]), .Z0_t (KeyMUX_MUXInst_4_U1_X), .Z0_f (new_AGEMA_signal_1658), .Z1_t (new_AGEMA_signal_1659), .Z1_f (new_AGEMA_signal_1660) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_4_U1_X), .B0_f (new_AGEMA_signal_1658), .B1_t (new_AGEMA_signal_1659), .B1_f (new_AGEMA_signal_1660), .Z0_t (KeyMUX_MUXInst_4_U1_Y), .Z0_f (new_AGEMA_signal_2463), .Z1_t (new_AGEMA_signal_2464), .Z1_f (new_AGEMA_signal_2465) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_4_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_4_U1_Y), .A0_f (new_AGEMA_signal_2463), .A1_t (new_AGEMA_signal_2464), .A1_f (new_AGEMA_signal_2465), .B0_t (Key_s0_t[68]), .B0_f (Key_s0_f[68]), .B1_t (Key_s1_t[68]), .B1_f (Key_s1_f[68]), .Z0_t (SelectedKey[4]), .Z0_f (new_AGEMA_signal_2850), .Z1_t (new_AGEMA_signal_2851), .Z1_f (new_AGEMA_signal_2852) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_5_U1_XOR1_U1 ( .A0_t (Key_s0_t[69]), .A0_f (Key_s0_f[69]), .A1_t (Key_s1_t[69]), .A1_f (Key_s1_f[69]), .B0_t (Key_s0_t[5]), .B0_f (Key_s0_f[5]), .B1_t (Key_s1_t[5]), .B1_f (Key_s1_f[5]), .Z0_t (KeyMUX_MUXInst_5_U1_X), .Z0_f (new_AGEMA_signal_1667), .Z1_t (new_AGEMA_signal_1668), .Z1_f (new_AGEMA_signal_1669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_5_U1_X), .B0_f (new_AGEMA_signal_1667), .B1_t (new_AGEMA_signal_1668), .B1_f (new_AGEMA_signal_1669), .Z0_t (KeyMUX_MUXInst_5_U1_Y), .Z0_f (new_AGEMA_signal_2466), .Z1_t (new_AGEMA_signal_2467), .Z1_f (new_AGEMA_signal_2468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_5_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_5_U1_Y), .A0_f (new_AGEMA_signal_2466), .A1_t (new_AGEMA_signal_2467), .A1_f (new_AGEMA_signal_2468), .B0_t (Key_s0_t[69]), .B0_f (Key_s0_f[69]), .B1_t (Key_s1_t[69]), .B1_f (Key_s1_f[69]), .Z0_t (SelectedKey[5]), .Z0_f (new_AGEMA_signal_2853), .Z1_t (new_AGEMA_signal_2854), .Z1_f (new_AGEMA_signal_2855) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_6_U1_XOR1_U1 ( .A0_t (Key_s0_t[70]), .A0_f (Key_s0_f[70]), .A1_t (Key_s1_t[70]), .A1_f (Key_s1_f[70]), .B0_t (Key_s0_t[6]), .B0_f (Key_s0_f[6]), .B1_t (Key_s1_t[6]), .B1_f (Key_s1_f[6]), .Z0_t (KeyMUX_MUXInst_6_U1_X), .Z0_f (new_AGEMA_signal_1676), .Z1_t (new_AGEMA_signal_1677), .Z1_f (new_AGEMA_signal_1678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_6_U1_X), .B0_f (new_AGEMA_signal_1676), .B1_t (new_AGEMA_signal_1677), .B1_f (new_AGEMA_signal_1678), .Z0_t (KeyMUX_MUXInst_6_U1_Y), .Z0_f (new_AGEMA_signal_2469), .Z1_t (new_AGEMA_signal_2470), .Z1_f (new_AGEMA_signal_2471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_6_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_6_U1_Y), .A0_f (new_AGEMA_signal_2469), .A1_t (new_AGEMA_signal_2470), .A1_f (new_AGEMA_signal_2471), .B0_t (Key_s0_t[70]), .B0_f (Key_s0_f[70]), .B1_t (Key_s1_t[70]), .B1_f (Key_s1_f[70]), .Z0_t (SelectedKey[6]), .Z0_f (new_AGEMA_signal_2856), .Z1_t (new_AGEMA_signal_2857), .Z1_f (new_AGEMA_signal_2858) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_7_U1_XOR1_U1 ( .A0_t (Key_s0_t[71]), .A0_f (Key_s0_f[71]), .A1_t (Key_s1_t[71]), .A1_f (Key_s1_f[71]), .B0_t (Key_s0_t[7]), .B0_f (Key_s0_f[7]), .B1_t (Key_s1_t[7]), .B1_f (Key_s1_f[7]), .Z0_t (KeyMUX_MUXInst_7_U1_X), .Z0_f (new_AGEMA_signal_1685), .Z1_t (new_AGEMA_signal_1686), .Z1_f (new_AGEMA_signal_1687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_7_U1_X), .B0_f (new_AGEMA_signal_1685), .B1_t (new_AGEMA_signal_1686), .B1_f (new_AGEMA_signal_1687), .Z0_t (KeyMUX_MUXInst_7_U1_Y), .Z0_f (new_AGEMA_signal_2472), .Z1_t (new_AGEMA_signal_2473), .Z1_f (new_AGEMA_signal_2474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_7_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_7_U1_Y), .A0_f (new_AGEMA_signal_2472), .A1_t (new_AGEMA_signal_2473), .A1_f (new_AGEMA_signal_2474), .B0_t (Key_s0_t[71]), .B0_f (Key_s0_f[71]), .B1_t (Key_s1_t[71]), .B1_f (Key_s1_f[71]), .Z0_t (SelectedKey[7]), .Z0_f (new_AGEMA_signal_2859), .Z1_t (new_AGEMA_signal_2860), .Z1_f (new_AGEMA_signal_2861) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_8_U1_XOR1_U1 ( .A0_t (Key_s0_t[72]), .A0_f (Key_s0_f[72]), .A1_t (Key_s1_t[72]), .A1_f (Key_s1_f[72]), .B0_t (Key_s0_t[8]), .B0_f (Key_s0_f[8]), .B1_t (Key_s1_t[8]), .B1_f (Key_s1_f[8]), .Z0_t (KeyMUX_MUXInst_8_U1_X), .Z0_f (new_AGEMA_signal_1694), .Z1_t (new_AGEMA_signal_1695), .Z1_f (new_AGEMA_signal_1696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_8_U1_X), .B0_f (new_AGEMA_signal_1694), .B1_t (new_AGEMA_signal_1695), .B1_f (new_AGEMA_signal_1696), .Z0_t (KeyMUX_MUXInst_8_U1_Y), .Z0_f (new_AGEMA_signal_2475), .Z1_t (new_AGEMA_signal_2476), .Z1_f (new_AGEMA_signal_2477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_8_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_8_U1_Y), .A0_f (new_AGEMA_signal_2475), .A1_t (new_AGEMA_signal_2476), .A1_f (new_AGEMA_signal_2477), .B0_t (Key_s0_t[72]), .B0_f (Key_s0_f[72]), .B1_t (Key_s1_t[72]), .B1_f (Key_s1_f[72]), .Z0_t (SelectedKey[8]), .Z0_f (new_AGEMA_signal_2862), .Z1_t (new_AGEMA_signal_2863), .Z1_f (new_AGEMA_signal_2864) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_9_U1_XOR1_U1 ( .A0_t (Key_s0_t[73]), .A0_f (Key_s0_f[73]), .A1_t (Key_s1_t[73]), .A1_f (Key_s1_f[73]), .B0_t (Key_s0_t[9]), .B0_f (Key_s0_f[9]), .B1_t (Key_s1_t[9]), .B1_f (Key_s1_f[9]), .Z0_t (KeyMUX_MUXInst_9_U1_X), .Z0_f (new_AGEMA_signal_1703), .Z1_t (new_AGEMA_signal_1704), .Z1_f (new_AGEMA_signal_1705) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_9_U1_X), .B0_f (new_AGEMA_signal_1703), .B1_t (new_AGEMA_signal_1704), .B1_f (new_AGEMA_signal_1705), .Z0_t (KeyMUX_MUXInst_9_U1_Y), .Z0_f (new_AGEMA_signal_2478), .Z1_t (new_AGEMA_signal_2479), .Z1_f (new_AGEMA_signal_2480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_9_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_9_U1_Y), .A0_f (new_AGEMA_signal_2478), .A1_t (new_AGEMA_signal_2479), .A1_f (new_AGEMA_signal_2480), .B0_t (Key_s0_t[73]), .B0_f (Key_s0_f[73]), .B1_t (Key_s1_t[73]), .B1_f (Key_s1_f[73]), .Z0_t (SelectedKey[9]), .Z0_f (new_AGEMA_signal_2865), .Z1_t (new_AGEMA_signal_2866), .Z1_f (new_AGEMA_signal_2867) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_10_U1_XOR1_U1 ( .A0_t (Key_s0_t[74]), .A0_f (Key_s0_f[74]), .A1_t (Key_s1_t[74]), .A1_f (Key_s1_f[74]), .B0_t (Key_s0_t[10]), .B0_f (Key_s0_f[10]), .B1_t (Key_s1_t[10]), .B1_f (Key_s1_f[10]), .Z0_t (KeyMUX_MUXInst_10_U1_X), .Z0_f (new_AGEMA_signal_1712), .Z1_t (new_AGEMA_signal_1713), .Z1_f (new_AGEMA_signal_1714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_10_U1_X), .B0_f (new_AGEMA_signal_1712), .B1_t (new_AGEMA_signal_1713), .B1_f (new_AGEMA_signal_1714), .Z0_t (KeyMUX_MUXInst_10_U1_Y), .Z0_f (new_AGEMA_signal_2481), .Z1_t (new_AGEMA_signal_2482), .Z1_f (new_AGEMA_signal_2483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_10_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_10_U1_Y), .A0_f (new_AGEMA_signal_2481), .A1_t (new_AGEMA_signal_2482), .A1_f (new_AGEMA_signal_2483), .B0_t (Key_s0_t[74]), .B0_f (Key_s0_f[74]), .B1_t (Key_s1_t[74]), .B1_f (Key_s1_f[74]), .Z0_t (SelectedKey[10]), .Z0_f (new_AGEMA_signal_2868), .Z1_t (new_AGEMA_signal_2869), .Z1_f (new_AGEMA_signal_2870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_11_U1_XOR1_U1 ( .A0_t (Key_s0_t[75]), .A0_f (Key_s0_f[75]), .A1_t (Key_s1_t[75]), .A1_f (Key_s1_f[75]), .B0_t (Key_s0_t[11]), .B0_f (Key_s0_f[11]), .B1_t (Key_s1_t[11]), .B1_f (Key_s1_f[11]), .Z0_t (KeyMUX_MUXInst_11_U1_X), .Z0_f (new_AGEMA_signal_1721), .Z1_t (new_AGEMA_signal_1722), .Z1_f (new_AGEMA_signal_1723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_11_U1_X), .B0_f (new_AGEMA_signal_1721), .B1_t (new_AGEMA_signal_1722), .B1_f (new_AGEMA_signal_1723), .Z0_t (KeyMUX_MUXInst_11_U1_Y), .Z0_f (new_AGEMA_signal_2484), .Z1_t (new_AGEMA_signal_2485), .Z1_f (new_AGEMA_signal_2486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_11_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_11_U1_Y), .A0_f (new_AGEMA_signal_2484), .A1_t (new_AGEMA_signal_2485), .A1_f (new_AGEMA_signal_2486), .B0_t (Key_s0_t[75]), .B0_f (Key_s0_f[75]), .B1_t (Key_s1_t[75]), .B1_f (Key_s1_f[75]), .Z0_t (SelectedKey[11]), .Z0_f (new_AGEMA_signal_2871), .Z1_t (new_AGEMA_signal_2872), .Z1_f (new_AGEMA_signal_2873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_12_U1_XOR1_U1 ( .A0_t (Key_s0_t[76]), .A0_f (Key_s0_f[76]), .A1_t (Key_s1_t[76]), .A1_f (Key_s1_f[76]), .B0_t (Key_s0_t[12]), .B0_f (Key_s0_f[12]), .B1_t (Key_s1_t[12]), .B1_f (Key_s1_f[12]), .Z0_t (KeyMUX_MUXInst_12_U1_X), .Z0_f (new_AGEMA_signal_1730), .Z1_t (new_AGEMA_signal_1731), .Z1_f (new_AGEMA_signal_1732) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_12_U1_X), .B0_f (new_AGEMA_signal_1730), .B1_t (new_AGEMA_signal_1731), .B1_f (new_AGEMA_signal_1732), .Z0_t (KeyMUX_MUXInst_12_U1_Y), .Z0_f (new_AGEMA_signal_2487), .Z1_t (new_AGEMA_signal_2488), .Z1_f (new_AGEMA_signal_2489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_12_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_12_U1_Y), .A0_f (new_AGEMA_signal_2487), .A1_t (new_AGEMA_signal_2488), .A1_f (new_AGEMA_signal_2489), .B0_t (Key_s0_t[76]), .B0_f (Key_s0_f[76]), .B1_t (Key_s1_t[76]), .B1_f (Key_s1_f[76]), .Z0_t (SelectedKey[12]), .Z0_f (new_AGEMA_signal_2874), .Z1_t (new_AGEMA_signal_2875), .Z1_f (new_AGEMA_signal_2876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_13_U1_XOR1_U1 ( .A0_t (Key_s0_t[77]), .A0_f (Key_s0_f[77]), .A1_t (Key_s1_t[77]), .A1_f (Key_s1_f[77]), .B0_t (Key_s0_t[13]), .B0_f (Key_s0_f[13]), .B1_t (Key_s1_t[13]), .B1_f (Key_s1_f[13]), .Z0_t (KeyMUX_MUXInst_13_U1_X), .Z0_f (new_AGEMA_signal_1739), .Z1_t (new_AGEMA_signal_1740), .Z1_f (new_AGEMA_signal_1741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_13_U1_X), .B0_f (new_AGEMA_signal_1739), .B1_t (new_AGEMA_signal_1740), .B1_f (new_AGEMA_signal_1741), .Z0_t (KeyMUX_MUXInst_13_U1_Y), .Z0_f (new_AGEMA_signal_2490), .Z1_t (new_AGEMA_signal_2491), .Z1_f (new_AGEMA_signal_2492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_13_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_13_U1_Y), .A0_f (new_AGEMA_signal_2490), .A1_t (new_AGEMA_signal_2491), .A1_f (new_AGEMA_signal_2492), .B0_t (Key_s0_t[77]), .B0_f (Key_s0_f[77]), .B1_t (Key_s1_t[77]), .B1_f (Key_s1_f[77]), .Z0_t (SelectedKey[13]), .Z0_f (new_AGEMA_signal_2877), .Z1_t (new_AGEMA_signal_2878), .Z1_f (new_AGEMA_signal_2879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_14_U1_XOR1_U1 ( .A0_t (Key_s0_t[78]), .A0_f (Key_s0_f[78]), .A1_t (Key_s1_t[78]), .A1_f (Key_s1_f[78]), .B0_t (Key_s0_t[14]), .B0_f (Key_s0_f[14]), .B1_t (Key_s1_t[14]), .B1_f (Key_s1_f[14]), .Z0_t (KeyMUX_MUXInst_14_U1_X), .Z0_f (new_AGEMA_signal_1748), .Z1_t (new_AGEMA_signal_1749), .Z1_f (new_AGEMA_signal_1750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_14_U1_X), .B0_f (new_AGEMA_signal_1748), .B1_t (new_AGEMA_signal_1749), .B1_f (new_AGEMA_signal_1750), .Z0_t (KeyMUX_MUXInst_14_U1_Y), .Z0_f (new_AGEMA_signal_2493), .Z1_t (new_AGEMA_signal_2494), .Z1_f (new_AGEMA_signal_2495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_14_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_14_U1_Y), .A0_f (new_AGEMA_signal_2493), .A1_t (new_AGEMA_signal_2494), .A1_f (new_AGEMA_signal_2495), .B0_t (Key_s0_t[78]), .B0_f (Key_s0_f[78]), .B1_t (Key_s1_t[78]), .B1_f (Key_s1_f[78]), .Z0_t (SelectedKey[14]), .Z0_f (new_AGEMA_signal_2880), .Z1_t (new_AGEMA_signal_2881), .Z1_f (new_AGEMA_signal_2882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_15_U1_XOR1_U1 ( .A0_t (Key_s0_t[79]), .A0_f (Key_s0_f[79]), .A1_t (Key_s1_t[79]), .A1_f (Key_s1_f[79]), .B0_t (Key_s0_t[15]), .B0_f (Key_s0_f[15]), .B1_t (Key_s1_t[15]), .B1_f (Key_s1_f[15]), .Z0_t (KeyMUX_MUXInst_15_U1_X), .Z0_f (new_AGEMA_signal_1757), .Z1_t (new_AGEMA_signal_1758), .Z1_f (new_AGEMA_signal_1759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_15_U1_X), .B0_f (new_AGEMA_signal_1757), .B1_t (new_AGEMA_signal_1758), .B1_f (new_AGEMA_signal_1759), .Z0_t (KeyMUX_MUXInst_15_U1_Y), .Z0_f (new_AGEMA_signal_2496), .Z1_t (new_AGEMA_signal_2497), .Z1_f (new_AGEMA_signal_2498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_15_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_15_U1_Y), .A0_f (new_AGEMA_signal_2496), .A1_t (new_AGEMA_signal_2497), .A1_f (new_AGEMA_signal_2498), .B0_t (Key_s0_t[79]), .B0_f (Key_s0_f[79]), .B1_t (Key_s1_t[79]), .B1_f (Key_s1_f[79]), .Z0_t (SelectedKey[15]), .Z0_f (new_AGEMA_signal_2883), .Z1_t (new_AGEMA_signal_2884), .Z1_f (new_AGEMA_signal_2885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_16_U1_XOR1_U1 ( .A0_t (Key_s0_t[80]), .A0_f (Key_s0_f[80]), .A1_t (Key_s1_t[80]), .A1_f (Key_s1_f[80]), .B0_t (Key_s0_t[16]), .B0_f (Key_s0_f[16]), .B1_t (Key_s1_t[16]), .B1_f (Key_s1_f[16]), .Z0_t (KeyMUX_MUXInst_16_U1_X), .Z0_f (new_AGEMA_signal_1766), .Z1_t (new_AGEMA_signal_1767), .Z1_f (new_AGEMA_signal_1768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_16_U1_X), .B0_f (new_AGEMA_signal_1766), .B1_t (new_AGEMA_signal_1767), .B1_f (new_AGEMA_signal_1768), .Z0_t (KeyMUX_MUXInst_16_U1_Y), .Z0_f (new_AGEMA_signal_2499), .Z1_t (new_AGEMA_signal_2500), .Z1_f (new_AGEMA_signal_2501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_16_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_16_U1_Y), .A0_f (new_AGEMA_signal_2499), .A1_t (new_AGEMA_signal_2500), .A1_f (new_AGEMA_signal_2501), .B0_t (Key_s0_t[80]), .B0_f (Key_s0_f[80]), .B1_t (Key_s1_t[80]), .B1_f (Key_s1_f[80]), .Z0_t (SelectedKey[16]), .Z0_f (new_AGEMA_signal_2886), .Z1_t (new_AGEMA_signal_2887), .Z1_f (new_AGEMA_signal_2888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_17_U1_XOR1_U1 ( .A0_t (Key_s0_t[81]), .A0_f (Key_s0_f[81]), .A1_t (Key_s1_t[81]), .A1_f (Key_s1_f[81]), .B0_t (Key_s0_t[17]), .B0_f (Key_s0_f[17]), .B1_t (Key_s1_t[17]), .B1_f (Key_s1_f[17]), .Z0_t (KeyMUX_MUXInst_17_U1_X), .Z0_f (new_AGEMA_signal_1775), .Z1_t (new_AGEMA_signal_1776), .Z1_f (new_AGEMA_signal_1777) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_17_U1_X), .B0_f (new_AGEMA_signal_1775), .B1_t (new_AGEMA_signal_1776), .B1_f (new_AGEMA_signal_1777), .Z0_t (KeyMUX_MUXInst_17_U1_Y), .Z0_f (new_AGEMA_signal_2502), .Z1_t (new_AGEMA_signal_2503), .Z1_f (new_AGEMA_signal_2504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_17_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_17_U1_Y), .A0_f (new_AGEMA_signal_2502), .A1_t (new_AGEMA_signal_2503), .A1_f (new_AGEMA_signal_2504), .B0_t (Key_s0_t[81]), .B0_f (Key_s0_f[81]), .B1_t (Key_s1_t[81]), .B1_f (Key_s1_f[81]), .Z0_t (SelectedKey[17]), .Z0_f (new_AGEMA_signal_2889), .Z1_t (new_AGEMA_signal_2890), .Z1_f (new_AGEMA_signal_2891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_18_U1_XOR1_U1 ( .A0_t (Key_s0_t[82]), .A0_f (Key_s0_f[82]), .A1_t (Key_s1_t[82]), .A1_f (Key_s1_f[82]), .B0_t (Key_s0_t[18]), .B0_f (Key_s0_f[18]), .B1_t (Key_s1_t[18]), .B1_f (Key_s1_f[18]), .Z0_t (KeyMUX_MUXInst_18_U1_X), .Z0_f (new_AGEMA_signal_1784), .Z1_t (new_AGEMA_signal_1785), .Z1_f (new_AGEMA_signal_1786) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_18_U1_X), .B0_f (new_AGEMA_signal_1784), .B1_t (new_AGEMA_signal_1785), .B1_f (new_AGEMA_signal_1786), .Z0_t (KeyMUX_MUXInst_18_U1_Y), .Z0_f (new_AGEMA_signal_2505), .Z1_t (new_AGEMA_signal_2506), .Z1_f (new_AGEMA_signal_2507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_18_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_18_U1_Y), .A0_f (new_AGEMA_signal_2505), .A1_t (new_AGEMA_signal_2506), .A1_f (new_AGEMA_signal_2507), .B0_t (Key_s0_t[82]), .B0_f (Key_s0_f[82]), .B1_t (Key_s1_t[82]), .B1_f (Key_s1_f[82]), .Z0_t (SelectedKey[18]), .Z0_f (new_AGEMA_signal_2892), .Z1_t (new_AGEMA_signal_2893), .Z1_f (new_AGEMA_signal_2894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_19_U1_XOR1_U1 ( .A0_t (Key_s0_t[83]), .A0_f (Key_s0_f[83]), .A1_t (Key_s1_t[83]), .A1_f (Key_s1_f[83]), .B0_t (Key_s0_t[19]), .B0_f (Key_s0_f[19]), .B1_t (Key_s1_t[19]), .B1_f (Key_s1_f[19]), .Z0_t (KeyMUX_MUXInst_19_U1_X), .Z0_f (new_AGEMA_signal_1793), .Z1_t (new_AGEMA_signal_1794), .Z1_f (new_AGEMA_signal_1795) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_19_U1_X), .B0_f (new_AGEMA_signal_1793), .B1_t (new_AGEMA_signal_1794), .B1_f (new_AGEMA_signal_1795), .Z0_t (KeyMUX_MUXInst_19_U1_Y), .Z0_f (new_AGEMA_signal_2508), .Z1_t (new_AGEMA_signal_2509), .Z1_f (new_AGEMA_signal_2510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_19_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_19_U1_Y), .A0_f (new_AGEMA_signal_2508), .A1_t (new_AGEMA_signal_2509), .A1_f (new_AGEMA_signal_2510), .B0_t (Key_s0_t[83]), .B0_f (Key_s0_f[83]), .B1_t (Key_s1_t[83]), .B1_f (Key_s1_f[83]), .Z0_t (SelectedKey[19]), .Z0_f (new_AGEMA_signal_2895), .Z1_t (new_AGEMA_signal_2896), .Z1_f (new_AGEMA_signal_2897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_20_U1_XOR1_U1 ( .A0_t (Key_s0_t[84]), .A0_f (Key_s0_f[84]), .A1_t (Key_s1_t[84]), .A1_f (Key_s1_f[84]), .B0_t (Key_s0_t[20]), .B0_f (Key_s0_f[20]), .B1_t (Key_s1_t[20]), .B1_f (Key_s1_f[20]), .Z0_t (KeyMUX_MUXInst_20_U1_X), .Z0_f (new_AGEMA_signal_1802), .Z1_t (new_AGEMA_signal_1803), .Z1_f (new_AGEMA_signal_1804) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_20_U1_X), .B0_f (new_AGEMA_signal_1802), .B1_t (new_AGEMA_signal_1803), .B1_f (new_AGEMA_signal_1804), .Z0_t (KeyMUX_MUXInst_20_U1_Y), .Z0_f (new_AGEMA_signal_2511), .Z1_t (new_AGEMA_signal_2512), .Z1_f (new_AGEMA_signal_2513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_20_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_20_U1_Y), .A0_f (new_AGEMA_signal_2511), .A1_t (new_AGEMA_signal_2512), .A1_f (new_AGEMA_signal_2513), .B0_t (Key_s0_t[84]), .B0_f (Key_s0_f[84]), .B1_t (Key_s1_t[84]), .B1_f (Key_s1_f[84]), .Z0_t (SelectedKey[20]), .Z0_f (new_AGEMA_signal_2898), .Z1_t (new_AGEMA_signal_2899), .Z1_f (new_AGEMA_signal_2900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_21_U1_XOR1_U1 ( .A0_t (Key_s0_t[85]), .A0_f (Key_s0_f[85]), .A1_t (Key_s1_t[85]), .A1_f (Key_s1_f[85]), .B0_t (Key_s0_t[21]), .B0_f (Key_s0_f[21]), .B1_t (Key_s1_t[21]), .B1_f (Key_s1_f[21]), .Z0_t (KeyMUX_MUXInst_21_U1_X), .Z0_f (new_AGEMA_signal_1811), .Z1_t (new_AGEMA_signal_1812), .Z1_f (new_AGEMA_signal_1813) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_21_U1_X), .B0_f (new_AGEMA_signal_1811), .B1_t (new_AGEMA_signal_1812), .B1_f (new_AGEMA_signal_1813), .Z0_t (KeyMUX_MUXInst_21_U1_Y), .Z0_f (new_AGEMA_signal_2514), .Z1_t (new_AGEMA_signal_2515), .Z1_f (new_AGEMA_signal_2516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_21_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_21_U1_Y), .A0_f (new_AGEMA_signal_2514), .A1_t (new_AGEMA_signal_2515), .A1_f (new_AGEMA_signal_2516), .B0_t (Key_s0_t[85]), .B0_f (Key_s0_f[85]), .B1_t (Key_s1_t[85]), .B1_f (Key_s1_f[85]), .Z0_t (SelectedKey[21]), .Z0_f (new_AGEMA_signal_2901), .Z1_t (new_AGEMA_signal_2902), .Z1_f (new_AGEMA_signal_2903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_22_U1_XOR1_U1 ( .A0_t (Key_s0_t[86]), .A0_f (Key_s0_f[86]), .A1_t (Key_s1_t[86]), .A1_f (Key_s1_f[86]), .B0_t (Key_s0_t[22]), .B0_f (Key_s0_f[22]), .B1_t (Key_s1_t[22]), .B1_f (Key_s1_f[22]), .Z0_t (KeyMUX_MUXInst_22_U1_X), .Z0_f (new_AGEMA_signal_1820), .Z1_t (new_AGEMA_signal_1821), .Z1_f (new_AGEMA_signal_1822) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_22_U1_X), .B0_f (new_AGEMA_signal_1820), .B1_t (new_AGEMA_signal_1821), .B1_f (new_AGEMA_signal_1822), .Z0_t (KeyMUX_MUXInst_22_U1_Y), .Z0_f (new_AGEMA_signal_2517), .Z1_t (new_AGEMA_signal_2518), .Z1_f (new_AGEMA_signal_2519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_22_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_22_U1_Y), .A0_f (new_AGEMA_signal_2517), .A1_t (new_AGEMA_signal_2518), .A1_f (new_AGEMA_signal_2519), .B0_t (Key_s0_t[86]), .B0_f (Key_s0_f[86]), .B1_t (Key_s1_t[86]), .B1_f (Key_s1_f[86]), .Z0_t (SelectedKey[22]), .Z0_f (new_AGEMA_signal_2904), .Z1_t (new_AGEMA_signal_2905), .Z1_f (new_AGEMA_signal_2906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_23_U1_XOR1_U1 ( .A0_t (Key_s0_t[87]), .A0_f (Key_s0_f[87]), .A1_t (Key_s1_t[87]), .A1_f (Key_s1_f[87]), .B0_t (Key_s0_t[23]), .B0_f (Key_s0_f[23]), .B1_t (Key_s1_t[23]), .B1_f (Key_s1_f[23]), .Z0_t (KeyMUX_MUXInst_23_U1_X), .Z0_f (new_AGEMA_signal_1829), .Z1_t (new_AGEMA_signal_1830), .Z1_f (new_AGEMA_signal_1831) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_23_U1_X), .B0_f (new_AGEMA_signal_1829), .B1_t (new_AGEMA_signal_1830), .B1_f (new_AGEMA_signal_1831), .Z0_t (KeyMUX_MUXInst_23_U1_Y), .Z0_f (new_AGEMA_signal_2520), .Z1_t (new_AGEMA_signal_2521), .Z1_f (new_AGEMA_signal_2522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_23_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_23_U1_Y), .A0_f (new_AGEMA_signal_2520), .A1_t (new_AGEMA_signal_2521), .A1_f (new_AGEMA_signal_2522), .B0_t (Key_s0_t[87]), .B0_f (Key_s0_f[87]), .B1_t (Key_s1_t[87]), .B1_f (Key_s1_f[87]), .Z0_t (SelectedKey[23]), .Z0_f (new_AGEMA_signal_2907), .Z1_t (new_AGEMA_signal_2908), .Z1_f (new_AGEMA_signal_2909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_24_U1_XOR1_U1 ( .A0_t (Key_s0_t[88]), .A0_f (Key_s0_f[88]), .A1_t (Key_s1_t[88]), .A1_f (Key_s1_f[88]), .B0_t (Key_s0_t[24]), .B0_f (Key_s0_f[24]), .B1_t (Key_s1_t[24]), .B1_f (Key_s1_f[24]), .Z0_t (KeyMUX_MUXInst_24_U1_X), .Z0_f (new_AGEMA_signal_1838), .Z1_t (new_AGEMA_signal_1839), .Z1_f (new_AGEMA_signal_1840) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_24_U1_X), .B0_f (new_AGEMA_signal_1838), .B1_t (new_AGEMA_signal_1839), .B1_f (new_AGEMA_signal_1840), .Z0_t (KeyMUX_MUXInst_24_U1_Y), .Z0_f (new_AGEMA_signal_2523), .Z1_t (new_AGEMA_signal_2524), .Z1_f (new_AGEMA_signal_2525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_24_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_24_U1_Y), .A0_f (new_AGEMA_signal_2523), .A1_t (new_AGEMA_signal_2524), .A1_f (new_AGEMA_signal_2525), .B0_t (Key_s0_t[88]), .B0_f (Key_s0_f[88]), .B1_t (Key_s1_t[88]), .B1_f (Key_s1_f[88]), .Z0_t (SelectedKey[24]), .Z0_f (new_AGEMA_signal_2910), .Z1_t (new_AGEMA_signal_2911), .Z1_f (new_AGEMA_signal_2912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_25_U1_XOR1_U1 ( .A0_t (Key_s0_t[89]), .A0_f (Key_s0_f[89]), .A1_t (Key_s1_t[89]), .A1_f (Key_s1_f[89]), .B0_t (Key_s0_t[25]), .B0_f (Key_s0_f[25]), .B1_t (Key_s1_t[25]), .B1_f (Key_s1_f[25]), .Z0_t (KeyMUX_MUXInst_25_U1_X), .Z0_f (new_AGEMA_signal_1847), .Z1_t (new_AGEMA_signal_1848), .Z1_f (new_AGEMA_signal_1849) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_25_U1_X), .B0_f (new_AGEMA_signal_1847), .B1_t (new_AGEMA_signal_1848), .B1_f (new_AGEMA_signal_1849), .Z0_t (KeyMUX_MUXInst_25_U1_Y), .Z0_f (new_AGEMA_signal_2526), .Z1_t (new_AGEMA_signal_2527), .Z1_f (new_AGEMA_signal_2528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_25_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_25_U1_Y), .A0_f (new_AGEMA_signal_2526), .A1_t (new_AGEMA_signal_2527), .A1_f (new_AGEMA_signal_2528), .B0_t (Key_s0_t[89]), .B0_f (Key_s0_f[89]), .B1_t (Key_s1_t[89]), .B1_f (Key_s1_f[89]), .Z0_t (SelectedKey[25]), .Z0_f (new_AGEMA_signal_2913), .Z1_t (new_AGEMA_signal_2914), .Z1_f (new_AGEMA_signal_2915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_26_U1_XOR1_U1 ( .A0_t (Key_s0_t[90]), .A0_f (Key_s0_f[90]), .A1_t (Key_s1_t[90]), .A1_f (Key_s1_f[90]), .B0_t (Key_s0_t[26]), .B0_f (Key_s0_f[26]), .B1_t (Key_s1_t[26]), .B1_f (Key_s1_f[26]), .Z0_t (KeyMUX_MUXInst_26_U1_X), .Z0_f (new_AGEMA_signal_1856), .Z1_t (new_AGEMA_signal_1857), .Z1_f (new_AGEMA_signal_1858) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_26_U1_X), .B0_f (new_AGEMA_signal_1856), .B1_t (new_AGEMA_signal_1857), .B1_f (new_AGEMA_signal_1858), .Z0_t (KeyMUX_MUXInst_26_U1_Y), .Z0_f (new_AGEMA_signal_2529), .Z1_t (new_AGEMA_signal_2530), .Z1_f (new_AGEMA_signal_2531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_26_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_26_U1_Y), .A0_f (new_AGEMA_signal_2529), .A1_t (new_AGEMA_signal_2530), .A1_f (new_AGEMA_signal_2531), .B0_t (Key_s0_t[90]), .B0_f (Key_s0_f[90]), .B1_t (Key_s1_t[90]), .B1_f (Key_s1_f[90]), .Z0_t (SelectedKey[26]), .Z0_f (new_AGEMA_signal_2916), .Z1_t (new_AGEMA_signal_2917), .Z1_f (new_AGEMA_signal_2918) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_27_U1_XOR1_U1 ( .A0_t (Key_s0_t[91]), .A0_f (Key_s0_f[91]), .A1_t (Key_s1_t[91]), .A1_f (Key_s1_f[91]), .B0_t (Key_s0_t[27]), .B0_f (Key_s0_f[27]), .B1_t (Key_s1_t[27]), .B1_f (Key_s1_f[27]), .Z0_t (KeyMUX_MUXInst_27_U1_X), .Z0_f (new_AGEMA_signal_1865), .Z1_t (new_AGEMA_signal_1866), .Z1_f (new_AGEMA_signal_1867) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_27_U1_X), .B0_f (new_AGEMA_signal_1865), .B1_t (new_AGEMA_signal_1866), .B1_f (new_AGEMA_signal_1867), .Z0_t (KeyMUX_MUXInst_27_U1_Y), .Z0_f (new_AGEMA_signal_2532), .Z1_t (new_AGEMA_signal_2533), .Z1_f (new_AGEMA_signal_2534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_27_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_27_U1_Y), .A0_f (new_AGEMA_signal_2532), .A1_t (new_AGEMA_signal_2533), .A1_f (new_AGEMA_signal_2534), .B0_t (Key_s0_t[91]), .B0_f (Key_s0_f[91]), .B1_t (Key_s1_t[91]), .B1_f (Key_s1_f[91]), .Z0_t (SelectedKey[27]), .Z0_f (new_AGEMA_signal_2919), .Z1_t (new_AGEMA_signal_2920), .Z1_f (new_AGEMA_signal_2921) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_28_U1_XOR1_U1 ( .A0_t (Key_s0_t[92]), .A0_f (Key_s0_f[92]), .A1_t (Key_s1_t[92]), .A1_f (Key_s1_f[92]), .B0_t (Key_s0_t[28]), .B0_f (Key_s0_f[28]), .B1_t (Key_s1_t[28]), .B1_f (Key_s1_f[28]), .Z0_t (KeyMUX_MUXInst_28_U1_X), .Z0_f (new_AGEMA_signal_1874), .Z1_t (new_AGEMA_signal_1875), .Z1_f (new_AGEMA_signal_1876) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_28_U1_X), .B0_f (new_AGEMA_signal_1874), .B1_t (new_AGEMA_signal_1875), .B1_f (new_AGEMA_signal_1876), .Z0_t (KeyMUX_MUXInst_28_U1_Y), .Z0_f (new_AGEMA_signal_2535), .Z1_t (new_AGEMA_signal_2536), .Z1_f (new_AGEMA_signal_2537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_28_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_28_U1_Y), .A0_f (new_AGEMA_signal_2535), .A1_t (new_AGEMA_signal_2536), .A1_f (new_AGEMA_signal_2537), .B0_t (Key_s0_t[92]), .B0_f (Key_s0_f[92]), .B1_t (Key_s1_t[92]), .B1_f (Key_s1_f[92]), .Z0_t (SelectedKey[28]), .Z0_f (new_AGEMA_signal_2922), .Z1_t (new_AGEMA_signal_2923), .Z1_f (new_AGEMA_signal_2924) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_29_U1_XOR1_U1 ( .A0_t (Key_s0_t[93]), .A0_f (Key_s0_f[93]), .A1_t (Key_s1_t[93]), .A1_f (Key_s1_f[93]), .B0_t (Key_s0_t[29]), .B0_f (Key_s0_f[29]), .B1_t (Key_s1_t[29]), .B1_f (Key_s1_f[29]), .Z0_t (KeyMUX_MUXInst_29_U1_X), .Z0_f (new_AGEMA_signal_1883), .Z1_t (new_AGEMA_signal_1884), .Z1_f (new_AGEMA_signal_1885) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_29_U1_X), .B0_f (new_AGEMA_signal_1883), .B1_t (new_AGEMA_signal_1884), .B1_f (new_AGEMA_signal_1885), .Z0_t (KeyMUX_MUXInst_29_U1_Y), .Z0_f (new_AGEMA_signal_2538), .Z1_t (new_AGEMA_signal_2539), .Z1_f (new_AGEMA_signal_2540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_29_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_29_U1_Y), .A0_f (new_AGEMA_signal_2538), .A1_t (new_AGEMA_signal_2539), .A1_f (new_AGEMA_signal_2540), .B0_t (Key_s0_t[93]), .B0_f (Key_s0_f[93]), .B1_t (Key_s1_t[93]), .B1_f (Key_s1_f[93]), .Z0_t (SelectedKey[29]), .Z0_f (new_AGEMA_signal_2925), .Z1_t (new_AGEMA_signal_2926), .Z1_f (new_AGEMA_signal_2927) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_30_U1_XOR1_U1 ( .A0_t (Key_s0_t[94]), .A0_f (Key_s0_f[94]), .A1_t (Key_s1_t[94]), .A1_f (Key_s1_f[94]), .B0_t (Key_s0_t[30]), .B0_f (Key_s0_f[30]), .B1_t (Key_s1_t[30]), .B1_f (Key_s1_f[30]), .Z0_t (KeyMUX_MUXInst_30_U1_X), .Z0_f (new_AGEMA_signal_1892), .Z1_t (new_AGEMA_signal_1893), .Z1_f (new_AGEMA_signal_1894) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_30_U1_X), .B0_f (new_AGEMA_signal_1892), .B1_t (new_AGEMA_signal_1893), .B1_f (new_AGEMA_signal_1894), .Z0_t (KeyMUX_MUXInst_30_U1_Y), .Z0_f (new_AGEMA_signal_2541), .Z1_t (new_AGEMA_signal_2542), .Z1_f (new_AGEMA_signal_2543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_30_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_30_U1_Y), .A0_f (new_AGEMA_signal_2541), .A1_t (new_AGEMA_signal_2542), .A1_f (new_AGEMA_signal_2543), .B0_t (Key_s0_t[94]), .B0_f (Key_s0_f[94]), .B1_t (Key_s1_t[94]), .B1_f (Key_s1_f[94]), .Z0_t (SelectedKey[30]), .Z0_f (new_AGEMA_signal_2928), .Z1_t (new_AGEMA_signal_2929), .Z1_f (new_AGEMA_signal_2930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_31_U1_XOR1_U1 ( .A0_t (Key_s0_t[95]), .A0_f (Key_s0_f[95]), .A1_t (Key_s1_t[95]), .A1_f (Key_s1_f[95]), .B0_t (Key_s0_t[31]), .B0_f (Key_s0_f[31]), .B1_t (Key_s1_t[31]), .B1_f (Key_s1_f[31]), .Z0_t (KeyMUX_MUXInst_31_U1_X), .Z0_f (new_AGEMA_signal_1901), .Z1_t (new_AGEMA_signal_1902), .Z1_f (new_AGEMA_signal_1903) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_31_U1_X), .B0_f (new_AGEMA_signal_1901), .B1_t (new_AGEMA_signal_1902), .B1_f (new_AGEMA_signal_1903), .Z0_t (KeyMUX_MUXInst_31_U1_Y), .Z0_f (new_AGEMA_signal_2544), .Z1_t (new_AGEMA_signal_2545), .Z1_f (new_AGEMA_signal_2546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_31_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_31_U1_Y), .A0_f (new_AGEMA_signal_2544), .A1_t (new_AGEMA_signal_2545), .A1_f (new_AGEMA_signal_2546), .B0_t (Key_s0_t[95]), .B0_f (Key_s0_f[95]), .B1_t (Key_s1_t[95]), .B1_f (Key_s1_f[95]), .Z0_t (SelectedKey[31]), .Z0_f (new_AGEMA_signal_2931), .Z1_t (new_AGEMA_signal_2932), .Z1_f (new_AGEMA_signal_2933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_32_U1_XOR1_U1 ( .A0_t (Key_s0_t[96]), .A0_f (Key_s0_f[96]), .A1_t (Key_s1_t[96]), .A1_f (Key_s1_f[96]), .B0_t (Key_s0_t[32]), .B0_f (Key_s0_f[32]), .B1_t (Key_s1_t[32]), .B1_f (Key_s1_f[32]), .Z0_t (KeyMUX_MUXInst_32_U1_X), .Z0_f (new_AGEMA_signal_1910), .Z1_t (new_AGEMA_signal_1911), .Z1_f (new_AGEMA_signal_1912) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_32_U1_X), .B0_f (new_AGEMA_signal_1910), .B1_t (new_AGEMA_signal_1911), .B1_f (new_AGEMA_signal_1912), .Z0_t (KeyMUX_MUXInst_32_U1_Y), .Z0_f (new_AGEMA_signal_2547), .Z1_t (new_AGEMA_signal_2548), .Z1_f (new_AGEMA_signal_2549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_32_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_32_U1_Y), .A0_f (new_AGEMA_signal_2547), .A1_t (new_AGEMA_signal_2548), .A1_f (new_AGEMA_signal_2549), .B0_t (Key_s0_t[96]), .B0_f (Key_s0_f[96]), .B1_t (Key_s1_t[96]), .B1_f (Key_s1_f[96]), .Z0_t (SelectedKey[32]), .Z0_f (new_AGEMA_signal_2934), .Z1_t (new_AGEMA_signal_2935), .Z1_f (new_AGEMA_signal_2936) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_33_U1_XOR1_U1 ( .A0_t (Key_s0_t[97]), .A0_f (Key_s0_f[97]), .A1_t (Key_s1_t[97]), .A1_f (Key_s1_f[97]), .B0_t (Key_s0_t[33]), .B0_f (Key_s0_f[33]), .B1_t (Key_s1_t[33]), .B1_f (Key_s1_f[33]), .Z0_t (KeyMUX_MUXInst_33_U1_X), .Z0_f (new_AGEMA_signal_1919), .Z1_t (new_AGEMA_signal_1920), .Z1_f (new_AGEMA_signal_1921) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_33_U1_X), .B0_f (new_AGEMA_signal_1919), .B1_t (new_AGEMA_signal_1920), .B1_f (new_AGEMA_signal_1921), .Z0_t (KeyMUX_MUXInst_33_U1_Y), .Z0_f (new_AGEMA_signal_2550), .Z1_t (new_AGEMA_signal_2551), .Z1_f (new_AGEMA_signal_2552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_33_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_33_U1_Y), .A0_f (new_AGEMA_signal_2550), .A1_t (new_AGEMA_signal_2551), .A1_f (new_AGEMA_signal_2552), .B0_t (Key_s0_t[97]), .B0_f (Key_s0_f[97]), .B1_t (Key_s1_t[97]), .B1_f (Key_s1_f[97]), .Z0_t (SelectedKey[33]), .Z0_f (new_AGEMA_signal_2937), .Z1_t (new_AGEMA_signal_2938), .Z1_f (new_AGEMA_signal_2939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_34_U1_XOR1_U1 ( .A0_t (Key_s0_t[98]), .A0_f (Key_s0_f[98]), .A1_t (Key_s1_t[98]), .A1_f (Key_s1_f[98]), .B0_t (Key_s0_t[34]), .B0_f (Key_s0_f[34]), .B1_t (Key_s1_t[34]), .B1_f (Key_s1_f[34]), .Z0_t (KeyMUX_MUXInst_34_U1_X), .Z0_f (new_AGEMA_signal_1928), .Z1_t (new_AGEMA_signal_1929), .Z1_f (new_AGEMA_signal_1930) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_34_U1_X), .B0_f (new_AGEMA_signal_1928), .B1_t (new_AGEMA_signal_1929), .B1_f (new_AGEMA_signal_1930), .Z0_t (KeyMUX_MUXInst_34_U1_Y), .Z0_f (new_AGEMA_signal_2553), .Z1_t (new_AGEMA_signal_2554), .Z1_f (new_AGEMA_signal_2555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_34_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_34_U1_Y), .A0_f (new_AGEMA_signal_2553), .A1_t (new_AGEMA_signal_2554), .A1_f (new_AGEMA_signal_2555), .B0_t (Key_s0_t[98]), .B0_f (Key_s0_f[98]), .B1_t (Key_s1_t[98]), .B1_f (Key_s1_f[98]), .Z0_t (SelectedKey[34]), .Z0_f (new_AGEMA_signal_2940), .Z1_t (new_AGEMA_signal_2941), .Z1_f (new_AGEMA_signal_2942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_35_U1_XOR1_U1 ( .A0_t (Key_s0_t[99]), .A0_f (Key_s0_f[99]), .A1_t (Key_s1_t[99]), .A1_f (Key_s1_f[99]), .B0_t (Key_s0_t[35]), .B0_f (Key_s0_f[35]), .B1_t (Key_s1_t[35]), .B1_f (Key_s1_f[35]), .Z0_t (KeyMUX_MUXInst_35_U1_X), .Z0_f (new_AGEMA_signal_1937), .Z1_t (new_AGEMA_signal_1938), .Z1_f (new_AGEMA_signal_1939) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_35_U1_X), .B0_f (new_AGEMA_signal_1937), .B1_t (new_AGEMA_signal_1938), .B1_f (new_AGEMA_signal_1939), .Z0_t (KeyMUX_MUXInst_35_U1_Y), .Z0_f (new_AGEMA_signal_2556), .Z1_t (new_AGEMA_signal_2557), .Z1_f (new_AGEMA_signal_2558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_35_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_35_U1_Y), .A0_f (new_AGEMA_signal_2556), .A1_t (new_AGEMA_signal_2557), .A1_f (new_AGEMA_signal_2558), .B0_t (Key_s0_t[99]), .B0_f (Key_s0_f[99]), .B1_t (Key_s1_t[99]), .B1_f (Key_s1_f[99]), .Z0_t (SelectedKey[35]), .Z0_f (new_AGEMA_signal_2943), .Z1_t (new_AGEMA_signal_2944), .Z1_f (new_AGEMA_signal_2945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_36_U1_XOR1_U1 ( .A0_t (Key_s0_t[100]), .A0_f (Key_s0_f[100]), .A1_t (Key_s1_t[100]), .A1_f (Key_s1_f[100]), .B0_t (Key_s0_t[36]), .B0_f (Key_s0_f[36]), .B1_t (Key_s1_t[36]), .B1_f (Key_s1_f[36]), .Z0_t (KeyMUX_MUXInst_36_U1_X), .Z0_f (new_AGEMA_signal_1946), .Z1_t (new_AGEMA_signal_1947), .Z1_f (new_AGEMA_signal_1948) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_36_U1_X), .B0_f (new_AGEMA_signal_1946), .B1_t (new_AGEMA_signal_1947), .B1_f (new_AGEMA_signal_1948), .Z0_t (KeyMUX_MUXInst_36_U1_Y), .Z0_f (new_AGEMA_signal_2559), .Z1_t (new_AGEMA_signal_2560), .Z1_f (new_AGEMA_signal_2561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_36_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_36_U1_Y), .A0_f (new_AGEMA_signal_2559), .A1_t (new_AGEMA_signal_2560), .A1_f (new_AGEMA_signal_2561), .B0_t (Key_s0_t[100]), .B0_f (Key_s0_f[100]), .B1_t (Key_s1_t[100]), .B1_f (Key_s1_f[100]), .Z0_t (SelectedKey[36]), .Z0_f (new_AGEMA_signal_2946), .Z1_t (new_AGEMA_signal_2947), .Z1_f (new_AGEMA_signal_2948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_37_U1_XOR1_U1 ( .A0_t (Key_s0_t[101]), .A0_f (Key_s0_f[101]), .A1_t (Key_s1_t[101]), .A1_f (Key_s1_f[101]), .B0_t (Key_s0_t[37]), .B0_f (Key_s0_f[37]), .B1_t (Key_s1_t[37]), .B1_f (Key_s1_f[37]), .Z0_t (KeyMUX_MUXInst_37_U1_X), .Z0_f (new_AGEMA_signal_1955), .Z1_t (new_AGEMA_signal_1956), .Z1_f (new_AGEMA_signal_1957) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_37_U1_X), .B0_f (new_AGEMA_signal_1955), .B1_t (new_AGEMA_signal_1956), .B1_f (new_AGEMA_signal_1957), .Z0_t (KeyMUX_MUXInst_37_U1_Y), .Z0_f (new_AGEMA_signal_2562), .Z1_t (new_AGEMA_signal_2563), .Z1_f (new_AGEMA_signal_2564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_37_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_37_U1_Y), .A0_f (new_AGEMA_signal_2562), .A1_t (new_AGEMA_signal_2563), .A1_f (new_AGEMA_signal_2564), .B0_t (Key_s0_t[101]), .B0_f (Key_s0_f[101]), .B1_t (Key_s1_t[101]), .B1_f (Key_s1_f[101]), .Z0_t (SelectedKey[37]), .Z0_f (new_AGEMA_signal_2949), .Z1_t (new_AGEMA_signal_2950), .Z1_f (new_AGEMA_signal_2951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_38_U1_XOR1_U1 ( .A0_t (Key_s0_t[102]), .A0_f (Key_s0_f[102]), .A1_t (Key_s1_t[102]), .A1_f (Key_s1_f[102]), .B0_t (Key_s0_t[38]), .B0_f (Key_s0_f[38]), .B1_t (Key_s1_t[38]), .B1_f (Key_s1_f[38]), .Z0_t (KeyMUX_MUXInst_38_U1_X), .Z0_f (new_AGEMA_signal_1964), .Z1_t (new_AGEMA_signal_1965), .Z1_f (new_AGEMA_signal_1966) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_38_U1_X), .B0_f (new_AGEMA_signal_1964), .B1_t (new_AGEMA_signal_1965), .B1_f (new_AGEMA_signal_1966), .Z0_t (KeyMUX_MUXInst_38_U1_Y), .Z0_f (new_AGEMA_signal_2565), .Z1_t (new_AGEMA_signal_2566), .Z1_f (new_AGEMA_signal_2567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_38_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_38_U1_Y), .A0_f (new_AGEMA_signal_2565), .A1_t (new_AGEMA_signal_2566), .A1_f (new_AGEMA_signal_2567), .B0_t (Key_s0_t[102]), .B0_f (Key_s0_f[102]), .B1_t (Key_s1_t[102]), .B1_f (Key_s1_f[102]), .Z0_t (SelectedKey[38]), .Z0_f (new_AGEMA_signal_2952), .Z1_t (new_AGEMA_signal_2953), .Z1_f (new_AGEMA_signal_2954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_39_U1_XOR1_U1 ( .A0_t (Key_s0_t[103]), .A0_f (Key_s0_f[103]), .A1_t (Key_s1_t[103]), .A1_f (Key_s1_f[103]), .B0_t (Key_s0_t[39]), .B0_f (Key_s0_f[39]), .B1_t (Key_s1_t[39]), .B1_f (Key_s1_f[39]), .Z0_t (KeyMUX_MUXInst_39_U1_X), .Z0_f (new_AGEMA_signal_1973), .Z1_t (new_AGEMA_signal_1974), .Z1_f (new_AGEMA_signal_1975) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_39_U1_X), .B0_f (new_AGEMA_signal_1973), .B1_t (new_AGEMA_signal_1974), .B1_f (new_AGEMA_signal_1975), .Z0_t (KeyMUX_MUXInst_39_U1_Y), .Z0_f (new_AGEMA_signal_2568), .Z1_t (new_AGEMA_signal_2569), .Z1_f (new_AGEMA_signal_2570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_39_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_39_U1_Y), .A0_f (new_AGEMA_signal_2568), .A1_t (new_AGEMA_signal_2569), .A1_f (new_AGEMA_signal_2570), .B0_t (Key_s0_t[103]), .B0_f (Key_s0_f[103]), .B1_t (Key_s1_t[103]), .B1_f (Key_s1_f[103]), .Z0_t (SelectedKey[39]), .Z0_f (new_AGEMA_signal_2955), .Z1_t (new_AGEMA_signal_2956), .Z1_f (new_AGEMA_signal_2957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_40_U1_XOR1_U1 ( .A0_t (Key_s0_t[104]), .A0_f (Key_s0_f[104]), .A1_t (Key_s1_t[104]), .A1_f (Key_s1_f[104]), .B0_t (Key_s0_t[40]), .B0_f (Key_s0_f[40]), .B1_t (Key_s1_t[40]), .B1_f (Key_s1_f[40]), .Z0_t (KeyMUX_MUXInst_40_U1_X), .Z0_f (new_AGEMA_signal_1982), .Z1_t (new_AGEMA_signal_1983), .Z1_f (new_AGEMA_signal_1984) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_40_U1_X), .B0_f (new_AGEMA_signal_1982), .B1_t (new_AGEMA_signal_1983), .B1_f (new_AGEMA_signal_1984), .Z0_t (KeyMUX_MUXInst_40_U1_Y), .Z0_f (new_AGEMA_signal_2571), .Z1_t (new_AGEMA_signal_2572), .Z1_f (new_AGEMA_signal_2573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_40_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_40_U1_Y), .A0_f (new_AGEMA_signal_2571), .A1_t (new_AGEMA_signal_2572), .A1_f (new_AGEMA_signal_2573), .B0_t (Key_s0_t[104]), .B0_f (Key_s0_f[104]), .B1_t (Key_s1_t[104]), .B1_f (Key_s1_f[104]), .Z0_t (SelectedKey[40]), .Z0_f (new_AGEMA_signal_2958), .Z1_t (new_AGEMA_signal_2959), .Z1_f (new_AGEMA_signal_2960) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_41_U1_XOR1_U1 ( .A0_t (Key_s0_t[105]), .A0_f (Key_s0_f[105]), .A1_t (Key_s1_t[105]), .A1_f (Key_s1_f[105]), .B0_t (Key_s0_t[41]), .B0_f (Key_s0_f[41]), .B1_t (Key_s1_t[41]), .B1_f (Key_s1_f[41]), .Z0_t (KeyMUX_MUXInst_41_U1_X), .Z0_f (new_AGEMA_signal_1991), .Z1_t (new_AGEMA_signal_1992), .Z1_f (new_AGEMA_signal_1993) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_41_U1_X), .B0_f (new_AGEMA_signal_1991), .B1_t (new_AGEMA_signal_1992), .B1_f (new_AGEMA_signal_1993), .Z0_t (KeyMUX_MUXInst_41_U1_Y), .Z0_f (new_AGEMA_signal_2574), .Z1_t (new_AGEMA_signal_2575), .Z1_f (new_AGEMA_signal_2576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_41_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_41_U1_Y), .A0_f (new_AGEMA_signal_2574), .A1_t (new_AGEMA_signal_2575), .A1_f (new_AGEMA_signal_2576), .B0_t (Key_s0_t[105]), .B0_f (Key_s0_f[105]), .B1_t (Key_s1_t[105]), .B1_f (Key_s1_f[105]), .Z0_t (SelectedKey[41]), .Z0_f (new_AGEMA_signal_2961), .Z1_t (new_AGEMA_signal_2962), .Z1_f (new_AGEMA_signal_2963) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_42_U1_XOR1_U1 ( .A0_t (Key_s0_t[106]), .A0_f (Key_s0_f[106]), .A1_t (Key_s1_t[106]), .A1_f (Key_s1_f[106]), .B0_t (Key_s0_t[42]), .B0_f (Key_s0_f[42]), .B1_t (Key_s1_t[42]), .B1_f (Key_s1_f[42]), .Z0_t (KeyMUX_MUXInst_42_U1_X), .Z0_f (new_AGEMA_signal_2000), .Z1_t (new_AGEMA_signal_2001), .Z1_f (new_AGEMA_signal_2002) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_42_U1_X), .B0_f (new_AGEMA_signal_2000), .B1_t (new_AGEMA_signal_2001), .B1_f (new_AGEMA_signal_2002), .Z0_t (KeyMUX_MUXInst_42_U1_Y), .Z0_f (new_AGEMA_signal_2577), .Z1_t (new_AGEMA_signal_2578), .Z1_f (new_AGEMA_signal_2579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_42_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_42_U1_Y), .A0_f (new_AGEMA_signal_2577), .A1_t (new_AGEMA_signal_2578), .A1_f (new_AGEMA_signal_2579), .B0_t (Key_s0_t[106]), .B0_f (Key_s0_f[106]), .B1_t (Key_s1_t[106]), .B1_f (Key_s1_f[106]), .Z0_t (SelectedKey[42]), .Z0_f (new_AGEMA_signal_2964), .Z1_t (new_AGEMA_signal_2965), .Z1_f (new_AGEMA_signal_2966) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_43_U1_XOR1_U1 ( .A0_t (Key_s0_t[107]), .A0_f (Key_s0_f[107]), .A1_t (Key_s1_t[107]), .A1_f (Key_s1_f[107]), .B0_t (Key_s0_t[43]), .B0_f (Key_s0_f[43]), .B1_t (Key_s1_t[43]), .B1_f (Key_s1_f[43]), .Z0_t (KeyMUX_MUXInst_43_U1_X), .Z0_f (new_AGEMA_signal_2009), .Z1_t (new_AGEMA_signal_2010), .Z1_f (new_AGEMA_signal_2011) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_43_U1_X), .B0_f (new_AGEMA_signal_2009), .B1_t (new_AGEMA_signal_2010), .B1_f (new_AGEMA_signal_2011), .Z0_t (KeyMUX_MUXInst_43_U1_Y), .Z0_f (new_AGEMA_signal_2580), .Z1_t (new_AGEMA_signal_2581), .Z1_f (new_AGEMA_signal_2582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_43_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_43_U1_Y), .A0_f (new_AGEMA_signal_2580), .A1_t (new_AGEMA_signal_2581), .A1_f (new_AGEMA_signal_2582), .B0_t (Key_s0_t[107]), .B0_f (Key_s0_f[107]), .B1_t (Key_s1_t[107]), .B1_f (Key_s1_f[107]), .Z0_t (SelectedKey[43]), .Z0_f (new_AGEMA_signal_2967), .Z1_t (new_AGEMA_signal_2968), .Z1_f (new_AGEMA_signal_2969) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_44_U1_XOR1_U1 ( .A0_t (Key_s0_t[108]), .A0_f (Key_s0_f[108]), .A1_t (Key_s1_t[108]), .A1_f (Key_s1_f[108]), .B0_t (Key_s0_t[44]), .B0_f (Key_s0_f[44]), .B1_t (Key_s1_t[44]), .B1_f (Key_s1_f[44]), .Z0_t (KeyMUX_MUXInst_44_U1_X), .Z0_f (new_AGEMA_signal_2018), .Z1_t (new_AGEMA_signal_2019), .Z1_f (new_AGEMA_signal_2020) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_44_U1_X), .B0_f (new_AGEMA_signal_2018), .B1_t (new_AGEMA_signal_2019), .B1_f (new_AGEMA_signal_2020), .Z0_t (KeyMUX_MUXInst_44_U1_Y), .Z0_f (new_AGEMA_signal_2583), .Z1_t (new_AGEMA_signal_2584), .Z1_f (new_AGEMA_signal_2585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_44_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_44_U1_Y), .A0_f (new_AGEMA_signal_2583), .A1_t (new_AGEMA_signal_2584), .A1_f (new_AGEMA_signal_2585), .B0_t (Key_s0_t[108]), .B0_f (Key_s0_f[108]), .B1_t (Key_s1_t[108]), .B1_f (Key_s1_f[108]), .Z0_t (SelectedKey[44]), .Z0_f (new_AGEMA_signal_2970), .Z1_t (new_AGEMA_signal_2971), .Z1_f (new_AGEMA_signal_2972) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_45_U1_XOR1_U1 ( .A0_t (Key_s0_t[109]), .A0_f (Key_s0_f[109]), .A1_t (Key_s1_t[109]), .A1_f (Key_s1_f[109]), .B0_t (Key_s0_t[45]), .B0_f (Key_s0_f[45]), .B1_t (Key_s1_t[45]), .B1_f (Key_s1_f[45]), .Z0_t (KeyMUX_MUXInst_45_U1_X), .Z0_f (new_AGEMA_signal_2027), .Z1_t (new_AGEMA_signal_2028), .Z1_f (new_AGEMA_signal_2029) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_45_U1_X), .B0_f (new_AGEMA_signal_2027), .B1_t (new_AGEMA_signal_2028), .B1_f (new_AGEMA_signal_2029), .Z0_t (KeyMUX_MUXInst_45_U1_Y), .Z0_f (new_AGEMA_signal_2586), .Z1_t (new_AGEMA_signal_2587), .Z1_f (new_AGEMA_signal_2588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_45_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_45_U1_Y), .A0_f (new_AGEMA_signal_2586), .A1_t (new_AGEMA_signal_2587), .A1_f (new_AGEMA_signal_2588), .B0_t (Key_s0_t[109]), .B0_f (Key_s0_f[109]), .B1_t (Key_s1_t[109]), .B1_f (Key_s1_f[109]), .Z0_t (SelectedKey[45]), .Z0_f (new_AGEMA_signal_2973), .Z1_t (new_AGEMA_signal_2974), .Z1_f (new_AGEMA_signal_2975) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_46_U1_XOR1_U1 ( .A0_t (Key_s0_t[110]), .A0_f (Key_s0_f[110]), .A1_t (Key_s1_t[110]), .A1_f (Key_s1_f[110]), .B0_t (Key_s0_t[46]), .B0_f (Key_s0_f[46]), .B1_t (Key_s1_t[46]), .B1_f (Key_s1_f[46]), .Z0_t (KeyMUX_MUXInst_46_U1_X), .Z0_f (new_AGEMA_signal_2036), .Z1_t (new_AGEMA_signal_2037), .Z1_f (new_AGEMA_signal_2038) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_46_U1_X), .B0_f (new_AGEMA_signal_2036), .B1_t (new_AGEMA_signal_2037), .B1_f (new_AGEMA_signal_2038), .Z0_t (KeyMUX_MUXInst_46_U1_Y), .Z0_f (new_AGEMA_signal_2589), .Z1_t (new_AGEMA_signal_2590), .Z1_f (new_AGEMA_signal_2591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_46_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_46_U1_Y), .A0_f (new_AGEMA_signal_2589), .A1_t (new_AGEMA_signal_2590), .A1_f (new_AGEMA_signal_2591), .B0_t (Key_s0_t[110]), .B0_f (Key_s0_f[110]), .B1_t (Key_s1_t[110]), .B1_f (Key_s1_f[110]), .Z0_t (SelectedKey[46]), .Z0_f (new_AGEMA_signal_2976), .Z1_t (new_AGEMA_signal_2977), .Z1_f (new_AGEMA_signal_2978) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_47_U1_XOR1_U1 ( .A0_t (Key_s0_t[111]), .A0_f (Key_s0_f[111]), .A1_t (Key_s1_t[111]), .A1_f (Key_s1_f[111]), .B0_t (Key_s0_t[47]), .B0_f (Key_s0_f[47]), .B1_t (Key_s1_t[47]), .B1_f (Key_s1_f[47]), .Z0_t (KeyMUX_MUXInst_47_U1_X), .Z0_f (new_AGEMA_signal_2045), .Z1_t (new_AGEMA_signal_2046), .Z1_f (new_AGEMA_signal_2047) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_47_U1_X), .B0_f (new_AGEMA_signal_2045), .B1_t (new_AGEMA_signal_2046), .B1_f (new_AGEMA_signal_2047), .Z0_t (KeyMUX_MUXInst_47_U1_Y), .Z0_f (new_AGEMA_signal_2592), .Z1_t (new_AGEMA_signal_2593), .Z1_f (new_AGEMA_signal_2594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_47_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_47_U1_Y), .A0_f (new_AGEMA_signal_2592), .A1_t (new_AGEMA_signal_2593), .A1_f (new_AGEMA_signal_2594), .B0_t (Key_s0_t[111]), .B0_f (Key_s0_f[111]), .B1_t (Key_s1_t[111]), .B1_f (Key_s1_f[111]), .Z0_t (SelectedKey[47]), .Z0_f (new_AGEMA_signal_2979), .Z1_t (new_AGEMA_signal_2980), .Z1_f (new_AGEMA_signal_2981) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_48_U1_XOR1_U1 ( .A0_t (Key_s0_t[112]), .A0_f (Key_s0_f[112]), .A1_t (Key_s1_t[112]), .A1_f (Key_s1_f[112]), .B0_t (Key_s0_t[48]), .B0_f (Key_s0_f[48]), .B1_t (Key_s1_t[48]), .B1_f (Key_s1_f[48]), .Z0_t (KeyMUX_MUXInst_48_U1_X), .Z0_f (new_AGEMA_signal_2054), .Z1_t (new_AGEMA_signal_2055), .Z1_f (new_AGEMA_signal_2056) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_48_U1_X), .B0_f (new_AGEMA_signal_2054), .B1_t (new_AGEMA_signal_2055), .B1_f (new_AGEMA_signal_2056), .Z0_t (KeyMUX_MUXInst_48_U1_Y), .Z0_f (new_AGEMA_signal_2595), .Z1_t (new_AGEMA_signal_2596), .Z1_f (new_AGEMA_signal_2597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_48_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_48_U1_Y), .A0_f (new_AGEMA_signal_2595), .A1_t (new_AGEMA_signal_2596), .A1_f (new_AGEMA_signal_2597), .B0_t (Key_s0_t[112]), .B0_f (Key_s0_f[112]), .B1_t (Key_s1_t[112]), .B1_f (Key_s1_f[112]), .Z0_t (SelectedKey[48]), .Z0_f (new_AGEMA_signal_2982), .Z1_t (new_AGEMA_signal_2983), .Z1_f (new_AGEMA_signal_2984) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_49_U1_XOR1_U1 ( .A0_t (Key_s0_t[113]), .A0_f (Key_s0_f[113]), .A1_t (Key_s1_t[113]), .A1_f (Key_s1_f[113]), .B0_t (Key_s0_t[49]), .B0_f (Key_s0_f[49]), .B1_t (Key_s1_t[49]), .B1_f (Key_s1_f[49]), .Z0_t (KeyMUX_MUXInst_49_U1_X), .Z0_f (new_AGEMA_signal_2063), .Z1_t (new_AGEMA_signal_2064), .Z1_f (new_AGEMA_signal_2065) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_49_U1_X), .B0_f (new_AGEMA_signal_2063), .B1_t (new_AGEMA_signal_2064), .B1_f (new_AGEMA_signal_2065), .Z0_t (KeyMUX_MUXInst_49_U1_Y), .Z0_f (new_AGEMA_signal_2598), .Z1_t (new_AGEMA_signal_2599), .Z1_f (new_AGEMA_signal_2600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_49_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_49_U1_Y), .A0_f (new_AGEMA_signal_2598), .A1_t (new_AGEMA_signal_2599), .A1_f (new_AGEMA_signal_2600), .B0_t (Key_s0_t[113]), .B0_f (Key_s0_f[113]), .B1_t (Key_s1_t[113]), .B1_f (Key_s1_f[113]), .Z0_t (SelectedKey[49]), .Z0_f (new_AGEMA_signal_2985), .Z1_t (new_AGEMA_signal_2986), .Z1_f (new_AGEMA_signal_2987) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_50_U1_XOR1_U1 ( .A0_t (Key_s0_t[114]), .A0_f (Key_s0_f[114]), .A1_t (Key_s1_t[114]), .A1_f (Key_s1_f[114]), .B0_t (Key_s0_t[50]), .B0_f (Key_s0_f[50]), .B1_t (Key_s1_t[50]), .B1_f (Key_s1_f[50]), .Z0_t (KeyMUX_MUXInst_50_U1_X), .Z0_f (new_AGEMA_signal_2072), .Z1_t (new_AGEMA_signal_2073), .Z1_f (new_AGEMA_signal_2074) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_50_U1_X), .B0_f (new_AGEMA_signal_2072), .B1_t (new_AGEMA_signal_2073), .B1_f (new_AGEMA_signal_2074), .Z0_t (KeyMUX_MUXInst_50_U1_Y), .Z0_f (new_AGEMA_signal_2601), .Z1_t (new_AGEMA_signal_2602), .Z1_f (new_AGEMA_signal_2603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_50_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_50_U1_Y), .A0_f (new_AGEMA_signal_2601), .A1_t (new_AGEMA_signal_2602), .A1_f (new_AGEMA_signal_2603), .B0_t (Key_s0_t[114]), .B0_f (Key_s0_f[114]), .B1_t (Key_s1_t[114]), .B1_f (Key_s1_f[114]), .Z0_t (SelectedKey[50]), .Z0_f (new_AGEMA_signal_2988), .Z1_t (new_AGEMA_signal_2989), .Z1_f (new_AGEMA_signal_2990) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_51_U1_XOR1_U1 ( .A0_t (Key_s0_t[115]), .A0_f (Key_s0_f[115]), .A1_t (Key_s1_t[115]), .A1_f (Key_s1_f[115]), .B0_t (Key_s0_t[51]), .B0_f (Key_s0_f[51]), .B1_t (Key_s1_t[51]), .B1_f (Key_s1_f[51]), .Z0_t (KeyMUX_MUXInst_51_U1_X), .Z0_f (new_AGEMA_signal_2081), .Z1_t (new_AGEMA_signal_2082), .Z1_f (new_AGEMA_signal_2083) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_51_U1_X), .B0_f (new_AGEMA_signal_2081), .B1_t (new_AGEMA_signal_2082), .B1_f (new_AGEMA_signal_2083), .Z0_t (KeyMUX_MUXInst_51_U1_Y), .Z0_f (new_AGEMA_signal_2604), .Z1_t (new_AGEMA_signal_2605), .Z1_f (new_AGEMA_signal_2606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_51_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_51_U1_Y), .A0_f (new_AGEMA_signal_2604), .A1_t (new_AGEMA_signal_2605), .A1_f (new_AGEMA_signal_2606), .B0_t (Key_s0_t[115]), .B0_f (Key_s0_f[115]), .B1_t (Key_s1_t[115]), .B1_f (Key_s1_f[115]), .Z0_t (SelectedKey[51]), .Z0_f (new_AGEMA_signal_2991), .Z1_t (new_AGEMA_signal_2992), .Z1_f (new_AGEMA_signal_2993) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_52_U1_XOR1_U1 ( .A0_t (Key_s0_t[116]), .A0_f (Key_s0_f[116]), .A1_t (Key_s1_t[116]), .A1_f (Key_s1_f[116]), .B0_t (Key_s0_t[52]), .B0_f (Key_s0_f[52]), .B1_t (Key_s1_t[52]), .B1_f (Key_s1_f[52]), .Z0_t (KeyMUX_MUXInst_52_U1_X), .Z0_f (new_AGEMA_signal_2090), .Z1_t (new_AGEMA_signal_2091), .Z1_f (new_AGEMA_signal_2092) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_52_U1_X), .B0_f (new_AGEMA_signal_2090), .B1_t (new_AGEMA_signal_2091), .B1_f (new_AGEMA_signal_2092), .Z0_t (KeyMUX_MUXInst_52_U1_Y), .Z0_f (new_AGEMA_signal_2607), .Z1_t (new_AGEMA_signal_2608), .Z1_f (new_AGEMA_signal_2609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_52_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_52_U1_Y), .A0_f (new_AGEMA_signal_2607), .A1_t (new_AGEMA_signal_2608), .A1_f (new_AGEMA_signal_2609), .B0_t (Key_s0_t[116]), .B0_f (Key_s0_f[116]), .B1_t (Key_s1_t[116]), .B1_f (Key_s1_f[116]), .Z0_t (SelectedKey[52]), .Z0_f (new_AGEMA_signal_2994), .Z1_t (new_AGEMA_signal_2995), .Z1_f (new_AGEMA_signal_2996) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_53_U1_XOR1_U1 ( .A0_t (Key_s0_t[117]), .A0_f (Key_s0_f[117]), .A1_t (Key_s1_t[117]), .A1_f (Key_s1_f[117]), .B0_t (Key_s0_t[53]), .B0_f (Key_s0_f[53]), .B1_t (Key_s1_t[53]), .B1_f (Key_s1_f[53]), .Z0_t (KeyMUX_MUXInst_53_U1_X), .Z0_f (new_AGEMA_signal_2099), .Z1_t (new_AGEMA_signal_2100), .Z1_f (new_AGEMA_signal_2101) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_53_U1_X), .B0_f (new_AGEMA_signal_2099), .B1_t (new_AGEMA_signal_2100), .B1_f (new_AGEMA_signal_2101), .Z0_t (KeyMUX_MUXInst_53_U1_Y), .Z0_f (new_AGEMA_signal_2610), .Z1_t (new_AGEMA_signal_2611), .Z1_f (new_AGEMA_signal_2612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_53_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_53_U1_Y), .A0_f (new_AGEMA_signal_2610), .A1_t (new_AGEMA_signal_2611), .A1_f (new_AGEMA_signal_2612), .B0_t (Key_s0_t[117]), .B0_f (Key_s0_f[117]), .B1_t (Key_s1_t[117]), .B1_f (Key_s1_f[117]), .Z0_t (SelectedKey[53]), .Z0_f (new_AGEMA_signal_2997), .Z1_t (new_AGEMA_signal_2998), .Z1_f (new_AGEMA_signal_2999) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_54_U1_XOR1_U1 ( .A0_t (Key_s0_t[118]), .A0_f (Key_s0_f[118]), .A1_t (Key_s1_t[118]), .A1_f (Key_s1_f[118]), .B0_t (Key_s0_t[54]), .B0_f (Key_s0_f[54]), .B1_t (Key_s1_t[54]), .B1_f (Key_s1_f[54]), .Z0_t (KeyMUX_MUXInst_54_U1_X), .Z0_f (new_AGEMA_signal_2108), .Z1_t (new_AGEMA_signal_2109), .Z1_f (new_AGEMA_signal_2110) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_54_U1_X), .B0_f (new_AGEMA_signal_2108), .B1_t (new_AGEMA_signal_2109), .B1_f (new_AGEMA_signal_2110), .Z0_t (KeyMUX_MUXInst_54_U1_Y), .Z0_f (new_AGEMA_signal_2613), .Z1_t (new_AGEMA_signal_2614), .Z1_f (new_AGEMA_signal_2615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_54_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_54_U1_Y), .A0_f (new_AGEMA_signal_2613), .A1_t (new_AGEMA_signal_2614), .A1_f (new_AGEMA_signal_2615), .B0_t (Key_s0_t[118]), .B0_f (Key_s0_f[118]), .B1_t (Key_s1_t[118]), .B1_f (Key_s1_f[118]), .Z0_t (SelectedKey[54]), .Z0_f (new_AGEMA_signal_3000), .Z1_t (new_AGEMA_signal_3001), .Z1_f (new_AGEMA_signal_3002) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_55_U1_XOR1_U1 ( .A0_t (Key_s0_t[119]), .A0_f (Key_s0_f[119]), .A1_t (Key_s1_t[119]), .A1_f (Key_s1_f[119]), .B0_t (Key_s0_t[55]), .B0_f (Key_s0_f[55]), .B1_t (Key_s1_t[55]), .B1_f (Key_s1_f[55]), .Z0_t (KeyMUX_MUXInst_55_U1_X), .Z0_f (new_AGEMA_signal_2117), .Z1_t (new_AGEMA_signal_2118), .Z1_f (new_AGEMA_signal_2119) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_55_U1_X), .B0_f (new_AGEMA_signal_2117), .B1_t (new_AGEMA_signal_2118), .B1_f (new_AGEMA_signal_2119), .Z0_t (KeyMUX_MUXInst_55_U1_Y), .Z0_f (new_AGEMA_signal_2616), .Z1_t (new_AGEMA_signal_2617), .Z1_f (new_AGEMA_signal_2618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_55_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_55_U1_Y), .A0_f (new_AGEMA_signal_2616), .A1_t (new_AGEMA_signal_2617), .A1_f (new_AGEMA_signal_2618), .B0_t (Key_s0_t[119]), .B0_f (Key_s0_f[119]), .B1_t (Key_s1_t[119]), .B1_f (Key_s1_f[119]), .Z0_t (SelectedKey[55]), .Z0_f (new_AGEMA_signal_3003), .Z1_t (new_AGEMA_signal_3004), .Z1_f (new_AGEMA_signal_3005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_56_U1_XOR1_U1 ( .A0_t (Key_s0_t[120]), .A0_f (Key_s0_f[120]), .A1_t (Key_s1_t[120]), .A1_f (Key_s1_f[120]), .B0_t (Key_s0_t[56]), .B0_f (Key_s0_f[56]), .B1_t (Key_s1_t[56]), .B1_f (Key_s1_f[56]), .Z0_t (KeyMUX_MUXInst_56_U1_X), .Z0_f (new_AGEMA_signal_2126), .Z1_t (new_AGEMA_signal_2127), .Z1_f (new_AGEMA_signal_2128) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_56_U1_X), .B0_f (new_AGEMA_signal_2126), .B1_t (new_AGEMA_signal_2127), .B1_f (new_AGEMA_signal_2128), .Z0_t (KeyMUX_MUXInst_56_U1_Y), .Z0_f (new_AGEMA_signal_2619), .Z1_t (new_AGEMA_signal_2620), .Z1_f (new_AGEMA_signal_2621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_56_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_56_U1_Y), .A0_f (new_AGEMA_signal_2619), .A1_t (new_AGEMA_signal_2620), .A1_f (new_AGEMA_signal_2621), .B0_t (Key_s0_t[120]), .B0_f (Key_s0_f[120]), .B1_t (Key_s1_t[120]), .B1_f (Key_s1_f[120]), .Z0_t (SelectedKey[56]), .Z0_f (new_AGEMA_signal_3006), .Z1_t (new_AGEMA_signal_3007), .Z1_f (new_AGEMA_signal_3008) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_57_U1_XOR1_U1 ( .A0_t (Key_s0_t[121]), .A0_f (Key_s0_f[121]), .A1_t (Key_s1_t[121]), .A1_f (Key_s1_f[121]), .B0_t (Key_s0_t[57]), .B0_f (Key_s0_f[57]), .B1_t (Key_s1_t[57]), .B1_f (Key_s1_f[57]), .Z0_t (KeyMUX_MUXInst_57_U1_X), .Z0_f (new_AGEMA_signal_2135), .Z1_t (new_AGEMA_signal_2136), .Z1_f (new_AGEMA_signal_2137) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_57_U1_X), .B0_f (new_AGEMA_signal_2135), .B1_t (new_AGEMA_signal_2136), .B1_f (new_AGEMA_signal_2137), .Z0_t (KeyMUX_MUXInst_57_U1_Y), .Z0_f (new_AGEMA_signal_2622), .Z1_t (new_AGEMA_signal_2623), .Z1_f (new_AGEMA_signal_2624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_57_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_57_U1_Y), .A0_f (new_AGEMA_signal_2622), .A1_t (new_AGEMA_signal_2623), .A1_f (new_AGEMA_signal_2624), .B0_t (Key_s0_t[121]), .B0_f (Key_s0_f[121]), .B1_t (Key_s1_t[121]), .B1_f (Key_s1_f[121]), .Z0_t (SelectedKey[57]), .Z0_f (new_AGEMA_signal_3009), .Z1_t (new_AGEMA_signal_3010), .Z1_f (new_AGEMA_signal_3011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_58_U1_XOR1_U1 ( .A0_t (Key_s0_t[122]), .A0_f (Key_s0_f[122]), .A1_t (Key_s1_t[122]), .A1_f (Key_s1_f[122]), .B0_t (Key_s0_t[58]), .B0_f (Key_s0_f[58]), .B1_t (Key_s1_t[58]), .B1_f (Key_s1_f[58]), .Z0_t (KeyMUX_MUXInst_58_U1_X), .Z0_f (new_AGEMA_signal_2144), .Z1_t (new_AGEMA_signal_2145), .Z1_f (new_AGEMA_signal_2146) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_58_U1_X), .B0_f (new_AGEMA_signal_2144), .B1_t (new_AGEMA_signal_2145), .B1_f (new_AGEMA_signal_2146), .Z0_t (KeyMUX_MUXInst_58_U1_Y), .Z0_f (new_AGEMA_signal_2625), .Z1_t (new_AGEMA_signal_2626), .Z1_f (new_AGEMA_signal_2627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_58_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_58_U1_Y), .A0_f (new_AGEMA_signal_2625), .A1_t (new_AGEMA_signal_2626), .A1_f (new_AGEMA_signal_2627), .B0_t (Key_s0_t[122]), .B0_f (Key_s0_f[122]), .B1_t (Key_s1_t[122]), .B1_f (Key_s1_f[122]), .Z0_t (SelectedKey[58]), .Z0_f (new_AGEMA_signal_3012), .Z1_t (new_AGEMA_signal_3013), .Z1_f (new_AGEMA_signal_3014) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_59_U1_XOR1_U1 ( .A0_t (Key_s0_t[123]), .A0_f (Key_s0_f[123]), .A1_t (Key_s1_t[123]), .A1_f (Key_s1_f[123]), .B0_t (Key_s0_t[59]), .B0_f (Key_s0_f[59]), .B1_t (Key_s1_t[59]), .B1_f (Key_s1_f[59]), .Z0_t (KeyMUX_MUXInst_59_U1_X), .Z0_f (new_AGEMA_signal_2153), .Z1_t (new_AGEMA_signal_2154), .Z1_f (new_AGEMA_signal_2155) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_59_U1_X), .B0_f (new_AGEMA_signal_2153), .B1_t (new_AGEMA_signal_2154), .B1_f (new_AGEMA_signal_2155), .Z0_t (KeyMUX_MUXInst_59_U1_Y), .Z0_f (new_AGEMA_signal_2628), .Z1_t (new_AGEMA_signal_2629), .Z1_f (new_AGEMA_signal_2630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_59_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_59_U1_Y), .A0_f (new_AGEMA_signal_2628), .A1_t (new_AGEMA_signal_2629), .A1_f (new_AGEMA_signal_2630), .B0_t (Key_s0_t[123]), .B0_f (Key_s0_f[123]), .B1_t (Key_s1_t[123]), .B1_f (Key_s1_f[123]), .Z0_t (SelectedKey[59]), .Z0_f (new_AGEMA_signal_3015), .Z1_t (new_AGEMA_signal_3016), .Z1_f (new_AGEMA_signal_3017) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_60_U1_XOR1_U1 ( .A0_t (Key_s0_t[124]), .A0_f (Key_s0_f[124]), .A1_t (Key_s1_t[124]), .A1_f (Key_s1_f[124]), .B0_t (Key_s0_t[60]), .B0_f (Key_s0_f[60]), .B1_t (Key_s1_t[60]), .B1_f (Key_s1_f[60]), .Z0_t (KeyMUX_MUXInst_60_U1_X), .Z0_f (new_AGEMA_signal_2162), .Z1_t (new_AGEMA_signal_2163), .Z1_f (new_AGEMA_signal_2164) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_60_U1_X), .B0_f (new_AGEMA_signal_2162), .B1_t (new_AGEMA_signal_2163), .B1_f (new_AGEMA_signal_2164), .Z0_t (KeyMUX_MUXInst_60_U1_Y), .Z0_f (new_AGEMA_signal_2631), .Z1_t (new_AGEMA_signal_2632), .Z1_f (new_AGEMA_signal_2633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_60_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_60_U1_Y), .A0_f (new_AGEMA_signal_2631), .A1_t (new_AGEMA_signal_2632), .A1_f (new_AGEMA_signal_2633), .B0_t (Key_s0_t[124]), .B0_f (Key_s0_f[124]), .B1_t (Key_s1_t[124]), .B1_f (Key_s1_f[124]), .Z0_t (SelectedKey[60]), .Z0_f (new_AGEMA_signal_3018), .Z1_t (new_AGEMA_signal_3019), .Z1_f (new_AGEMA_signal_3020) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_61_U1_XOR1_U1 ( .A0_t (Key_s0_t[125]), .A0_f (Key_s0_f[125]), .A1_t (Key_s1_t[125]), .A1_f (Key_s1_f[125]), .B0_t (Key_s0_t[61]), .B0_f (Key_s0_f[61]), .B1_t (Key_s1_t[61]), .B1_f (Key_s1_f[61]), .Z0_t (KeyMUX_MUXInst_61_U1_X), .Z0_f (new_AGEMA_signal_2171), .Z1_t (new_AGEMA_signal_2172), .Z1_f (new_AGEMA_signal_2173) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_61_U1_X), .B0_f (new_AGEMA_signal_2171), .B1_t (new_AGEMA_signal_2172), .B1_f (new_AGEMA_signal_2173), .Z0_t (KeyMUX_MUXInst_61_U1_Y), .Z0_f (new_AGEMA_signal_2634), .Z1_t (new_AGEMA_signal_2635), .Z1_f (new_AGEMA_signal_2636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_61_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_61_U1_Y), .A0_f (new_AGEMA_signal_2634), .A1_t (new_AGEMA_signal_2635), .A1_f (new_AGEMA_signal_2636), .B0_t (Key_s0_t[125]), .B0_f (Key_s0_f[125]), .B1_t (Key_s1_t[125]), .B1_f (Key_s1_f[125]), .Z0_t (SelectedKey[61]), .Z0_f (new_AGEMA_signal_3021), .Z1_t (new_AGEMA_signal_3022), .Z1_f (new_AGEMA_signal_3023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_62_U1_XOR1_U1 ( .A0_t (Key_s0_t[126]), .A0_f (Key_s0_f[126]), .A1_t (Key_s1_t[126]), .A1_f (Key_s1_f[126]), .B0_t (Key_s0_t[62]), .B0_f (Key_s0_f[62]), .B1_t (Key_s1_t[62]), .B1_f (Key_s1_f[62]), .Z0_t (KeyMUX_MUXInst_62_U1_X), .Z0_f (new_AGEMA_signal_2180), .Z1_t (new_AGEMA_signal_2181), .Z1_f (new_AGEMA_signal_2182) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_62_U1_X), .B0_f (new_AGEMA_signal_2180), .B1_t (new_AGEMA_signal_2181), .B1_f (new_AGEMA_signal_2182), .Z0_t (KeyMUX_MUXInst_62_U1_Y), .Z0_f (new_AGEMA_signal_2637), .Z1_t (new_AGEMA_signal_2638), .Z1_f (new_AGEMA_signal_2639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_62_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_62_U1_Y), .A0_f (new_AGEMA_signal_2637), .A1_t (new_AGEMA_signal_2638), .A1_f (new_AGEMA_signal_2639), .B0_t (Key_s0_t[126]), .B0_f (Key_s0_f[126]), .B1_t (Key_s1_t[126]), .B1_f (Key_s1_f[126]), .Z0_t (SelectedKey[62]), .Z0_f (new_AGEMA_signal_3024), .Z1_t (new_AGEMA_signal_3025), .Z1_f (new_AGEMA_signal_3026) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_63_U1_XOR1_U1 ( .A0_t (Key_s0_t[127]), .A0_f (Key_s0_f[127]), .A1_t (Key_s1_t[127]), .A1_f (Key_s1_f[127]), .B0_t (Key_s0_t[63]), .B0_f (Key_s0_f[63]), .B1_t (Key_s1_t[63]), .B1_f (Key_s1_f[63]), .Z0_t (KeyMUX_MUXInst_63_U1_X), .Z0_f (new_AGEMA_signal_2189), .Z1_t (new_AGEMA_signal_2190), .Z1_f (new_AGEMA_signal_2191) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selects[0]), .A1_f (new_AGEMA_signal_2208), .B0_t (KeyMUX_MUXInst_63_U1_X), .B0_f (new_AGEMA_signal_2189), .B1_t (new_AGEMA_signal_2190), .B1_f (new_AGEMA_signal_2191), .Z0_t (KeyMUX_MUXInst_63_U1_Y), .Z0_f (new_AGEMA_signal_2640), .Z1_t (new_AGEMA_signal_2641), .Z1_f (new_AGEMA_signal_2642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyMUX_MUXInst_63_U1_XOR2_U1 ( .A0_t (KeyMUX_MUXInst_63_U1_Y), .A0_f (new_AGEMA_signal_2640), .A1_t (new_AGEMA_signal_2641), .A1_f (new_AGEMA_signal_2642), .B0_t (Key_s0_t[127]), .B0_f (Key_s0_f[127]), .B1_t (Key_s1_t[127]), .B1_f (Key_s1_f[127]), .Z0_t (SelectedKey[63]), .Z0_f (new_AGEMA_signal_3027), .Z1_t (new_AGEMA_signal_3028), .Z1_f (new_AGEMA_signal_3029) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_0_U1 ( .A0_t (FSMReg[0]), .A0_f (new_AGEMA_signal_2192), .B0_t (rst_t), .B0_f (rst_f), .Z0_t (RoundConstant_0), .Z0_f (new_AGEMA_signal_2194) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_1_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (FSMReg[1]), .B0_f (new_AGEMA_signal_2195), .Z0_t (FSMUpdate[0]), .Z0_f (new_AGEMA_signal_2196) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_2_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (FSMReg[2]), .B0_f (new_AGEMA_signal_2197), .Z0_t (FSMUpdate[1]), .Z0_f (new_AGEMA_signal_2198) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_3_U1 ( .A0_t (FSMReg[3]), .A0_f (new_AGEMA_signal_2199), .B0_t (rst_t), .B0_f (rst_f), .Z0_t (RoundConstant_4_), .Z0_f (new_AGEMA_signal_2200) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_4_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (FSMReg[4]), .B0_f (new_AGEMA_signal_2201), .Z0_t (FSMUpdate[3]), .Z0_f (new_AGEMA_signal_2202) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_5_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (FSMReg[5]), .B0_f (new_AGEMA_signal_2203), .Z0_t (FSMUpdate[4]), .Z0_f (new_AGEMA_signal_2204) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMMUX_MUXInst_6_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (FSMReg[6]), .B0_f (new_AGEMA_signal_2205), .Z0_t (FSMUpdate[5]), .Z0_f (new_AGEMA_signal_2206) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) FSMUpdateInst_U2 ( .A0_t (FSMUpdate[0]), .A0_f (new_AGEMA_signal_2196), .B0_t (RoundConstant_0), .B0_f (new_AGEMA_signal_2194), .Z0_t (FSMReg[2]), .Z0_f (new_AGEMA_signal_2197) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) FSMUpdateInst_U1 ( .A0_t (FSMUpdate[3]), .A0_f (new_AGEMA_signal_2202), .B0_t (RoundConstant_4_), .B0_f (new_AGEMA_signal_2200), .Z0_t (FSMReg[6]), .Z0_f (new_AGEMA_signal_2205) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMSignalsInst_U6 ( .A0_t (RoundConstant_0), .A0_f (new_AGEMA_signal_2194), .B0_t (FSMSignalsInst_n5), .B0_f (new_AGEMA_signal_3319), .Z0_t (done_t), .Z0_f (done_f) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_U5 ( .A0_t (FSMSignalsInst_n4), .A0_f (new_AGEMA_signal_2645), .B0_t (FSMSignalsInst_n3), .B0_f (new_AGEMA_signal_3030), .Z0_t (FSMSignalsInst_n5), .Z0_f (new_AGEMA_signal_3319) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_U4 ( .A0_t (FSMSignalsInst_n2), .A0_f (new_AGEMA_signal_2644), .B0_t (FSMSignalsInst_n1), .B0_f (new_AGEMA_signal_2643), .Z0_t (FSMSignalsInst_n3), .Z0_f (new_AGEMA_signal_3030) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_U3 ( .A0_t (RoundConstant_4_), .A0_f (new_AGEMA_signal_2200), .B0_t (FSMUpdate[0]), .B0_f (new_AGEMA_signal_2196), .Z0_t (FSMSignalsInst_n1), .Z0_f (new_AGEMA_signal_2643) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_U2 ( .A0_t (FSMUpdate[4]), .A0_f (new_AGEMA_signal_2204), .B0_t (FSMUpdate[3]), .B0_f (new_AGEMA_signal_2202), .Z0_t (FSMSignalsInst_n2), .Z0_f (new_AGEMA_signal_2644) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_U1 ( .A0_t (FSMUpdate[1]), .A0_f (new_AGEMA_signal_2198), .B0_t (FSMUpdate[5]), .B0_f (new_AGEMA_signal_2206), .Z0_t (FSMSignalsInst_n4), .Z0_f (new_AGEMA_signal_2645) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) selectsMUX_MUXInst_0_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (selectsReg[0]), .B0_f (new_AGEMA_signal_2207), .Z0_t (selects[0]), .Z0_f (new_AGEMA_signal_2208) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) selectsMUX_MUXInst_1_U2 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (selectsReg[1]), .B0_f (new_AGEMA_signal_2209), .Z0_t (selects[1]), .Z0_f (new_AGEMA_signal_2210) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b0)) selectsUpdateInst_U2 ( .A0_t (selects[1]), .A0_f (new_AGEMA_signal_2210), .B0_t (selects[0]), .B0_f (new_AGEMA_signal_2208), .Z0_t (selectsReg[1]), .Z0_f (new_AGEMA_signal_2209) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_984 ( .A0_t (FSMUpdate[5]), .A0_f (new_AGEMA_signal_2206), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (FSMReg[5]), .Z0_f (new_AGEMA_signal_2203) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_985 ( .A0_t (FSMUpdate[4]), .A0_f (new_AGEMA_signal_2204), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (FSMReg[4]), .Z0_f (new_AGEMA_signal_2201) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_986 ( .A0_t (FSMUpdate[3]), .A0_f (new_AGEMA_signal_2202), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (FSMReg[3]), .Z0_f (new_AGEMA_signal_2199) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_987 ( .A0_t (FSMUpdate[1]), .A0_f (new_AGEMA_signal_2198), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (FSMReg[1]), .Z0_f (new_AGEMA_signal_2195) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_988 ( .A0_t (FSMUpdate[0]), .A0_f (new_AGEMA_signal_2196), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (FSMReg[0]), .Z0_f (new_AGEMA_signal_2192) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_989 ( .A0_t (selects[0]), .A0_f (new_AGEMA_signal_2208), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (selectsReg[0]), .Z0_f (new_AGEMA_signal_2207) ) ;

    /* register cells */
endmodule
